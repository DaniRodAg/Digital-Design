`timescale 1ns/1ps

module FA_8B_TB();

reg[7:0] A, B;
wire[7:0] S;
wire Cout;
wire Cin = 1'b0;

FA_8B duv
(
	.A(A),
	.B(B),
	.S(S),
	
	.Cin(Cin),
	.Cout(Cout)
);

initial
begin
A = 8'h0; B = 8'h0; #100;
A = 8'h0; B = 8'h1; #100;
A = 8'h0; B = 8'h2; #100;
A = 8'h0; B = 8'h3; #100;
A = 8'h0; B = 8'h4; #100;
A = 8'h0; B = 8'h5; #100;
A = 8'h0; B = 8'h6; #100;
A = 8'h0; B = 8'h7; #100;
A = 8'h0; B = 8'h8; #100;
A = 8'h0; B = 8'h9; #100;
A = 8'h0; B = 8'hA; #100;
A = 8'h0; B = 8'hB; #100;
A = 8'h0; B = 8'hC; #100;
A = 8'h0; B = 8'hD; #100;
A = 8'h0; B = 8'hE; #100;
A = 8'h0; B = 8'hF; #100;
A = 8'h0; B = 8'h10; #100;
A = 8'h0; B = 8'h11; #100;
A = 8'h0; B = 8'h12; #100;
A = 8'h0; B = 8'h13; #100;
A = 8'h0; B = 8'h14; #100;
A = 8'h0; B = 8'h15; #100;
A = 8'h0; B = 8'h16; #100;
A = 8'h0; B = 8'h17; #100;
A = 8'h0; B = 8'h18; #100;
A = 8'h0; B = 8'h19; #100;
A = 8'h0; B = 8'h1A; #100;
A = 8'h0; B = 8'h1B; #100;
A = 8'h0; B = 8'h1C; #100;
A = 8'h0; B = 8'h1D; #100;
A = 8'h0; B = 8'h1E; #100;
A = 8'h0; B = 8'h1F; #100;
A = 8'h0; B = 8'h20; #100;
A = 8'h0; B = 8'h21; #100;
A = 8'h0; B = 8'h22; #100;
A = 8'h0; B = 8'h23; #100;
A = 8'h0; B = 8'h24; #100;
A = 8'h0; B = 8'h25; #100;
A = 8'h0; B = 8'h26; #100;
A = 8'h0; B = 8'h27; #100;
A = 8'h0; B = 8'h28; #100;
A = 8'h0; B = 8'h29; #100;
A = 8'h0; B = 8'h2A; #100;
A = 8'h0; B = 8'h2B; #100;
A = 8'h0; B = 8'h2C; #100;
A = 8'h0; B = 8'h2D; #100;
A = 8'h0; B = 8'h2E; #100;
A = 8'h0; B = 8'h2F; #100;
A = 8'h0; B = 8'h30; #100;
A = 8'h0; B = 8'h31; #100;
A = 8'h0; B = 8'h32; #100;
A = 8'h0; B = 8'h33; #100;
A = 8'h0; B = 8'h34; #100;
A = 8'h0; B = 8'h35; #100;
A = 8'h0; B = 8'h36; #100;
A = 8'h0; B = 8'h37; #100;
A = 8'h0; B = 8'h38; #100;
A = 8'h0; B = 8'h39; #100;
A = 8'h0; B = 8'h3A; #100;
A = 8'h0; B = 8'h3B; #100;
A = 8'h0; B = 8'h3C; #100;
A = 8'h0; B = 8'h3D; #100;
A = 8'h0; B = 8'h3E; #100;
A = 8'h0; B = 8'h3F; #100;
A = 8'h0; B = 8'h40; #100;
A = 8'h0; B = 8'h41; #100;
A = 8'h0; B = 8'h42; #100;
A = 8'h0; B = 8'h43; #100;
A = 8'h0; B = 8'h44; #100;
A = 8'h0; B = 8'h45; #100;
A = 8'h0; B = 8'h46; #100;
A = 8'h0; B = 8'h47; #100;
A = 8'h0; B = 8'h48; #100;
A = 8'h0; B = 8'h49; #100;
A = 8'h0; B = 8'h4A; #100;
A = 8'h0; B = 8'h4B; #100;
A = 8'h0; B = 8'h4C; #100;
A = 8'h0; B = 8'h4D; #100;
A = 8'h0; B = 8'h4E; #100;
A = 8'h0; B = 8'h4F; #100;
A = 8'h0; B = 8'h50; #100;
A = 8'h0; B = 8'h51; #100;
A = 8'h0; B = 8'h52; #100;
A = 8'h0; B = 8'h53; #100;
A = 8'h0; B = 8'h54; #100;
A = 8'h0; B = 8'h55; #100;
A = 8'h0; B = 8'h56; #100;
A = 8'h0; B = 8'h57; #100;
A = 8'h0; B = 8'h58; #100;
A = 8'h0; B = 8'h59; #100;
A = 8'h0; B = 8'h5A; #100;
A = 8'h0; B = 8'h5B; #100;
A = 8'h0; B = 8'h5C; #100;
A = 8'h0; B = 8'h5D; #100;
A = 8'h0; B = 8'h5E; #100;
A = 8'h0; B = 8'h5F; #100;
A = 8'h0; B = 8'h60; #100;
A = 8'h0; B = 8'h61; #100;
A = 8'h0; B = 8'h62; #100;
A = 8'h0; B = 8'h63; #100;
A = 8'h0; B = 8'h64; #100;
A = 8'h0; B = 8'h65; #100;
A = 8'h0; B = 8'h66; #100;
A = 8'h0; B = 8'h67; #100;
A = 8'h0; B = 8'h68; #100;
A = 8'h0; B = 8'h69; #100;
A = 8'h0; B = 8'h6A; #100;
A = 8'h0; B = 8'h6B; #100;
A = 8'h0; B = 8'h6C; #100;
A = 8'h0; B = 8'h6D; #100;
A = 8'h0; B = 8'h6E; #100;
A = 8'h0; B = 8'h6F; #100;
A = 8'h0; B = 8'h70; #100;
A = 8'h0; B = 8'h71; #100;
A = 8'h0; B = 8'h72; #100;
A = 8'h0; B = 8'h73; #100;
A = 8'h0; B = 8'h74; #100;
A = 8'h0; B = 8'h75; #100;
A = 8'h0; B = 8'h76; #100;
A = 8'h0; B = 8'h77; #100;
A = 8'h0; B = 8'h78; #100;
A = 8'h0; B = 8'h79; #100;
A = 8'h0; B = 8'h7A; #100;
A = 8'h0; B = 8'h7B; #100;
A = 8'h0; B = 8'h7C; #100;
A = 8'h0; B = 8'h7D; #100;
A = 8'h0; B = 8'h7E; #100;
A = 8'h0; B = 8'h7F; #100;
A = 8'h0; B = 8'h80; #100;
A = 8'h0; B = 8'h81; #100;
A = 8'h0; B = 8'h82; #100;
A = 8'h0; B = 8'h83; #100;
A = 8'h0; B = 8'h84; #100;
A = 8'h0; B = 8'h85; #100;
A = 8'h0; B = 8'h86; #100;
A = 8'h0; B = 8'h87; #100;
A = 8'h0; B = 8'h88; #100;
A = 8'h0; B = 8'h89; #100;
A = 8'h0; B = 8'h8A; #100;
A = 8'h0; B = 8'h8B; #100;
A = 8'h0; B = 8'h8C; #100;
A = 8'h0; B = 8'h8D; #100;
A = 8'h0; B = 8'h8E; #100;
A = 8'h0; B = 8'h8F; #100;
A = 8'h0; B = 8'h90; #100;
A = 8'h0; B = 8'h91; #100;
A = 8'h0; B = 8'h92; #100;
A = 8'h0; B = 8'h93; #100;
A = 8'h0; B = 8'h94; #100;
A = 8'h0; B = 8'h95; #100;
A = 8'h0; B = 8'h96; #100;
A = 8'h0; B = 8'h97; #100;
A = 8'h0; B = 8'h98; #100;
A = 8'h0; B = 8'h99; #100;
A = 8'h0; B = 8'h9A; #100;
A = 8'h0; B = 8'h9B; #100;
A = 8'h0; B = 8'h9C; #100;
A = 8'h0; B = 8'h9D; #100;
A = 8'h0; B = 8'h9E; #100;
A = 8'h0; B = 8'h9F; #100;
A = 8'h0; B = 8'hA0; #100;
A = 8'h0; B = 8'hA1; #100;
A = 8'h0; B = 8'hA2; #100;
A = 8'h0; B = 8'hA3; #100;
A = 8'h0; B = 8'hA4; #100;
A = 8'h0; B = 8'hA5; #100;
A = 8'h0; B = 8'hA6; #100;
A = 8'h0; B = 8'hA7; #100;
A = 8'h0; B = 8'hA8; #100;
A = 8'h0; B = 8'hA9; #100;
A = 8'h0; B = 8'hAA; #100;
A = 8'h0; B = 8'hAB; #100;
A = 8'h0; B = 8'hAC; #100;
A = 8'h0; B = 8'hAD; #100;
A = 8'h0; B = 8'hAE; #100;
A = 8'h0; B = 8'hAF; #100;
A = 8'h0; B = 8'hB0; #100;
A = 8'h0; B = 8'hB1; #100;
A = 8'h0; B = 8'hB2; #100;
A = 8'h0; B = 8'hB3; #100;
A = 8'h0; B = 8'hB4; #100;
A = 8'h0; B = 8'hB5; #100;
A = 8'h0; B = 8'hB6; #100;
A = 8'h0; B = 8'hB7; #100;
A = 8'h0; B = 8'hB8; #100;
A = 8'h0; B = 8'hB9; #100;
A = 8'h0; B = 8'hBA; #100;
A = 8'h0; B = 8'hBB; #100;
A = 8'h0; B = 8'hBC; #100;
A = 8'h0; B = 8'hBD; #100;
A = 8'h0; B = 8'hBE; #100;
A = 8'h0; B = 8'hBF; #100;
A = 8'h0; B = 8'hC0; #100;
A = 8'h0; B = 8'hC1; #100;
A = 8'h0; B = 8'hC2; #100;
A = 8'h0; B = 8'hC3; #100;
A = 8'h0; B = 8'hC4; #100;
A = 8'h0; B = 8'hC5; #100;
A = 8'h0; B = 8'hC6; #100;
A = 8'h0; B = 8'hC7; #100;
A = 8'h0; B = 8'hC8; #100;
A = 8'h0; B = 8'hC9; #100;
A = 8'h0; B = 8'hCA; #100;
A = 8'h0; B = 8'hCB; #100;
A = 8'h0; B = 8'hCC; #100;
A = 8'h0; B = 8'hCD; #100;
A = 8'h0; B = 8'hCE; #100;
A = 8'h0; B = 8'hCF; #100;
A = 8'h0; B = 8'hD0; #100;
A = 8'h0; B = 8'hD1; #100;
A = 8'h0; B = 8'hD2; #100;
A = 8'h0; B = 8'hD3; #100;
A = 8'h0; B = 8'hD4; #100;
A = 8'h0; B = 8'hD5; #100;
A = 8'h0; B = 8'hD6; #100;
A = 8'h0; B = 8'hD7; #100;
A = 8'h0; B = 8'hD8; #100;
A = 8'h0; B = 8'hD9; #100;
A = 8'h0; B = 8'hDA; #100;
A = 8'h0; B = 8'hDB; #100;
A = 8'h0; B = 8'hDC; #100;
A = 8'h0; B = 8'hDD; #100;
A = 8'h0; B = 8'hDE; #100;
A = 8'h0; B = 8'hDF; #100;
A = 8'h0; B = 8'hE0; #100;
A = 8'h0; B = 8'hE1; #100;
A = 8'h0; B = 8'hE2; #100;
A = 8'h0; B = 8'hE3; #100;
A = 8'h0; B = 8'hE4; #100;
A = 8'h0; B = 8'hE5; #100;
A = 8'h0; B = 8'hE6; #100;
A = 8'h0; B = 8'hE7; #100;
A = 8'h0; B = 8'hE8; #100;
A = 8'h0; B = 8'hE9; #100;
A = 8'h0; B = 8'hEA; #100;
A = 8'h0; B = 8'hEB; #100;
A = 8'h0; B = 8'hEC; #100;
A = 8'h0; B = 8'hED; #100;
A = 8'h0; B = 8'hEE; #100;
A = 8'h0; B = 8'hEF; #100;
A = 8'h0; B = 8'hF0; #100;
A = 8'h0; B = 8'hF1; #100;
A = 8'h0; B = 8'hF2; #100;
A = 8'h0; B = 8'hF3; #100;
A = 8'h0; B = 8'hF4; #100;
A = 8'h0; B = 8'hF5; #100;
A = 8'h0; B = 8'hF6; #100;
A = 8'h0; B = 8'hF7; #100;
A = 8'h0; B = 8'hF8; #100;
A = 8'h0; B = 8'hF9; #100;
A = 8'h0; B = 8'hFA; #100;
A = 8'h0; B = 8'hFB; #100;
A = 8'h0; B = 8'hFC; #100;
A = 8'h0; B = 8'hFD; #100;
A = 8'h0; B = 8'hFE; #100;
A = 8'h0; B = 8'hFF; #100;
A = 8'h1; B = 8'h0; #100;
A = 8'h1; B = 8'h1; #100;
A = 8'h1; B = 8'h2; #100;
A = 8'h1; B = 8'h3; #100;
A = 8'h1; B = 8'h4; #100;
A = 8'h1; B = 8'h5; #100;
A = 8'h1; B = 8'h6; #100;
A = 8'h1; B = 8'h7; #100;
A = 8'h1; B = 8'h8; #100;
A = 8'h1; B = 8'h9; #100;
A = 8'h1; B = 8'hA; #100;
A = 8'h1; B = 8'hB; #100;
A = 8'h1; B = 8'hC; #100;
A = 8'h1; B = 8'hD; #100;
A = 8'h1; B = 8'hE; #100;
A = 8'h1; B = 8'hF; #100;
A = 8'h1; B = 8'h10; #100;
A = 8'h1; B = 8'h11; #100;
A = 8'h1; B = 8'h12; #100;
A = 8'h1; B = 8'h13; #100;
A = 8'h1; B = 8'h14; #100;
A = 8'h1; B = 8'h15; #100;
A = 8'h1; B = 8'h16; #100;
A = 8'h1; B = 8'h17; #100;
A = 8'h1; B = 8'h18; #100;
A = 8'h1; B = 8'h19; #100;
A = 8'h1; B = 8'h1A; #100;
A = 8'h1; B = 8'h1B; #100;
A = 8'h1; B = 8'h1C; #100;
A = 8'h1; B = 8'h1D; #100;
A = 8'h1; B = 8'h1E; #100;
A = 8'h1; B = 8'h1F; #100;
A = 8'h1; B = 8'h20; #100;
A = 8'h1; B = 8'h21; #100;
A = 8'h1; B = 8'h22; #100;
A = 8'h1; B = 8'h23; #100;
A = 8'h1; B = 8'h24; #100;
A = 8'h1; B = 8'h25; #100;
A = 8'h1; B = 8'h26; #100;
A = 8'h1; B = 8'h27; #100;
A = 8'h1; B = 8'h28; #100;
A = 8'h1; B = 8'h29; #100;
A = 8'h1; B = 8'h2A; #100;
A = 8'h1; B = 8'h2B; #100;
A = 8'h1; B = 8'h2C; #100;
A = 8'h1; B = 8'h2D; #100;
A = 8'h1; B = 8'h2E; #100;
A = 8'h1; B = 8'h2F; #100;
A = 8'h1; B = 8'h30; #100;
A = 8'h1; B = 8'h31; #100;
A = 8'h1; B = 8'h32; #100;
A = 8'h1; B = 8'h33; #100;
A = 8'h1; B = 8'h34; #100;
A = 8'h1; B = 8'h35; #100;
A = 8'h1; B = 8'h36; #100;
A = 8'h1; B = 8'h37; #100;
A = 8'h1; B = 8'h38; #100;
A = 8'h1; B = 8'h39; #100;
A = 8'h1; B = 8'h3A; #100;
A = 8'h1; B = 8'h3B; #100;
A = 8'h1; B = 8'h3C; #100;
A = 8'h1; B = 8'h3D; #100;
A = 8'h1; B = 8'h3E; #100;
A = 8'h1; B = 8'h3F; #100;
A = 8'h1; B = 8'h40; #100;
A = 8'h1; B = 8'h41; #100;
A = 8'h1; B = 8'h42; #100;
A = 8'h1; B = 8'h43; #100;
A = 8'h1; B = 8'h44; #100;
A = 8'h1; B = 8'h45; #100;
A = 8'h1; B = 8'h46; #100;
A = 8'h1; B = 8'h47; #100;
A = 8'h1; B = 8'h48; #100;
A = 8'h1; B = 8'h49; #100;
A = 8'h1; B = 8'h4A; #100;
A = 8'h1; B = 8'h4B; #100;
A = 8'h1; B = 8'h4C; #100;
A = 8'h1; B = 8'h4D; #100;
A = 8'h1; B = 8'h4E; #100;
A = 8'h1; B = 8'h4F; #100;
A = 8'h1; B = 8'h50; #100;
A = 8'h1; B = 8'h51; #100;
A = 8'h1; B = 8'h52; #100;
A = 8'h1; B = 8'h53; #100;
A = 8'h1; B = 8'h54; #100;
A = 8'h1; B = 8'h55; #100;
A = 8'h1; B = 8'h56; #100;
A = 8'h1; B = 8'h57; #100;
A = 8'h1; B = 8'h58; #100;
A = 8'h1; B = 8'h59; #100;
A = 8'h1; B = 8'h5A; #100;
A = 8'h1; B = 8'h5B; #100;
A = 8'h1; B = 8'h5C; #100;
A = 8'h1; B = 8'h5D; #100;
A = 8'h1; B = 8'h5E; #100;
A = 8'h1; B = 8'h5F; #100;
A = 8'h1; B = 8'h60; #100;
A = 8'h1; B = 8'h61; #100;
A = 8'h1; B = 8'h62; #100;
A = 8'h1; B = 8'h63; #100;
A = 8'h1; B = 8'h64; #100;
A = 8'h1; B = 8'h65; #100;
A = 8'h1; B = 8'h66; #100;
A = 8'h1; B = 8'h67; #100;
A = 8'h1; B = 8'h68; #100;
A = 8'h1; B = 8'h69; #100;
A = 8'h1; B = 8'h6A; #100;
A = 8'h1; B = 8'h6B; #100;
A = 8'h1; B = 8'h6C; #100;
A = 8'h1; B = 8'h6D; #100;
A = 8'h1; B = 8'h6E; #100;
A = 8'h1; B = 8'h6F; #100;
A = 8'h1; B = 8'h70; #100;
A = 8'h1; B = 8'h71; #100;
A = 8'h1; B = 8'h72; #100;
A = 8'h1; B = 8'h73; #100;
A = 8'h1; B = 8'h74; #100;
A = 8'h1; B = 8'h75; #100;
A = 8'h1; B = 8'h76; #100;
A = 8'h1; B = 8'h77; #100;
A = 8'h1; B = 8'h78; #100;
A = 8'h1; B = 8'h79; #100;
A = 8'h1; B = 8'h7A; #100;
A = 8'h1; B = 8'h7B; #100;
A = 8'h1; B = 8'h7C; #100;
A = 8'h1; B = 8'h7D; #100;
A = 8'h1; B = 8'h7E; #100;
A = 8'h1; B = 8'h7F; #100;
A = 8'h1; B = 8'h80; #100;
A = 8'h1; B = 8'h81; #100;
A = 8'h1; B = 8'h82; #100;
A = 8'h1; B = 8'h83; #100;
A = 8'h1; B = 8'h84; #100;
A = 8'h1; B = 8'h85; #100;
A = 8'h1; B = 8'h86; #100;
A = 8'h1; B = 8'h87; #100;
A = 8'h1; B = 8'h88; #100;
A = 8'h1; B = 8'h89; #100;
A = 8'h1; B = 8'h8A; #100;
A = 8'h1; B = 8'h8B; #100;
A = 8'h1; B = 8'h8C; #100;
A = 8'h1; B = 8'h8D; #100;
A = 8'h1; B = 8'h8E; #100;
A = 8'h1; B = 8'h8F; #100;
A = 8'h1; B = 8'h90; #100;
A = 8'h1; B = 8'h91; #100;
A = 8'h1; B = 8'h92; #100;
A = 8'h1; B = 8'h93; #100;
A = 8'h1; B = 8'h94; #100;
A = 8'h1; B = 8'h95; #100;
A = 8'h1; B = 8'h96; #100;
A = 8'h1; B = 8'h97; #100;
A = 8'h1; B = 8'h98; #100;
A = 8'h1; B = 8'h99; #100;
A = 8'h1; B = 8'h9A; #100;
A = 8'h1; B = 8'h9B; #100;
A = 8'h1; B = 8'h9C; #100;
A = 8'h1; B = 8'h9D; #100;
A = 8'h1; B = 8'h9E; #100;
A = 8'h1; B = 8'h9F; #100;
A = 8'h1; B = 8'hA0; #100;
A = 8'h1; B = 8'hA1; #100;
A = 8'h1; B = 8'hA2; #100;
A = 8'h1; B = 8'hA3; #100;
A = 8'h1; B = 8'hA4; #100;
A = 8'h1; B = 8'hA5; #100;
A = 8'h1; B = 8'hA6; #100;
A = 8'h1; B = 8'hA7; #100;
A = 8'h1; B = 8'hA8; #100;
A = 8'h1; B = 8'hA9; #100;
A = 8'h1; B = 8'hAA; #100;
A = 8'h1; B = 8'hAB; #100;
A = 8'h1; B = 8'hAC; #100;
A = 8'h1; B = 8'hAD; #100;
A = 8'h1; B = 8'hAE; #100;
A = 8'h1; B = 8'hAF; #100;
A = 8'h1; B = 8'hB0; #100;
A = 8'h1; B = 8'hB1; #100;
A = 8'h1; B = 8'hB2; #100;
A = 8'h1; B = 8'hB3; #100;
A = 8'h1; B = 8'hB4; #100;
A = 8'h1; B = 8'hB5; #100;
A = 8'h1; B = 8'hB6; #100;
A = 8'h1; B = 8'hB7; #100;
A = 8'h1; B = 8'hB8; #100;
A = 8'h1; B = 8'hB9; #100;
A = 8'h1; B = 8'hBA; #100;
A = 8'h1; B = 8'hBB; #100;
A = 8'h1; B = 8'hBC; #100;
A = 8'h1; B = 8'hBD; #100;
A = 8'h1; B = 8'hBE; #100;
A = 8'h1; B = 8'hBF; #100;
A = 8'h1; B = 8'hC0; #100;
A = 8'h1; B = 8'hC1; #100;
A = 8'h1; B = 8'hC2; #100;
A = 8'h1; B = 8'hC3; #100;
A = 8'h1; B = 8'hC4; #100;
A = 8'h1; B = 8'hC5; #100;
A = 8'h1; B = 8'hC6; #100;
A = 8'h1; B = 8'hC7; #100;
A = 8'h1; B = 8'hC8; #100;
A = 8'h1; B = 8'hC9; #100;
A = 8'h1; B = 8'hCA; #100;
A = 8'h1; B = 8'hCB; #100;
A = 8'h1; B = 8'hCC; #100;
A = 8'h1; B = 8'hCD; #100;
A = 8'h1; B = 8'hCE; #100;
A = 8'h1; B = 8'hCF; #100;
A = 8'h1; B = 8'hD0; #100;
A = 8'h1; B = 8'hD1; #100;
A = 8'h1; B = 8'hD2; #100;
A = 8'h1; B = 8'hD3; #100;
A = 8'h1; B = 8'hD4; #100;
A = 8'h1; B = 8'hD5; #100;
A = 8'h1; B = 8'hD6; #100;
A = 8'h1; B = 8'hD7; #100;
A = 8'h1; B = 8'hD8; #100;
A = 8'h1; B = 8'hD9; #100;
A = 8'h1; B = 8'hDA; #100;
A = 8'h1; B = 8'hDB; #100;
A = 8'h1; B = 8'hDC; #100;
A = 8'h1; B = 8'hDD; #100;
A = 8'h1; B = 8'hDE; #100;
A = 8'h1; B = 8'hDF; #100;
A = 8'h1; B = 8'hE0; #100;
A = 8'h1; B = 8'hE1; #100;
A = 8'h1; B = 8'hE2; #100;
A = 8'h1; B = 8'hE3; #100;
A = 8'h1; B = 8'hE4; #100;
A = 8'h1; B = 8'hE5; #100;
A = 8'h1; B = 8'hE6; #100;
A = 8'h1; B = 8'hE7; #100;
A = 8'h1; B = 8'hE8; #100;
A = 8'h1; B = 8'hE9; #100;
A = 8'h1; B = 8'hEA; #100;
A = 8'h1; B = 8'hEB; #100;
A = 8'h1; B = 8'hEC; #100;
A = 8'h1; B = 8'hED; #100;
A = 8'h1; B = 8'hEE; #100;
A = 8'h1; B = 8'hEF; #100;
A = 8'h1; B = 8'hF0; #100;
A = 8'h1; B = 8'hF1; #100;
A = 8'h1; B = 8'hF2; #100;
A = 8'h1; B = 8'hF3; #100;
A = 8'h1; B = 8'hF4; #100;
A = 8'h1; B = 8'hF5; #100;
A = 8'h1; B = 8'hF6; #100;
A = 8'h1; B = 8'hF7; #100;
A = 8'h1; B = 8'hF8; #100;
A = 8'h1; B = 8'hF9; #100;
A = 8'h1; B = 8'hFA; #100;
A = 8'h1; B = 8'hFB; #100;
A = 8'h1; B = 8'hFC; #100;
A = 8'h1; B = 8'hFD; #100;
A = 8'h1; B = 8'hFE; #100;
A = 8'h1; B = 8'hFF; #100;
A = 8'h2; B = 8'h0; #100;
A = 8'h2; B = 8'h1; #100;
A = 8'h2; B = 8'h2; #100;
A = 8'h2; B = 8'h3; #100;
A = 8'h2; B = 8'h4; #100;
A = 8'h2; B = 8'h5; #100;
A = 8'h2; B = 8'h6; #100;
A = 8'h2; B = 8'h7; #100;
A = 8'h2; B = 8'h8; #100;
A = 8'h2; B = 8'h9; #100;
A = 8'h2; B = 8'hA; #100;
A = 8'h2; B = 8'hB; #100;
A = 8'h2; B = 8'hC; #100;
A = 8'h2; B = 8'hD; #100;
A = 8'h2; B = 8'hE; #100;
A = 8'h2; B = 8'hF; #100;
A = 8'h2; B = 8'h10; #100;
A = 8'h2; B = 8'h11; #100;
A = 8'h2; B = 8'h12; #100;
A = 8'h2; B = 8'h13; #100;
A = 8'h2; B = 8'h14; #100;
A = 8'h2; B = 8'h15; #100;
A = 8'h2; B = 8'h16; #100;
A = 8'h2; B = 8'h17; #100;
A = 8'h2; B = 8'h18; #100;
A = 8'h2; B = 8'h19; #100;
A = 8'h2; B = 8'h1A; #100;
A = 8'h2; B = 8'h1B; #100;
A = 8'h2; B = 8'h1C; #100;
A = 8'h2; B = 8'h1D; #100;
A = 8'h2; B = 8'h1E; #100;
A = 8'h2; B = 8'h1F; #100;
A = 8'h2; B = 8'h20; #100;
A = 8'h2; B = 8'h21; #100;
A = 8'h2; B = 8'h22; #100;
A = 8'h2; B = 8'h23; #100;
A = 8'h2; B = 8'h24; #100;
A = 8'h2; B = 8'h25; #100;
A = 8'h2; B = 8'h26; #100;
A = 8'h2; B = 8'h27; #100;
A = 8'h2; B = 8'h28; #100;
A = 8'h2; B = 8'h29; #100;
A = 8'h2; B = 8'h2A; #100;
A = 8'h2; B = 8'h2B; #100;
A = 8'h2; B = 8'h2C; #100;
A = 8'h2; B = 8'h2D; #100;
A = 8'h2; B = 8'h2E; #100;
A = 8'h2; B = 8'h2F; #100;
A = 8'h2; B = 8'h30; #100;
A = 8'h2; B = 8'h31; #100;
A = 8'h2; B = 8'h32; #100;
A = 8'h2; B = 8'h33; #100;
A = 8'h2; B = 8'h34; #100;
A = 8'h2; B = 8'h35; #100;
A = 8'h2; B = 8'h36; #100;
A = 8'h2; B = 8'h37; #100;
A = 8'h2; B = 8'h38; #100;
A = 8'h2; B = 8'h39; #100;
A = 8'h2; B = 8'h3A; #100;
A = 8'h2; B = 8'h3B; #100;
A = 8'h2; B = 8'h3C; #100;
A = 8'h2; B = 8'h3D; #100;
A = 8'h2; B = 8'h3E; #100;
A = 8'h2; B = 8'h3F; #100;
A = 8'h2; B = 8'h40; #100;
A = 8'h2; B = 8'h41; #100;
A = 8'h2; B = 8'h42; #100;
A = 8'h2; B = 8'h43; #100;
A = 8'h2; B = 8'h44; #100;
A = 8'h2; B = 8'h45; #100;
A = 8'h2; B = 8'h46; #100;
A = 8'h2; B = 8'h47; #100;
A = 8'h2; B = 8'h48; #100;
A = 8'h2; B = 8'h49; #100;
A = 8'h2; B = 8'h4A; #100;
A = 8'h2; B = 8'h4B; #100;
A = 8'h2; B = 8'h4C; #100;
A = 8'h2; B = 8'h4D; #100;
A = 8'h2; B = 8'h4E; #100;
A = 8'h2; B = 8'h4F; #100;
A = 8'h2; B = 8'h50; #100;
A = 8'h2; B = 8'h51; #100;
A = 8'h2; B = 8'h52; #100;
A = 8'h2; B = 8'h53; #100;
A = 8'h2; B = 8'h54; #100;
A = 8'h2; B = 8'h55; #100;
A = 8'h2; B = 8'h56; #100;
A = 8'h2; B = 8'h57; #100;
A = 8'h2; B = 8'h58; #100;
A = 8'h2; B = 8'h59; #100;
A = 8'h2; B = 8'h5A; #100;
A = 8'h2; B = 8'h5B; #100;
A = 8'h2; B = 8'h5C; #100;
A = 8'h2; B = 8'h5D; #100;
A = 8'h2; B = 8'h5E; #100;
A = 8'h2; B = 8'h5F; #100;
A = 8'h2; B = 8'h60; #100;
A = 8'h2; B = 8'h61; #100;
A = 8'h2; B = 8'h62; #100;
A = 8'h2; B = 8'h63; #100;
A = 8'h2; B = 8'h64; #100;
A = 8'h2; B = 8'h65; #100;
A = 8'h2; B = 8'h66; #100;
A = 8'h2; B = 8'h67; #100;
A = 8'h2; B = 8'h68; #100;
A = 8'h2; B = 8'h69; #100;
A = 8'h2; B = 8'h6A; #100;
A = 8'h2; B = 8'h6B; #100;
A = 8'h2; B = 8'h6C; #100;
A = 8'h2; B = 8'h6D; #100;
A = 8'h2; B = 8'h6E; #100;
A = 8'h2; B = 8'h6F; #100;
A = 8'h2; B = 8'h70; #100;
A = 8'h2; B = 8'h71; #100;
A = 8'h2; B = 8'h72; #100;
A = 8'h2; B = 8'h73; #100;
A = 8'h2; B = 8'h74; #100;
A = 8'h2; B = 8'h75; #100;
A = 8'h2; B = 8'h76; #100;
A = 8'h2; B = 8'h77; #100;
A = 8'h2; B = 8'h78; #100;
A = 8'h2; B = 8'h79; #100;
A = 8'h2; B = 8'h7A; #100;
A = 8'h2; B = 8'h7B; #100;
A = 8'h2; B = 8'h7C; #100;
A = 8'h2; B = 8'h7D; #100;
A = 8'h2; B = 8'h7E; #100;
A = 8'h2; B = 8'h7F; #100;
A = 8'h2; B = 8'h80; #100;
A = 8'h2; B = 8'h81; #100;
A = 8'h2; B = 8'h82; #100;
A = 8'h2; B = 8'h83; #100;
A = 8'h2; B = 8'h84; #100;
A = 8'h2; B = 8'h85; #100;
A = 8'h2; B = 8'h86; #100;
A = 8'h2; B = 8'h87; #100;
A = 8'h2; B = 8'h88; #100;
A = 8'h2; B = 8'h89; #100;
A = 8'h2; B = 8'h8A; #100;
A = 8'h2; B = 8'h8B; #100;
A = 8'h2; B = 8'h8C; #100;
A = 8'h2; B = 8'h8D; #100;
A = 8'h2; B = 8'h8E; #100;
A = 8'h2; B = 8'h8F; #100;
A = 8'h2; B = 8'h90; #100;
A = 8'h2; B = 8'h91; #100;
A = 8'h2; B = 8'h92; #100;
A = 8'h2; B = 8'h93; #100;
A = 8'h2; B = 8'h94; #100;
A = 8'h2; B = 8'h95; #100;
A = 8'h2; B = 8'h96; #100;
A = 8'h2; B = 8'h97; #100;
A = 8'h2; B = 8'h98; #100;
A = 8'h2; B = 8'h99; #100;
A = 8'h2; B = 8'h9A; #100;
A = 8'h2; B = 8'h9B; #100;
A = 8'h2; B = 8'h9C; #100;
A = 8'h2; B = 8'h9D; #100;
A = 8'h2; B = 8'h9E; #100;
A = 8'h2; B = 8'h9F; #100;
A = 8'h2; B = 8'hA0; #100;
A = 8'h2; B = 8'hA1; #100;
A = 8'h2; B = 8'hA2; #100;
A = 8'h2; B = 8'hA3; #100;
A = 8'h2; B = 8'hA4; #100;
A = 8'h2; B = 8'hA5; #100;
A = 8'h2; B = 8'hA6; #100;
A = 8'h2; B = 8'hA7; #100;
A = 8'h2; B = 8'hA8; #100;
A = 8'h2; B = 8'hA9; #100;
A = 8'h2; B = 8'hAA; #100;
A = 8'h2; B = 8'hAB; #100;
A = 8'h2; B = 8'hAC; #100;
A = 8'h2; B = 8'hAD; #100;
A = 8'h2; B = 8'hAE; #100;
A = 8'h2; B = 8'hAF; #100;
A = 8'h2; B = 8'hB0; #100;
A = 8'h2; B = 8'hB1; #100;
A = 8'h2; B = 8'hB2; #100;
A = 8'h2; B = 8'hB3; #100;
A = 8'h2; B = 8'hB4; #100;
A = 8'h2; B = 8'hB5; #100;
A = 8'h2; B = 8'hB6; #100;
A = 8'h2; B = 8'hB7; #100;
A = 8'h2; B = 8'hB8; #100;
A = 8'h2; B = 8'hB9; #100;
A = 8'h2; B = 8'hBA; #100;
A = 8'h2; B = 8'hBB; #100;
A = 8'h2; B = 8'hBC; #100;
A = 8'h2; B = 8'hBD; #100;
A = 8'h2; B = 8'hBE; #100;
A = 8'h2; B = 8'hBF; #100;
A = 8'h2; B = 8'hC0; #100;
A = 8'h2; B = 8'hC1; #100;
A = 8'h2; B = 8'hC2; #100;
A = 8'h2; B = 8'hC3; #100;
A = 8'h2; B = 8'hC4; #100;
A = 8'h2; B = 8'hC5; #100;
A = 8'h2; B = 8'hC6; #100;
A = 8'h2; B = 8'hC7; #100;
A = 8'h2; B = 8'hC8; #100;
A = 8'h2; B = 8'hC9; #100;
A = 8'h2; B = 8'hCA; #100;
A = 8'h2; B = 8'hCB; #100;
A = 8'h2; B = 8'hCC; #100;
A = 8'h2; B = 8'hCD; #100;
A = 8'h2; B = 8'hCE; #100;
A = 8'h2; B = 8'hCF; #100;
A = 8'h2; B = 8'hD0; #100;
A = 8'h2; B = 8'hD1; #100;
A = 8'h2; B = 8'hD2; #100;
A = 8'h2; B = 8'hD3; #100;
A = 8'h2; B = 8'hD4; #100;
A = 8'h2; B = 8'hD5; #100;
A = 8'h2; B = 8'hD6; #100;
A = 8'h2; B = 8'hD7; #100;
A = 8'h2; B = 8'hD8; #100;
A = 8'h2; B = 8'hD9; #100;
A = 8'h2; B = 8'hDA; #100;
A = 8'h2; B = 8'hDB; #100;
A = 8'h2; B = 8'hDC; #100;
A = 8'h2; B = 8'hDD; #100;
A = 8'h2; B = 8'hDE; #100;
A = 8'h2; B = 8'hDF; #100;
A = 8'h2; B = 8'hE0; #100;
A = 8'h2; B = 8'hE1; #100;
A = 8'h2; B = 8'hE2; #100;
A = 8'h2; B = 8'hE3; #100;
A = 8'h2; B = 8'hE4; #100;
A = 8'h2; B = 8'hE5; #100;
A = 8'h2; B = 8'hE6; #100;
A = 8'h2; B = 8'hE7; #100;
A = 8'h2; B = 8'hE8; #100;
A = 8'h2; B = 8'hE9; #100;
A = 8'h2; B = 8'hEA; #100;
A = 8'h2; B = 8'hEB; #100;
A = 8'h2; B = 8'hEC; #100;
A = 8'h2; B = 8'hED; #100;
A = 8'h2; B = 8'hEE; #100;
A = 8'h2; B = 8'hEF; #100;
A = 8'h2; B = 8'hF0; #100;
A = 8'h2; B = 8'hF1; #100;
A = 8'h2; B = 8'hF2; #100;
A = 8'h2; B = 8'hF3; #100;
A = 8'h2; B = 8'hF4; #100;
A = 8'h2; B = 8'hF5; #100;
A = 8'h2; B = 8'hF6; #100;
A = 8'h2; B = 8'hF7; #100;
A = 8'h2; B = 8'hF8; #100;
A = 8'h2; B = 8'hF9; #100;
A = 8'h2; B = 8'hFA; #100;
A = 8'h2; B = 8'hFB; #100;
A = 8'h2; B = 8'hFC; #100;
A = 8'h2; B = 8'hFD; #100;
A = 8'h2; B = 8'hFE; #100;
A = 8'h2; B = 8'hFF; #100;
A = 8'h3; B = 8'h0; #100;
A = 8'h3; B = 8'h1; #100;
A = 8'h3; B = 8'h2; #100;
A = 8'h3; B = 8'h3; #100;
A = 8'h3; B = 8'h4; #100;
A = 8'h3; B = 8'h5; #100;
A = 8'h3; B = 8'h6; #100;
A = 8'h3; B = 8'h7; #100;
A = 8'h3; B = 8'h8; #100;
A = 8'h3; B = 8'h9; #100;
A = 8'h3; B = 8'hA; #100;
A = 8'h3; B = 8'hB; #100;
A = 8'h3; B = 8'hC; #100;
A = 8'h3; B = 8'hD; #100;
A = 8'h3; B = 8'hE; #100;
A = 8'h3; B = 8'hF; #100;
A = 8'h3; B = 8'h10; #100;
A = 8'h3; B = 8'h11; #100;
A = 8'h3; B = 8'h12; #100;
A = 8'h3; B = 8'h13; #100;
A = 8'h3; B = 8'h14; #100;
A = 8'h3; B = 8'h15; #100;
A = 8'h3; B = 8'h16; #100;
A = 8'h3; B = 8'h17; #100;
A = 8'h3; B = 8'h18; #100;
A = 8'h3; B = 8'h19; #100;
A = 8'h3; B = 8'h1A; #100;
A = 8'h3; B = 8'h1B; #100;
A = 8'h3; B = 8'h1C; #100;
A = 8'h3; B = 8'h1D; #100;
A = 8'h3; B = 8'h1E; #100;
A = 8'h3; B = 8'h1F; #100;
A = 8'h3; B = 8'h20; #100;
A = 8'h3; B = 8'h21; #100;
A = 8'h3; B = 8'h22; #100;
A = 8'h3; B = 8'h23; #100;
A = 8'h3; B = 8'h24; #100;
A = 8'h3; B = 8'h25; #100;
A = 8'h3; B = 8'h26; #100;
A = 8'h3; B = 8'h27; #100;
A = 8'h3; B = 8'h28; #100;
A = 8'h3; B = 8'h29; #100;
A = 8'h3; B = 8'h2A; #100;
A = 8'h3; B = 8'h2B; #100;
A = 8'h3; B = 8'h2C; #100;
A = 8'h3; B = 8'h2D; #100;
A = 8'h3; B = 8'h2E; #100;
A = 8'h3; B = 8'h2F; #100;
A = 8'h3; B = 8'h30; #100;
A = 8'h3; B = 8'h31; #100;
A = 8'h3; B = 8'h32; #100;
A = 8'h3; B = 8'h33; #100;
A = 8'h3; B = 8'h34; #100;
A = 8'h3; B = 8'h35; #100;
A = 8'h3; B = 8'h36; #100;
A = 8'h3; B = 8'h37; #100;
A = 8'h3; B = 8'h38; #100;
A = 8'h3; B = 8'h39; #100;
A = 8'h3; B = 8'h3A; #100;
A = 8'h3; B = 8'h3B; #100;
A = 8'h3; B = 8'h3C; #100;
A = 8'h3; B = 8'h3D; #100;
A = 8'h3; B = 8'h3E; #100;
A = 8'h3; B = 8'h3F; #100;
A = 8'h3; B = 8'h40; #100;
A = 8'h3; B = 8'h41; #100;
A = 8'h3; B = 8'h42; #100;
A = 8'h3; B = 8'h43; #100;
A = 8'h3; B = 8'h44; #100;
A = 8'h3; B = 8'h45; #100;
A = 8'h3; B = 8'h46; #100;
A = 8'h3; B = 8'h47; #100;
A = 8'h3; B = 8'h48; #100;
A = 8'h3; B = 8'h49; #100;
A = 8'h3; B = 8'h4A; #100;
A = 8'h3; B = 8'h4B; #100;
A = 8'h3; B = 8'h4C; #100;
A = 8'h3; B = 8'h4D; #100;
A = 8'h3; B = 8'h4E; #100;
A = 8'h3; B = 8'h4F; #100;
A = 8'h3; B = 8'h50; #100;
A = 8'h3; B = 8'h51; #100;
A = 8'h3; B = 8'h52; #100;
A = 8'h3; B = 8'h53; #100;
A = 8'h3; B = 8'h54; #100;
A = 8'h3; B = 8'h55; #100;
A = 8'h3; B = 8'h56; #100;
A = 8'h3; B = 8'h57; #100;
A = 8'h3; B = 8'h58; #100;
A = 8'h3; B = 8'h59; #100;
A = 8'h3; B = 8'h5A; #100;
A = 8'h3; B = 8'h5B; #100;
A = 8'h3; B = 8'h5C; #100;
A = 8'h3; B = 8'h5D; #100;
A = 8'h3; B = 8'h5E; #100;
A = 8'h3; B = 8'h5F; #100;
A = 8'h3; B = 8'h60; #100;
A = 8'h3; B = 8'h61; #100;
A = 8'h3; B = 8'h62; #100;
A = 8'h3; B = 8'h63; #100;
A = 8'h3; B = 8'h64; #100;
A = 8'h3; B = 8'h65; #100;
A = 8'h3; B = 8'h66; #100;
A = 8'h3; B = 8'h67; #100;
A = 8'h3; B = 8'h68; #100;
A = 8'h3; B = 8'h69; #100;
A = 8'h3; B = 8'h6A; #100;
A = 8'h3; B = 8'h6B; #100;
A = 8'h3; B = 8'h6C; #100;
A = 8'h3; B = 8'h6D; #100;
A = 8'h3; B = 8'h6E; #100;
A = 8'h3; B = 8'h6F; #100;
A = 8'h3; B = 8'h70; #100;
A = 8'h3; B = 8'h71; #100;
A = 8'h3; B = 8'h72; #100;
A = 8'h3; B = 8'h73; #100;
A = 8'h3; B = 8'h74; #100;
A = 8'h3; B = 8'h75; #100;
A = 8'h3; B = 8'h76; #100;
A = 8'h3; B = 8'h77; #100;
A = 8'h3; B = 8'h78; #100;
A = 8'h3; B = 8'h79; #100;
A = 8'h3; B = 8'h7A; #100;
A = 8'h3; B = 8'h7B; #100;
A = 8'h3; B = 8'h7C; #100;
A = 8'h3; B = 8'h7D; #100;
A = 8'h3; B = 8'h7E; #100;
A = 8'h3; B = 8'h7F; #100;
A = 8'h3; B = 8'h80; #100;
A = 8'h3; B = 8'h81; #100;
A = 8'h3; B = 8'h82; #100;
A = 8'h3; B = 8'h83; #100;
A = 8'h3; B = 8'h84; #100;
A = 8'h3; B = 8'h85; #100;
A = 8'h3; B = 8'h86; #100;
A = 8'h3; B = 8'h87; #100;
A = 8'h3; B = 8'h88; #100;
A = 8'h3; B = 8'h89; #100;
A = 8'h3; B = 8'h8A; #100;
A = 8'h3; B = 8'h8B; #100;
A = 8'h3; B = 8'h8C; #100;
A = 8'h3; B = 8'h8D; #100;
A = 8'h3; B = 8'h8E; #100;
A = 8'h3; B = 8'h8F; #100;
A = 8'h3; B = 8'h90; #100;
A = 8'h3; B = 8'h91; #100;
A = 8'h3; B = 8'h92; #100;
A = 8'h3; B = 8'h93; #100;
A = 8'h3; B = 8'h94; #100;
A = 8'h3; B = 8'h95; #100;
A = 8'h3; B = 8'h96; #100;
A = 8'h3; B = 8'h97; #100;
A = 8'h3; B = 8'h98; #100;
A = 8'h3; B = 8'h99; #100;
A = 8'h3; B = 8'h9A; #100;
A = 8'h3; B = 8'h9B; #100;
A = 8'h3; B = 8'h9C; #100;
A = 8'h3; B = 8'h9D; #100;
A = 8'h3; B = 8'h9E; #100;
A = 8'h3; B = 8'h9F; #100;
A = 8'h3; B = 8'hA0; #100;
A = 8'h3; B = 8'hA1; #100;
A = 8'h3; B = 8'hA2; #100;
A = 8'h3; B = 8'hA3; #100;
A = 8'h3; B = 8'hA4; #100;
A = 8'h3; B = 8'hA5; #100;
A = 8'h3; B = 8'hA6; #100;
A = 8'h3; B = 8'hA7; #100;
A = 8'h3; B = 8'hA8; #100;
A = 8'h3; B = 8'hA9; #100;
A = 8'h3; B = 8'hAA; #100;
A = 8'h3; B = 8'hAB; #100;
A = 8'h3; B = 8'hAC; #100;
A = 8'h3; B = 8'hAD; #100;
A = 8'h3; B = 8'hAE; #100;
A = 8'h3; B = 8'hAF; #100;
A = 8'h3; B = 8'hB0; #100;
A = 8'h3; B = 8'hB1; #100;
A = 8'h3; B = 8'hB2; #100;
A = 8'h3; B = 8'hB3; #100;
A = 8'h3; B = 8'hB4; #100;
A = 8'h3; B = 8'hB5; #100;
A = 8'h3; B = 8'hB6; #100;
A = 8'h3; B = 8'hB7; #100;
A = 8'h3; B = 8'hB8; #100;
A = 8'h3; B = 8'hB9; #100;
A = 8'h3; B = 8'hBA; #100;
A = 8'h3; B = 8'hBB; #100;
A = 8'h3; B = 8'hBC; #100;
A = 8'h3; B = 8'hBD; #100;
A = 8'h3; B = 8'hBE; #100;
A = 8'h3; B = 8'hBF; #100;
A = 8'h3; B = 8'hC0; #100;
A = 8'h3; B = 8'hC1; #100;
A = 8'h3; B = 8'hC2; #100;
A = 8'h3; B = 8'hC3; #100;
A = 8'h3; B = 8'hC4; #100;
A = 8'h3; B = 8'hC5; #100;
A = 8'h3; B = 8'hC6; #100;
A = 8'h3; B = 8'hC7; #100;
A = 8'h3; B = 8'hC8; #100;
A = 8'h3; B = 8'hC9; #100;
A = 8'h3; B = 8'hCA; #100;
A = 8'h3; B = 8'hCB; #100;
A = 8'h3; B = 8'hCC; #100;
A = 8'h3; B = 8'hCD; #100;
A = 8'h3; B = 8'hCE; #100;
A = 8'h3; B = 8'hCF; #100;
A = 8'h3; B = 8'hD0; #100;
A = 8'h3; B = 8'hD1; #100;
A = 8'h3; B = 8'hD2; #100;
A = 8'h3; B = 8'hD3; #100;
A = 8'h3; B = 8'hD4; #100;
A = 8'h3; B = 8'hD5; #100;
A = 8'h3; B = 8'hD6; #100;
A = 8'h3; B = 8'hD7; #100;
A = 8'h3; B = 8'hD8; #100;
A = 8'h3; B = 8'hD9; #100;
A = 8'h3; B = 8'hDA; #100;
A = 8'h3; B = 8'hDB; #100;
A = 8'h3; B = 8'hDC; #100;
A = 8'h3; B = 8'hDD; #100;
A = 8'h3; B = 8'hDE; #100;
A = 8'h3; B = 8'hDF; #100;
A = 8'h3; B = 8'hE0; #100;
A = 8'h3; B = 8'hE1; #100;
A = 8'h3; B = 8'hE2; #100;
A = 8'h3; B = 8'hE3; #100;
A = 8'h3; B = 8'hE4; #100;
A = 8'h3; B = 8'hE5; #100;
A = 8'h3; B = 8'hE6; #100;
A = 8'h3; B = 8'hE7; #100;
A = 8'h3; B = 8'hE8; #100;
A = 8'h3; B = 8'hE9; #100;
A = 8'h3; B = 8'hEA; #100;
A = 8'h3; B = 8'hEB; #100;
A = 8'h3; B = 8'hEC; #100;
A = 8'h3; B = 8'hED; #100;
A = 8'h3; B = 8'hEE; #100;
A = 8'h3; B = 8'hEF; #100;
A = 8'h3; B = 8'hF0; #100;
A = 8'h3; B = 8'hF1; #100;
A = 8'h3; B = 8'hF2; #100;
A = 8'h3; B = 8'hF3; #100;
A = 8'h3; B = 8'hF4; #100;
A = 8'h3; B = 8'hF5; #100;
A = 8'h3; B = 8'hF6; #100;
A = 8'h3; B = 8'hF7; #100;
A = 8'h3; B = 8'hF8; #100;
A = 8'h3; B = 8'hF9; #100;
A = 8'h3; B = 8'hFA; #100;
A = 8'h3; B = 8'hFB; #100;
A = 8'h3; B = 8'hFC; #100;
A = 8'h3; B = 8'hFD; #100;
A = 8'h3; B = 8'hFE; #100;
A = 8'h3; B = 8'hFF; #100;
A = 8'h4; B = 8'h0; #100;
A = 8'h4; B = 8'h1; #100;
A = 8'h4; B = 8'h2; #100;
A = 8'h4; B = 8'h3; #100;
A = 8'h4; B = 8'h4; #100;
A = 8'h4; B = 8'h5; #100;
A = 8'h4; B = 8'h6; #100;
A = 8'h4; B = 8'h7; #100;
A = 8'h4; B = 8'h8; #100;
A = 8'h4; B = 8'h9; #100;
A = 8'h4; B = 8'hA; #100;
A = 8'h4; B = 8'hB; #100;
A = 8'h4; B = 8'hC; #100;
A = 8'h4; B = 8'hD; #100;
A = 8'h4; B = 8'hE; #100;
A = 8'h4; B = 8'hF; #100;
A = 8'h4; B = 8'h10; #100;
A = 8'h4; B = 8'h11; #100;
A = 8'h4; B = 8'h12; #100;
A = 8'h4; B = 8'h13; #100;
A = 8'h4; B = 8'h14; #100;
A = 8'h4; B = 8'h15; #100;
A = 8'h4; B = 8'h16; #100;
A = 8'h4; B = 8'h17; #100;
A = 8'h4; B = 8'h18; #100;
A = 8'h4; B = 8'h19; #100;
A = 8'h4; B = 8'h1A; #100;
A = 8'h4; B = 8'h1B; #100;
A = 8'h4; B = 8'h1C; #100;
A = 8'h4; B = 8'h1D; #100;
A = 8'h4; B = 8'h1E; #100;
A = 8'h4; B = 8'h1F; #100;
A = 8'h4; B = 8'h20; #100;
A = 8'h4; B = 8'h21; #100;
A = 8'h4; B = 8'h22; #100;
A = 8'h4; B = 8'h23; #100;
A = 8'h4; B = 8'h24; #100;
A = 8'h4; B = 8'h25; #100;
A = 8'h4; B = 8'h26; #100;
A = 8'h4; B = 8'h27; #100;
A = 8'h4; B = 8'h28; #100;
A = 8'h4; B = 8'h29; #100;
A = 8'h4; B = 8'h2A; #100;
A = 8'h4; B = 8'h2B; #100;
A = 8'h4; B = 8'h2C; #100;
A = 8'h4; B = 8'h2D; #100;
A = 8'h4; B = 8'h2E; #100;
A = 8'h4; B = 8'h2F; #100;
A = 8'h4; B = 8'h30; #100;
A = 8'h4; B = 8'h31; #100;
A = 8'h4; B = 8'h32; #100;
A = 8'h4; B = 8'h33; #100;
A = 8'h4; B = 8'h34; #100;
A = 8'h4; B = 8'h35; #100;
A = 8'h4; B = 8'h36; #100;
A = 8'h4; B = 8'h37; #100;
A = 8'h4; B = 8'h38; #100;
A = 8'h4; B = 8'h39; #100;
A = 8'h4; B = 8'h3A; #100;
A = 8'h4; B = 8'h3B; #100;
A = 8'h4; B = 8'h3C; #100;
A = 8'h4; B = 8'h3D; #100;
A = 8'h4; B = 8'h3E; #100;
A = 8'h4; B = 8'h3F; #100;
A = 8'h4; B = 8'h40; #100;
A = 8'h4; B = 8'h41; #100;
A = 8'h4; B = 8'h42; #100;
A = 8'h4; B = 8'h43; #100;
A = 8'h4; B = 8'h44; #100;
A = 8'h4; B = 8'h45; #100;
A = 8'h4; B = 8'h46; #100;
A = 8'h4; B = 8'h47; #100;
A = 8'h4; B = 8'h48; #100;
A = 8'h4; B = 8'h49; #100;
A = 8'h4; B = 8'h4A; #100;
A = 8'h4; B = 8'h4B; #100;
A = 8'h4; B = 8'h4C; #100;
A = 8'h4; B = 8'h4D; #100;
A = 8'h4; B = 8'h4E; #100;
A = 8'h4; B = 8'h4F; #100;
A = 8'h4; B = 8'h50; #100;
A = 8'h4; B = 8'h51; #100;
A = 8'h4; B = 8'h52; #100;
A = 8'h4; B = 8'h53; #100;
A = 8'h4; B = 8'h54; #100;
A = 8'h4; B = 8'h55; #100;
A = 8'h4; B = 8'h56; #100;
A = 8'h4; B = 8'h57; #100;
A = 8'h4; B = 8'h58; #100;
A = 8'h4; B = 8'h59; #100;
A = 8'h4; B = 8'h5A; #100;
A = 8'h4; B = 8'h5B; #100;
A = 8'h4; B = 8'h5C; #100;
A = 8'h4; B = 8'h5D; #100;
A = 8'h4; B = 8'h5E; #100;
A = 8'h4; B = 8'h5F; #100;
A = 8'h4; B = 8'h60; #100;
A = 8'h4; B = 8'h61; #100;
A = 8'h4; B = 8'h62; #100;
A = 8'h4; B = 8'h63; #100;
A = 8'h4; B = 8'h64; #100;
A = 8'h4; B = 8'h65; #100;
A = 8'h4; B = 8'h66; #100;
A = 8'h4; B = 8'h67; #100;
A = 8'h4; B = 8'h68; #100;
A = 8'h4; B = 8'h69; #100;
A = 8'h4; B = 8'h6A; #100;
A = 8'h4; B = 8'h6B; #100;
A = 8'h4; B = 8'h6C; #100;
A = 8'h4; B = 8'h6D; #100;
A = 8'h4; B = 8'h6E; #100;
A = 8'h4; B = 8'h6F; #100;
A = 8'h4; B = 8'h70; #100;
A = 8'h4; B = 8'h71; #100;
A = 8'h4; B = 8'h72; #100;
A = 8'h4; B = 8'h73; #100;
A = 8'h4; B = 8'h74; #100;
A = 8'h4; B = 8'h75; #100;
A = 8'h4; B = 8'h76; #100;
A = 8'h4; B = 8'h77; #100;
A = 8'h4; B = 8'h78; #100;
A = 8'h4; B = 8'h79; #100;
A = 8'h4; B = 8'h7A; #100;
A = 8'h4; B = 8'h7B; #100;
A = 8'h4; B = 8'h7C; #100;
A = 8'h4; B = 8'h7D; #100;
A = 8'h4; B = 8'h7E; #100;
A = 8'h4; B = 8'h7F; #100;
A = 8'h4; B = 8'h80; #100;
A = 8'h4; B = 8'h81; #100;
A = 8'h4; B = 8'h82; #100;
A = 8'h4; B = 8'h83; #100;
A = 8'h4; B = 8'h84; #100;
A = 8'h4; B = 8'h85; #100;
A = 8'h4; B = 8'h86; #100;
A = 8'h4; B = 8'h87; #100;
A = 8'h4; B = 8'h88; #100;
A = 8'h4; B = 8'h89; #100;
A = 8'h4; B = 8'h8A; #100;
A = 8'h4; B = 8'h8B; #100;
A = 8'h4; B = 8'h8C; #100;
A = 8'h4; B = 8'h8D; #100;
A = 8'h4; B = 8'h8E; #100;
A = 8'h4; B = 8'h8F; #100;
A = 8'h4; B = 8'h90; #100;
A = 8'h4; B = 8'h91; #100;
A = 8'h4; B = 8'h92; #100;
A = 8'h4; B = 8'h93; #100;
A = 8'h4; B = 8'h94; #100;
A = 8'h4; B = 8'h95; #100;
A = 8'h4; B = 8'h96; #100;
A = 8'h4; B = 8'h97; #100;
A = 8'h4; B = 8'h98; #100;
A = 8'h4; B = 8'h99; #100;
A = 8'h4; B = 8'h9A; #100;
A = 8'h4; B = 8'h9B; #100;
A = 8'h4; B = 8'h9C; #100;
A = 8'h4; B = 8'h9D; #100;
A = 8'h4; B = 8'h9E; #100;
A = 8'h4; B = 8'h9F; #100;
A = 8'h4; B = 8'hA0; #100;
A = 8'h4; B = 8'hA1; #100;
A = 8'h4; B = 8'hA2; #100;
A = 8'h4; B = 8'hA3; #100;
A = 8'h4; B = 8'hA4; #100;
A = 8'h4; B = 8'hA5; #100;
A = 8'h4; B = 8'hA6; #100;
A = 8'h4; B = 8'hA7; #100;
A = 8'h4; B = 8'hA8; #100;
A = 8'h4; B = 8'hA9; #100;
A = 8'h4; B = 8'hAA; #100;
A = 8'h4; B = 8'hAB; #100;
A = 8'h4; B = 8'hAC; #100;
A = 8'h4; B = 8'hAD; #100;
A = 8'h4; B = 8'hAE; #100;
A = 8'h4; B = 8'hAF; #100;
A = 8'h4; B = 8'hB0; #100;
A = 8'h4; B = 8'hB1; #100;
A = 8'h4; B = 8'hB2; #100;
A = 8'h4; B = 8'hB3; #100;
A = 8'h4; B = 8'hB4; #100;
A = 8'h4; B = 8'hB5; #100;
A = 8'h4; B = 8'hB6; #100;
A = 8'h4; B = 8'hB7; #100;
A = 8'h4; B = 8'hB8; #100;
A = 8'h4; B = 8'hB9; #100;
A = 8'h4; B = 8'hBA; #100;
A = 8'h4; B = 8'hBB; #100;
A = 8'h4; B = 8'hBC; #100;
A = 8'h4; B = 8'hBD; #100;
A = 8'h4; B = 8'hBE; #100;
A = 8'h4; B = 8'hBF; #100;
A = 8'h4; B = 8'hC0; #100;
A = 8'h4; B = 8'hC1; #100;
A = 8'h4; B = 8'hC2; #100;
A = 8'h4; B = 8'hC3; #100;
A = 8'h4; B = 8'hC4; #100;
A = 8'h4; B = 8'hC5; #100;
A = 8'h4; B = 8'hC6; #100;
A = 8'h4; B = 8'hC7; #100;
A = 8'h4; B = 8'hC8; #100;
A = 8'h4; B = 8'hC9; #100;
A = 8'h4; B = 8'hCA; #100;
A = 8'h4; B = 8'hCB; #100;
A = 8'h4; B = 8'hCC; #100;
A = 8'h4; B = 8'hCD; #100;
A = 8'h4; B = 8'hCE; #100;
A = 8'h4; B = 8'hCF; #100;
A = 8'h4; B = 8'hD0; #100;
A = 8'h4; B = 8'hD1; #100;
A = 8'h4; B = 8'hD2; #100;
A = 8'h4; B = 8'hD3; #100;
A = 8'h4; B = 8'hD4; #100;
A = 8'h4; B = 8'hD5; #100;
A = 8'h4; B = 8'hD6; #100;
A = 8'h4; B = 8'hD7; #100;
A = 8'h4; B = 8'hD8; #100;
A = 8'h4; B = 8'hD9; #100;
A = 8'h4; B = 8'hDA; #100;
A = 8'h4; B = 8'hDB; #100;
A = 8'h4; B = 8'hDC; #100;
A = 8'h4; B = 8'hDD; #100;
A = 8'h4; B = 8'hDE; #100;
A = 8'h4; B = 8'hDF; #100;
A = 8'h4; B = 8'hE0; #100;
A = 8'h4; B = 8'hE1; #100;
A = 8'h4; B = 8'hE2; #100;
A = 8'h4; B = 8'hE3; #100;
A = 8'h4; B = 8'hE4; #100;
A = 8'h4; B = 8'hE5; #100;
A = 8'h4; B = 8'hE6; #100;
A = 8'h4; B = 8'hE7; #100;
A = 8'h4; B = 8'hE8; #100;
A = 8'h4; B = 8'hE9; #100;
A = 8'h4; B = 8'hEA; #100;
A = 8'h4; B = 8'hEB; #100;
A = 8'h4; B = 8'hEC; #100;
A = 8'h4; B = 8'hED; #100;
A = 8'h4; B = 8'hEE; #100;
A = 8'h4; B = 8'hEF; #100;
A = 8'h4; B = 8'hF0; #100;
A = 8'h4; B = 8'hF1; #100;
A = 8'h4; B = 8'hF2; #100;
A = 8'h4; B = 8'hF3; #100;
A = 8'h4; B = 8'hF4; #100;
A = 8'h4; B = 8'hF5; #100;
A = 8'h4; B = 8'hF6; #100;
A = 8'h4; B = 8'hF7; #100;
A = 8'h4; B = 8'hF8; #100;
A = 8'h4; B = 8'hF9; #100;
A = 8'h4; B = 8'hFA; #100;
A = 8'h4; B = 8'hFB; #100;
A = 8'h4; B = 8'hFC; #100;
A = 8'h4; B = 8'hFD; #100;
A = 8'h4; B = 8'hFE; #100;
A = 8'h4; B = 8'hFF; #100;
A = 8'h5; B = 8'h0; #100;
A = 8'h5; B = 8'h1; #100;
A = 8'h5; B = 8'h2; #100;
A = 8'h5; B = 8'h3; #100;
A = 8'h5; B = 8'h4; #100;
A = 8'h5; B = 8'h5; #100;
A = 8'h5; B = 8'h6; #100;
A = 8'h5; B = 8'h7; #100;
A = 8'h5; B = 8'h8; #100;
A = 8'h5; B = 8'h9; #100;
A = 8'h5; B = 8'hA; #100;
A = 8'h5; B = 8'hB; #100;
A = 8'h5; B = 8'hC; #100;
A = 8'h5; B = 8'hD; #100;
A = 8'h5; B = 8'hE; #100;
A = 8'h5; B = 8'hF; #100;
A = 8'h5; B = 8'h10; #100;
A = 8'h5; B = 8'h11; #100;
A = 8'h5; B = 8'h12; #100;
A = 8'h5; B = 8'h13; #100;
A = 8'h5; B = 8'h14; #100;
A = 8'h5; B = 8'h15; #100;
A = 8'h5; B = 8'h16; #100;
A = 8'h5; B = 8'h17; #100;
A = 8'h5; B = 8'h18; #100;
A = 8'h5; B = 8'h19; #100;
A = 8'h5; B = 8'h1A; #100;
A = 8'h5; B = 8'h1B; #100;
A = 8'h5; B = 8'h1C; #100;
A = 8'h5; B = 8'h1D; #100;
A = 8'h5; B = 8'h1E; #100;
A = 8'h5; B = 8'h1F; #100;
A = 8'h5; B = 8'h20; #100;
A = 8'h5; B = 8'h21; #100;
A = 8'h5; B = 8'h22; #100;
A = 8'h5; B = 8'h23; #100;
A = 8'h5; B = 8'h24; #100;
A = 8'h5; B = 8'h25; #100;
A = 8'h5; B = 8'h26; #100;
A = 8'h5; B = 8'h27; #100;
A = 8'h5; B = 8'h28; #100;
A = 8'h5; B = 8'h29; #100;
A = 8'h5; B = 8'h2A; #100;
A = 8'h5; B = 8'h2B; #100;
A = 8'h5; B = 8'h2C; #100;
A = 8'h5; B = 8'h2D; #100;
A = 8'h5; B = 8'h2E; #100;
A = 8'h5; B = 8'h2F; #100;
A = 8'h5; B = 8'h30; #100;
A = 8'h5; B = 8'h31; #100;
A = 8'h5; B = 8'h32; #100;
A = 8'h5; B = 8'h33; #100;
A = 8'h5; B = 8'h34; #100;
A = 8'h5; B = 8'h35; #100;
A = 8'h5; B = 8'h36; #100;
A = 8'h5; B = 8'h37; #100;
A = 8'h5; B = 8'h38; #100;
A = 8'h5; B = 8'h39; #100;
A = 8'h5; B = 8'h3A; #100;
A = 8'h5; B = 8'h3B; #100;
A = 8'h5; B = 8'h3C; #100;
A = 8'h5; B = 8'h3D; #100;
A = 8'h5; B = 8'h3E; #100;
A = 8'h5; B = 8'h3F; #100;
A = 8'h5; B = 8'h40; #100;
A = 8'h5; B = 8'h41; #100;
A = 8'h5; B = 8'h42; #100;
A = 8'h5; B = 8'h43; #100;
A = 8'h5; B = 8'h44; #100;
A = 8'h5; B = 8'h45; #100;
A = 8'h5; B = 8'h46; #100;
A = 8'h5; B = 8'h47; #100;
A = 8'h5; B = 8'h48; #100;
A = 8'h5; B = 8'h49; #100;
A = 8'h5; B = 8'h4A; #100;
A = 8'h5; B = 8'h4B; #100;
A = 8'h5; B = 8'h4C; #100;
A = 8'h5; B = 8'h4D; #100;
A = 8'h5; B = 8'h4E; #100;
A = 8'h5; B = 8'h4F; #100;
A = 8'h5; B = 8'h50; #100;
A = 8'h5; B = 8'h51; #100;
A = 8'h5; B = 8'h52; #100;
A = 8'h5; B = 8'h53; #100;
A = 8'h5; B = 8'h54; #100;
A = 8'h5; B = 8'h55; #100;
A = 8'h5; B = 8'h56; #100;
A = 8'h5; B = 8'h57; #100;
A = 8'h5; B = 8'h58; #100;
A = 8'h5; B = 8'h59; #100;
A = 8'h5; B = 8'h5A; #100;
A = 8'h5; B = 8'h5B; #100;
A = 8'h5; B = 8'h5C; #100;
A = 8'h5; B = 8'h5D; #100;
A = 8'h5; B = 8'h5E; #100;
A = 8'h5; B = 8'h5F; #100;
A = 8'h5; B = 8'h60; #100;
A = 8'h5; B = 8'h61; #100;
A = 8'h5; B = 8'h62; #100;
A = 8'h5; B = 8'h63; #100;
A = 8'h5; B = 8'h64; #100;
A = 8'h5; B = 8'h65; #100;
A = 8'h5; B = 8'h66; #100;
A = 8'h5; B = 8'h67; #100;
A = 8'h5; B = 8'h68; #100;
A = 8'h5; B = 8'h69; #100;
A = 8'h5; B = 8'h6A; #100;
A = 8'h5; B = 8'h6B; #100;
A = 8'h5; B = 8'h6C; #100;
A = 8'h5; B = 8'h6D; #100;
A = 8'h5; B = 8'h6E; #100;
A = 8'h5; B = 8'h6F; #100;
A = 8'h5; B = 8'h70; #100;
A = 8'h5; B = 8'h71; #100;
A = 8'h5; B = 8'h72; #100;
A = 8'h5; B = 8'h73; #100;
A = 8'h5; B = 8'h74; #100;
A = 8'h5; B = 8'h75; #100;
A = 8'h5; B = 8'h76; #100;
A = 8'h5; B = 8'h77; #100;
A = 8'h5; B = 8'h78; #100;
A = 8'h5; B = 8'h79; #100;
A = 8'h5; B = 8'h7A; #100;
A = 8'h5; B = 8'h7B; #100;
A = 8'h5; B = 8'h7C; #100;
A = 8'h5; B = 8'h7D; #100;
A = 8'h5; B = 8'h7E; #100;
A = 8'h5; B = 8'h7F; #100;
A = 8'h5; B = 8'h80; #100;
A = 8'h5; B = 8'h81; #100;
A = 8'h5; B = 8'h82; #100;
A = 8'h5; B = 8'h83; #100;
A = 8'h5; B = 8'h84; #100;
A = 8'h5; B = 8'h85; #100;
A = 8'h5; B = 8'h86; #100;
A = 8'h5; B = 8'h87; #100;
A = 8'h5; B = 8'h88; #100;
A = 8'h5; B = 8'h89; #100;
A = 8'h5; B = 8'h8A; #100;
A = 8'h5; B = 8'h8B; #100;
A = 8'h5; B = 8'h8C; #100;
A = 8'h5; B = 8'h8D; #100;
A = 8'h5; B = 8'h8E; #100;
A = 8'h5; B = 8'h8F; #100;
A = 8'h5; B = 8'h90; #100;
A = 8'h5; B = 8'h91; #100;
A = 8'h5; B = 8'h92; #100;
A = 8'h5; B = 8'h93; #100;
A = 8'h5; B = 8'h94; #100;
A = 8'h5; B = 8'h95; #100;
A = 8'h5; B = 8'h96; #100;
A = 8'h5; B = 8'h97; #100;
A = 8'h5; B = 8'h98; #100;
A = 8'h5; B = 8'h99; #100;
A = 8'h5; B = 8'h9A; #100;
A = 8'h5; B = 8'h9B; #100;
A = 8'h5; B = 8'h9C; #100;
A = 8'h5; B = 8'h9D; #100;
A = 8'h5; B = 8'h9E; #100;
A = 8'h5; B = 8'h9F; #100;
A = 8'h5; B = 8'hA0; #100;
A = 8'h5; B = 8'hA1; #100;
A = 8'h5; B = 8'hA2; #100;
A = 8'h5; B = 8'hA3; #100;
A = 8'h5; B = 8'hA4; #100;
A = 8'h5; B = 8'hA5; #100;
A = 8'h5; B = 8'hA6; #100;
A = 8'h5; B = 8'hA7; #100;
A = 8'h5; B = 8'hA8; #100;
A = 8'h5; B = 8'hA9; #100;
A = 8'h5; B = 8'hAA; #100;
A = 8'h5; B = 8'hAB; #100;
A = 8'h5; B = 8'hAC; #100;
A = 8'h5; B = 8'hAD; #100;
A = 8'h5; B = 8'hAE; #100;
A = 8'h5; B = 8'hAF; #100;
A = 8'h5; B = 8'hB0; #100;
A = 8'h5; B = 8'hB1; #100;
A = 8'h5; B = 8'hB2; #100;
A = 8'h5; B = 8'hB3; #100;
A = 8'h5; B = 8'hB4; #100;
A = 8'h5; B = 8'hB5; #100;
A = 8'h5; B = 8'hB6; #100;
A = 8'h5; B = 8'hB7; #100;
A = 8'h5; B = 8'hB8; #100;
A = 8'h5; B = 8'hB9; #100;
A = 8'h5; B = 8'hBA; #100;
A = 8'h5; B = 8'hBB; #100;
A = 8'h5; B = 8'hBC; #100;
A = 8'h5; B = 8'hBD; #100;
A = 8'h5; B = 8'hBE; #100;
A = 8'h5; B = 8'hBF; #100;
A = 8'h5; B = 8'hC0; #100;
A = 8'h5; B = 8'hC1; #100;
A = 8'h5; B = 8'hC2; #100;
A = 8'h5; B = 8'hC3; #100;
A = 8'h5; B = 8'hC4; #100;
A = 8'h5; B = 8'hC5; #100;
A = 8'h5; B = 8'hC6; #100;
A = 8'h5; B = 8'hC7; #100;
A = 8'h5; B = 8'hC8; #100;
A = 8'h5; B = 8'hC9; #100;
A = 8'h5; B = 8'hCA; #100;
A = 8'h5; B = 8'hCB; #100;
A = 8'h5; B = 8'hCC; #100;
A = 8'h5; B = 8'hCD; #100;
A = 8'h5; B = 8'hCE; #100;
A = 8'h5; B = 8'hCF; #100;
A = 8'h5; B = 8'hD0; #100;
A = 8'h5; B = 8'hD1; #100;
A = 8'h5; B = 8'hD2; #100;
A = 8'h5; B = 8'hD3; #100;
A = 8'h5; B = 8'hD4; #100;
A = 8'h5; B = 8'hD5; #100;
A = 8'h5; B = 8'hD6; #100;
A = 8'h5; B = 8'hD7; #100;
A = 8'h5; B = 8'hD8; #100;
A = 8'h5; B = 8'hD9; #100;
A = 8'h5; B = 8'hDA; #100;
A = 8'h5; B = 8'hDB; #100;
A = 8'h5; B = 8'hDC; #100;
A = 8'h5; B = 8'hDD; #100;
A = 8'h5; B = 8'hDE; #100;
A = 8'h5; B = 8'hDF; #100;
A = 8'h5; B = 8'hE0; #100;
A = 8'h5; B = 8'hE1; #100;
A = 8'h5; B = 8'hE2; #100;
A = 8'h5; B = 8'hE3; #100;
A = 8'h5; B = 8'hE4; #100;
A = 8'h5; B = 8'hE5; #100;
A = 8'h5; B = 8'hE6; #100;
A = 8'h5; B = 8'hE7; #100;
A = 8'h5; B = 8'hE8; #100;
A = 8'h5; B = 8'hE9; #100;
A = 8'h5; B = 8'hEA; #100;
A = 8'h5; B = 8'hEB; #100;
A = 8'h5; B = 8'hEC; #100;
A = 8'h5; B = 8'hED; #100;
A = 8'h5; B = 8'hEE; #100;
A = 8'h5; B = 8'hEF; #100;
A = 8'h5; B = 8'hF0; #100;
A = 8'h5; B = 8'hF1; #100;
A = 8'h5; B = 8'hF2; #100;
A = 8'h5; B = 8'hF3; #100;
A = 8'h5; B = 8'hF4; #100;
A = 8'h5; B = 8'hF5; #100;
A = 8'h5; B = 8'hF6; #100;
A = 8'h5; B = 8'hF7; #100;
A = 8'h5; B = 8'hF8; #100;
A = 8'h5; B = 8'hF9; #100;
A = 8'h5; B = 8'hFA; #100;
A = 8'h5; B = 8'hFB; #100;
A = 8'h5; B = 8'hFC; #100;
A = 8'h5; B = 8'hFD; #100;
A = 8'h5; B = 8'hFE; #100;
A = 8'h5; B = 8'hFF; #100;
A = 8'h6; B = 8'h0; #100;
A = 8'h6; B = 8'h1; #100;
A = 8'h6; B = 8'h2; #100;
A = 8'h6; B = 8'h3; #100;
A = 8'h6; B = 8'h4; #100;
A = 8'h6; B = 8'h5; #100;
A = 8'h6; B = 8'h6; #100;
A = 8'h6; B = 8'h7; #100;
A = 8'h6; B = 8'h8; #100;
A = 8'h6; B = 8'h9; #100;
A = 8'h6; B = 8'hA; #100;
A = 8'h6; B = 8'hB; #100;
A = 8'h6; B = 8'hC; #100;
A = 8'h6; B = 8'hD; #100;
A = 8'h6; B = 8'hE; #100;
A = 8'h6; B = 8'hF; #100;
A = 8'h6; B = 8'h10; #100;
A = 8'h6; B = 8'h11; #100;
A = 8'h6; B = 8'h12; #100;
A = 8'h6; B = 8'h13; #100;
A = 8'h6; B = 8'h14; #100;
A = 8'h6; B = 8'h15; #100;
A = 8'h6; B = 8'h16; #100;
A = 8'h6; B = 8'h17; #100;
A = 8'h6; B = 8'h18; #100;
A = 8'h6; B = 8'h19; #100;
A = 8'h6; B = 8'h1A; #100;
A = 8'h6; B = 8'h1B; #100;
A = 8'h6; B = 8'h1C; #100;
A = 8'h6; B = 8'h1D; #100;
A = 8'h6; B = 8'h1E; #100;
A = 8'h6; B = 8'h1F; #100;
A = 8'h6; B = 8'h20; #100;
A = 8'h6; B = 8'h21; #100;
A = 8'h6; B = 8'h22; #100;
A = 8'h6; B = 8'h23; #100;
A = 8'h6; B = 8'h24; #100;
A = 8'h6; B = 8'h25; #100;
A = 8'h6; B = 8'h26; #100;
A = 8'h6; B = 8'h27; #100;
A = 8'h6; B = 8'h28; #100;
A = 8'h6; B = 8'h29; #100;
A = 8'h6; B = 8'h2A; #100;
A = 8'h6; B = 8'h2B; #100;
A = 8'h6; B = 8'h2C; #100;
A = 8'h6; B = 8'h2D; #100;
A = 8'h6; B = 8'h2E; #100;
A = 8'h6; B = 8'h2F; #100;
A = 8'h6; B = 8'h30; #100;
A = 8'h6; B = 8'h31; #100;
A = 8'h6; B = 8'h32; #100;
A = 8'h6; B = 8'h33; #100;
A = 8'h6; B = 8'h34; #100;
A = 8'h6; B = 8'h35; #100;
A = 8'h6; B = 8'h36; #100;
A = 8'h6; B = 8'h37; #100;
A = 8'h6; B = 8'h38; #100;
A = 8'h6; B = 8'h39; #100;
A = 8'h6; B = 8'h3A; #100;
A = 8'h6; B = 8'h3B; #100;
A = 8'h6; B = 8'h3C; #100;
A = 8'h6; B = 8'h3D; #100;
A = 8'h6; B = 8'h3E; #100;
A = 8'h6; B = 8'h3F; #100;
A = 8'h6; B = 8'h40; #100;
A = 8'h6; B = 8'h41; #100;
A = 8'h6; B = 8'h42; #100;
A = 8'h6; B = 8'h43; #100;
A = 8'h6; B = 8'h44; #100;
A = 8'h6; B = 8'h45; #100;
A = 8'h6; B = 8'h46; #100;
A = 8'h6; B = 8'h47; #100;
A = 8'h6; B = 8'h48; #100;
A = 8'h6; B = 8'h49; #100;
A = 8'h6; B = 8'h4A; #100;
A = 8'h6; B = 8'h4B; #100;
A = 8'h6; B = 8'h4C; #100;
A = 8'h6; B = 8'h4D; #100;
A = 8'h6; B = 8'h4E; #100;
A = 8'h6; B = 8'h4F; #100;
A = 8'h6; B = 8'h50; #100;
A = 8'h6; B = 8'h51; #100;
A = 8'h6; B = 8'h52; #100;
A = 8'h6; B = 8'h53; #100;
A = 8'h6; B = 8'h54; #100;
A = 8'h6; B = 8'h55; #100;
A = 8'h6; B = 8'h56; #100;
A = 8'h6; B = 8'h57; #100;
A = 8'h6; B = 8'h58; #100;
A = 8'h6; B = 8'h59; #100;
A = 8'h6; B = 8'h5A; #100;
A = 8'h6; B = 8'h5B; #100;
A = 8'h6; B = 8'h5C; #100;
A = 8'h6; B = 8'h5D; #100;
A = 8'h6; B = 8'h5E; #100;
A = 8'h6; B = 8'h5F; #100;
A = 8'h6; B = 8'h60; #100;
A = 8'h6; B = 8'h61; #100;
A = 8'h6; B = 8'h62; #100;
A = 8'h6; B = 8'h63; #100;
A = 8'h6; B = 8'h64; #100;
A = 8'h6; B = 8'h65; #100;
A = 8'h6; B = 8'h66; #100;
A = 8'h6; B = 8'h67; #100;
A = 8'h6; B = 8'h68; #100;
A = 8'h6; B = 8'h69; #100;
A = 8'h6; B = 8'h6A; #100;
A = 8'h6; B = 8'h6B; #100;
A = 8'h6; B = 8'h6C; #100;
A = 8'h6; B = 8'h6D; #100;
A = 8'h6; B = 8'h6E; #100;
A = 8'h6; B = 8'h6F; #100;
A = 8'h6; B = 8'h70; #100;
A = 8'h6; B = 8'h71; #100;
A = 8'h6; B = 8'h72; #100;
A = 8'h6; B = 8'h73; #100;
A = 8'h6; B = 8'h74; #100;
A = 8'h6; B = 8'h75; #100;
A = 8'h6; B = 8'h76; #100;
A = 8'h6; B = 8'h77; #100;
A = 8'h6; B = 8'h78; #100;
A = 8'h6; B = 8'h79; #100;
A = 8'h6; B = 8'h7A; #100;
A = 8'h6; B = 8'h7B; #100;
A = 8'h6; B = 8'h7C; #100;
A = 8'h6; B = 8'h7D; #100;
A = 8'h6; B = 8'h7E; #100;
A = 8'h6; B = 8'h7F; #100;
A = 8'h6; B = 8'h80; #100;
A = 8'h6; B = 8'h81; #100;
A = 8'h6; B = 8'h82; #100;
A = 8'h6; B = 8'h83; #100;
A = 8'h6; B = 8'h84; #100;
A = 8'h6; B = 8'h85; #100;
A = 8'h6; B = 8'h86; #100;
A = 8'h6; B = 8'h87; #100;
A = 8'h6; B = 8'h88; #100;
A = 8'h6; B = 8'h89; #100;
A = 8'h6; B = 8'h8A; #100;
A = 8'h6; B = 8'h8B; #100;
A = 8'h6; B = 8'h8C; #100;
A = 8'h6; B = 8'h8D; #100;
A = 8'h6; B = 8'h8E; #100;
A = 8'h6; B = 8'h8F; #100;
A = 8'h6; B = 8'h90; #100;
A = 8'h6; B = 8'h91; #100;
A = 8'h6; B = 8'h92; #100;
A = 8'h6; B = 8'h93; #100;
A = 8'h6; B = 8'h94; #100;
A = 8'h6; B = 8'h95; #100;
A = 8'h6; B = 8'h96; #100;
A = 8'h6; B = 8'h97; #100;
A = 8'h6; B = 8'h98; #100;
A = 8'h6; B = 8'h99; #100;
A = 8'h6; B = 8'h9A; #100;
A = 8'h6; B = 8'h9B; #100;
A = 8'h6; B = 8'h9C; #100;
A = 8'h6; B = 8'h9D; #100;
A = 8'h6; B = 8'h9E; #100;
A = 8'h6; B = 8'h9F; #100;
A = 8'h6; B = 8'hA0; #100;
A = 8'h6; B = 8'hA1; #100;
A = 8'h6; B = 8'hA2; #100;
A = 8'h6; B = 8'hA3; #100;
A = 8'h6; B = 8'hA4; #100;
A = 8'h6; B = 8'hA5; #100;
A = 8'h6; B = 8'hA6; #100;
A = 8'h6; B = 8'hA7; #100;
A = 8'h6; B = 8'hA8; #100;
A = 8'h6; B = 8'hA9; #100;
A = 8'h6; B = 8'hAA; #100;
A = 8'h6; B = 8'hAB; #100;
A = 8'h6; B = 8'hAC; #100;
A = 8'h6; B = 8'hAD; #100;
A = 8'h6; B = 8'hAE; #100;
A = 8'h6; B = 8'hAF; #100;
A = 8'h6; B = 8'hB0; #100;
A = 8'h6; B = 8'hB1; #100;
A = 8'h6; B = 8'hB2; #100;
A = 8'h6; B = 8'hB3; #100;
A = 8'h6; B = 8'hB4; #100;
A = 8'h6; B = 8'hB5; #100;
A = 8'h6; B = 8'hB6; #100;
A = 8'h6; B = 8'hB7; #100;
A = 8'h6; B = 8'hB8; #100;
A = 8'h6; B = 8'hB9; #100;
A = 8'h6; B = 8'hBA; #100;
A = 8'h6; B = 8'hBB; #100;
A = 8'h6; B = 8'hBC; #100;
A = 8'h6; B = 8'hBD; #100;
A = 8'h6; B = 8'hBE; #100;
A = 8'h6; B = 8'hBF; #100;
A = 8'h6; B = 8'hC0; #100;
A = 8'h6; B = 8'hC1; #100;
A = 8'h6; B = 8'hC2; #100;
A = 8'h6; B = 8'hC3; #100;
A = 8'h6; B = 8'hC4; #100;
A = 8'h6; B = 8'hC5; #100;
A = 8'h6; B = 8'hC6; #100;
A = 8'h6; B = 8'hC7; #100;
A = 8'h6; B = 8'hC8; #100;
A = 8'h6; B = 8'hC9; #100;
A = 8'h6; B = 8'hCA; #100;
A = 8'h6; B = 8'hCB; #100;
A = 8'h6; B = 8'hCC; #100;
A = 8'h6; B = 8'hCD; #100;
A = 8'h6; B = 8'hCE; #100;
A = 8'h6; B = 8'hCF; #100;
A = 8'h6; B = 8'hD0; #100;
A = 8'h6; B = 8'hD1; #100;
A = 8'h6; B = 8'hD2; #100;
A = 8'h6; B = 8'hD3; #100;
A = 8'h6; B = 8'hD4; #100;
A = 8'h6; B = 8'hD5; #100;
A = 8'h6; B = 8'hD6; #100;
A = 8'h6; B = 8'hD7; #100;
A = 8'h6; B = 8'hD8; #100;
A = 8'h6; B = 8'hD9; #100;
A = 8'h6; B = 8'hDA; #100;
A = 8'h6; B = 8'hDB; #100;
A = 8'h6; B = 8'hDC; #100;
A = 8'h6; B = 8'hDD; #100;
A = 8'h6; B = 8'hDE; #100;
A = 8'h6; B = 8'hDF; #100;
A = 8'h6; B = 8'hE0; #100;
A = 8'h6; B = 8'hE1; #100;
A = 8'h6; B = 8'hE2; #100;
A = 8'h6; B = 8'hE3; #100;
A = 8'h6; B = 8'hE4; #100;
A = 8'h6; B = 8'hE5; #100;
A = 8'h6; B = 8'hE6; #100;
A = 8'h6; B = 8'hE7; #100;
A = 8'h6; B = 8'hE8; #100;
A = 8'h6; B = 8'hE9; #100;
A = 8'h6; B = 8'hEA; #100;
A = 8'h6; B = 8'hEB; #100;
A = 8'h6; B = 8'hEC; #100;
A = 8'h6; B = 8'hED; #100;
A = 8'h6; B = 8'hEE; #100;
A = 8'h6; B = 8'hEF; #100;
A = 8'h6; B = 8'hF0; #100;
A = 8'h6; B = 8'hF1; #100;
A = 8'h6; B = 8'hF2; #100;
A = 8'h6; B = 8'hF3; #100;
A = 8'h6; B = 8'hF4; #100;
A = 8'h6; B = 8'hF5; #100;
A = 8'h6; B = 8'hF6; #100;
A = 8'h6; B = 8'hF7; #100;
A = 8'h6; B = 8'hF8; #100;
A = 8'h6; B = 8'hF9; #100;
A = 8'h6; B = 8'hFA; #100;
A = 8'h6; B = 8'hFB; #100;
A = 8'h6; B = 8'hFC; #100;
A = 8'h6; B = 8'hFD; #100;
A = 8'h6; B = 8'hFE; #100;
A = 8'h6; B = 8'hFF; #100;
A = 8'h7; B = 8'h0; #100;
A = 8'h7; B = 8'h1; #100;
A = 8'h7; B = 8'h2; #100;
A = 8'h7; B = 8'h3; #100;
A = 8'h7; B = 8'h4; #100;
A = 8'h7; B = 8'h5; #100;
A = 8'h7; B = 8'h6; #100;
A = 8'h7; B = 8'h7; #100;
A = 8'h7; B = 8'h8; #100;
A = 8'h7; B = 8'h9; #100;
A = 8'h7; B = 8'hA; #100;
A = 8'h7; B = 8'hB; #100;
A = 8'h7; B = 8'hC; #100;
A = 8'h7; B = 8'hD; #100;
A = 8'h7; B = 8'hE; #100;
A = 8'h7; B = 8'hF; #100;
A = 8'h7; B = 8'h10; #100;
A = 8'h7; B = 8'h11; #100;
A = 8'h7; B = 8'h12; #100;
A = 8'h7; B = 8'h13; #100;
A = 8'h7; B = 8'h14; #100;
A = 8'h7; B = 8'h15; #100;
A = 8'h7; B = 8'h16; #100;
A = 8'h7; B = 8'h17; #100;
A = 8'h7; B = 8'h18; #100;
A = 8'h7; B = 8'h19; #100;
A = 8'h7; B = 8'h1A; #100;
A = 8'h7; B = 8'h1B; #100;
A = 8'h7; B = 8'h1C; #100;
A = 8'h7; B = 8'h1D; #100;
A = 8'h7; B = 8'h1E; #100;
A = 8'h7; B = 8'h1F; #100;
A = 8'h7; B = 8'h20; #100;
A = 8'h7; B = 8'h21; #100;
A = 8'h7; B = 8'h22; #100;
A = 8'h7; B = 8'h23; #100;
A = 8'h7; B = 8'h24; #100;
A = 8'h7; B = 8'h25; #100;
A = 8'h7; B = 8'h26; #100;
A = 8'h7; B = 8'h27; #100;
A = 8'h7; B = 8'h28; #100;
A = 8'h7; B = 8'h29; #100;
A = 8'h7; B = 8'h2A; #100;
A = 8'h7; B = 8'h2B; #100;
A = 8'h7; B = 8'h2C; #100;
A = 8'h7; B = 8'h2D; #100;
A = 8'h7; B = 8'h2E; #100;
A = 8'h7; B = 8'h2F; #100;
A = 8'h7; B = 8'h30; #100;
A = 8'h7; B = 8'h31; #100;
A = 8'h7; B = 8'h32; #100;
A = 8'h7; B = 8'h33; #100;
A = 8'h7; B = 8'h34; #100;
A = 8'h7; B = 8'h35; #100;
A = 8'h7; B = 8'h36; #100;
A = 8'h7; B = 8'h37; #100;
A = 8'h7; B = 8'h38; #100;
A = 8'h7; B = 8'h39; #100;
A = 8'h7; B = 8'h3A; #100;
A = 8'h7; B = 8'h3B; #100;
A = 8'h7; B = 8'h3C; #100;
A = 8'h7; B = 8'h3D; #100;
A = 8'h7; B = 8'h3E; #100;
A = 8'h7; B = 8'h3F; #100;
A = 8'h7; B = 8'h40; #100;
A = 8'h7; B = 8'h41; #100;
A = 8'h7; B = 8'h42; #100;
A = 8'h7; B = 8'h43; #100;
A = 8'h7; B = 8'h44; #100;
A = 8'h7; B = 8'h45; #100;
A = 8'h7; B = 8'h46; #100;
A = 8'h7; B = 8'h47; #100;
A = 8'h7; B = 8'h48; #100;
A = 8'h7; B = 8'h49; #100;
A = 8'h7; B = 8'h4A; #100;
A = 8'h7; B = 8'h4B; #100;
A = 8'h7; B = 8'h4C; #100;
A = 8'h7; B = 8'h4D; #100;
A = 8'h7; B = 8'h4E; #100;
A = 8'h7; B = 8'h4F; #100;
A = 8'h7; B = 8'h50; #100;
A = 8'h7; B = 8'h51; #100;
A = 8'h7; B = 8'h52; #100;
A = 8'h7; B = 8'h53; #100;
A = 8'h7; B = 8'h54; #100;
A = 8'h7; B = 8'h55; #100;
A = 8'h7; B = 8'h56; #100;
A = 8'h7; B = 8'h57; #100;
A = 8'h7; B = 8'h58; #100;
A = 8'h7; B = 8'h59; #100;
A = 8'h7; B = 8'h5A; #100;
A = 8'h7; B = 8'h5B; #100;
A = 8'h7; B = 8'h5C; #100;
A = 8'h7; B = 8'h5D; #100;
A = 8'h7; B = 8'h5E; #100;
A = 8'h7; B = 8'h5F; #100;
A = 8'h7; B = 8'h60; #100;
A = 8'h7; B = 8'h61; #100;
A = 8'h7; B = 8'h62; #100;
A = 8'h7; B = 8'h63; #100;
A = 8'h7; B = 8'h64; #100;
A = 8'h7; B = 8'h65; #100;
A = 8'h7; B = 8'h66; #100;
A = 8'h7; B = 8'h67; #100;
A = 8'h7; B = 8'h68; #100;
A = 8'h7; B = 8'h69; #100;
A = 8'h7; B = 8'h6A; #100;
A = 8'h7; B = 8'h6B; #100;
A = 8'h7; B = 8'h6C; #100;
A = 8'h7; B = 8'h6D; #100;
A = 8'h7; B = 8'h6E; #100;
A = 8'h7; B = 8'h6F; #100;
A = 8'h7; B = 8'h70; #100;
A = 8'h7; B = 8'h71; #100;
A = 8'h7; B = 8'h72; #100;
A = 8'h7; B = 8'h73; #100;
A = 8'h7; B = 8'h74; #100;
A = 8'h7; B = 8'h75; #100;
A = 8'h7; B = 8'h76; #100;
A = 8'h7; B = 8'h77; #100;
A = 8'h7; B = 8'h78; #100;
A = 8'h7; B = 8'h79; #100;
A = 8'h7; B = 8'h7A; #100;
A = 8'h7; B = 8'h7B; #100;
A = 8'h7; B = 8'h7C; #100;
A = 8'h7; B = 8'h7D; #100;
A = 8'h7; B = 8'h7E; #100;
A = 8'h7; B = 8'h7F; #100;
A = 8'h7; B = 8'h80; #100;
A = 8'h7; B = 8'h81; #100;
A = 8'h7; B = 8'h82; #100;
A = 8'h7; B = 8'h83; #100;
A = 8'h7; B = 8'h84; #100;
A = 8'h7; B = 8'h85; #100;
A = 8'h7; B = 8'h86; #100;
A = 8'h7; B = 8'h87; #100;
A = 8'h7; B = 8'h88; #100;
A = 8'h7; B = 8'h89; #100;
A = 8'h7; B = 8'h8A; #100;
A = 8'h7; B = 8'h8B; #100;
A = 8'h7; B = 8'h8C; #100;
A = 8'h7; B = 8'h8D; #100;
A = 8'h7; B = 8'h8E; #100;
A = 8'h7; B = 8'h8F; #100;
A = 8'h7; B = 8'h90; #100;
A = 8'h7; B = 8'h91; #100;
A = 8'h7; B = 8'h92; #100;
A = 8'h7; B = 8'h93; #100;
A = 8'h7; B = 8'h94; #100;
A = 8'h7; B = 8'h95; #100;
A = 8'h7; B = 8'h96; #100;
A = 8'h7; B = 8'h97; #100;
A = 8'h7; B = 8'h98; #100;
A = 8'h7; B = 8'h99; #100;
A = 8'h7; B = 8'h9A; #100;
A = 8'h7; B = 8'h9B; #100;
A = 8'h7; B = 8'h9C; #100;
A = 8'h7; B = 8'h9D; #100;
A = 8'h7; B = 8'h9E; #100;
A = 8'h7; B = 8'h9F; #100;
A = 8'h7; B = 8'hA0; #100;
A = 8'h7; B = 8'hA1; #100;
A = 8'h7; B = 8'hA2; #100;
A = 8'h7; B = 8'hA3; #100;
A = 8'h7; B = 8'hA4; #100;
A = 8'h7; B = 8'hA5; #100;
A = 8'h7; B = 8'hA6; #100;
A = 8'h7; B = 8'hA7; #100;
A = 8'h7; B = 8'hA8; #100;
A = 8'h7; B = 8'hA9; #100;
A = 8'h7; B = 8'hAA; #100;
A = 8'h7; B = 8'hAB; #100;
A = 8'h7; B = 8'hAC; #100;
A = 8'h7; B = 8'hAD; #100;
A = 8'h7; B = 8'hAE; #100;
A = 8'h7; B = 8'hAF; #100;
A = 8'h7; B = 8'hB0; #100;
A = 8'h7; B = 8'hB1; #100;
A = 8'h7; B = 8'hB2; #100;
A = 8'h7; B = 8'hB3; #100;
A = 8'h7; B = 8'hB4; #100;
A = 8'h7; B = 8'hB5; #100;
A = 8'h7; B = 8'hB6; #100;
A = 8'h7; B = 8'hB7; #100;
A = 8'h7; B = 8'hB8; #100;
A = 8'h7; B = 8'hB9; #100;
A = 8'h7; B = 8'hBA; #100;
A = 8'h7; B = 8'hBB; #100;
A = 8'h7; B = 8'hBC; #100;
A = 8'h7; B = 8'hBD; #100;
A = 8'h7; B = 8'hBE; #100;
A = 8'h7; B = 8'hBF; #100;
A = 8'h7; B = 8'hC0; #100;
A = 8'h7; B = 8'hC1; #100;
A = 8'h7; B = 8'hC2; #100;
A = 8'h7; B = 8'hC3; #100;
A = 8'h7; B = 8'hC4; #100;
A = 8'h7; B = 8'hC5; #100;
A = 8'h7; B = 8'hC6; #100;
A = 8'h7; B = 8'hC7; #100;
A = 8'h7; B = 8'hC8; #100;
A = 8'h7; B = 8'hC9; #100;
A = 8'h7; B = 8'hCA; #100;
A = 8'h7; B = 8'hCB; #100;
A = 8'h7; B = 8'hCC; #100;
A = 8'h7; B = 8'hCD; #100;
A = 8'h7; B = 8'hCE; #100;
A = 8'h7; B = 8'hCF; #100;
A = 8'h7; B = 8'hD0; #100;
A = 8'h7; B = 8'hD1; #100;
A = 8'h7; B = 8'hD2; #100;
A = 8'h7; B = 8'hD3; #100;
A = 8'h7; B = 8'hD4; #100;
A = 8'h7; B = 8'hD5; #100;
A = 8'h7; B = 8'hD6; #100;
A = 8'h7; B = 8'hD7; #100;
A = 8'h7; B = 8'hD8; #100;
A = 8'h7; B = 8'hD9; #100;
A = 8'h7; B = 8'hDA; #100;
A = 8'h7; B = 8'hDB; #100;
A = 8'h7; B = 8'hDC; #100;
A = 8'h7; B = 8'hDD; #100;
A = 8'h7; B = 8'hDE; #100;
A = 8'h7; B = 8'hDF; #100;
A = 8'h7; B = 8'hE0; #100;
A = 8'h7; B = 8'hE1; #100;
A = 8'h7; B = 8'hE2; #100;
A = 8'h7; B = 8'hE3; #100;
A = 8'h7; B = 8'hE4; #100;
A = 8'h7; B = 8'hE5; #100;
A = 8'h7; B = 8'hE6; #100;
A = 8'h7; B = 8'hE7; #100;
A = 8'h7; B = 8'hE8; #100;
A = 8'h7; B = 8'hE9; #100;
A = 8'h7; B = 8'hEA; #100;
A = 8'h7; B = 8'hEB; #100;
A = 8'h7; B = 8'hEC; #100;
A = 8'h7; B = 8'hED; #100;
A = 8'h7; B = 8'hEE; #100;
A = 8'h7; B = 8'hEF; #100;
A = 8'h7; B = 8'hF0; #100;
A = 8'h7; B = 8'hF1; #100;
A = 8'h7; B = 8'hF2; #100;
A = 8'h7; B = 8'hF3; #100;
A = 8'h7; B = 8'hF4; #100;
A = 8'h7; B = 8'hF5; #100;
A = 8'h7; B = 8'hF6; #100;
A = 8'h7; B = 8'hF7; #100;
A = 8'h7; B = 8'hF8; #100;
A = 8'h7; B = 8'hF9; #100;
A = 8'h7; B = 8'hFA; #100;
A = 8'h7; B = 8'hFB; #100;
A = 8'h7; B = 8'hFC; #100;
A = 8'h7; B = 8'hFD; #100;
A = 8'h7; B = 8'hFE; #100;
A = 8'h7; B = 8'hFF; #100;
A = 8'h8; B = 8'h0; #100;
A = 8'h8; B = 8'h1; #100;
A = 8'h8; B = 8'h2; #100;
A = 8'h8; B = 8'h3; #100;
A = 8'h8; B = 8'h4; #100;
A = 8'h8; B = 8'h5; #100;
A = 8'h8; B = 8'h6; #100;
A = 8'h8; B = 8'h7; #100;
A = 8'h8; B = 8'h8; #100;
A = 8'h8; B = 8'h9; #100;
A = 8'h8; B = 8'hA; #100;
A = 8'h8; B = 8'hB; #100;
A = 8'h8; B = 8'hC; #100;
A = 8'h8; B = 8'hD; #100;
A = 8'h8; B = 8'hE; #100;
A = 8'h8; B = 8'hF; #100;
A = 8'h8; B = 8'h10; #100;
A = 8'h8; B = 8'h11; #100;
A = 8'h8; B = 8'h12; #100;
A = 8'h8; B = 8'h13; #100;
A = 8'h8; B = 8'h14; #100;
A = 8'h8; B = 8'h15; #100;
A = 8'h8; B = 8'h16; #100;
A = 8'h8; B = 8'h17; #100;
A = 8'h8; B = 8'h18; #100;
A = 8'h8; B = 8'h19; #100;
A = 8'h8; B = 8'h1A; #100;
A = 8'h8; B = 8'h1B; #100;
A = 8'h8; B = 8'h1C; #100;
A = 8'h8; B = 8'h1D; #100;
A = 8'h8; B = 8'h1E; #100;
A = 8'h8; B = 8'h1F; #100;
A = 8'h8; B = 8'h20; #100;
A = 8'h8; B = 8'h21; #100;
A = 8'h8; B = 8'h22; #100;
A = 8'h8; B = 8'h23; #100;
A = 8'h8; B = 8'h24; #100;
A = 8'h8; B = 8'h25; #100;
A = 8'h8; B = 8'h26; #100;
A = 8'h8; B = 8'h27; #100;
A = 8'h8; B = 8'h28; #100;
A = 8'h8; B = 8'h29; #100;
A = 8'h8; B = 8'h2A; #100;
A = 8'h8; B = 8'h2B; #100;
A = 8'h8; B = 8'h2C; #100;
A = 8'h8; B = 8'h2D; #100;
A = 8'h8; B = 8'h2E; #100;
A = 8'h8; B = 8'h2F; #100;
A = 8'h8; B = 8'h30; #100;
A = 8'h8; B = 8'h31; #100;
A = 8'h8; B = 8'h32; #100;
A = 8'h8; B = 8'h33; #100;
A = 8'h8; B = 8'h34; #100;
A = 8'h8; B = 8'h35; #100;
A = 8'h8; B = 8'h36; #100;
A = 8'h8; B = 8'h37; #100;
A = 8'h8; B = 8'h38; #100;
A = 8'h8; B = 8'h39; #100;
A = 8'h8; B = 8'h3A; #100;
A = 8'h8; B = 8'h3B; #100;
A = 8'h8; B = 8'h3C; #100;
A = 8'h8; B = 8'h3D; #100;
A = 8'h8; B = 8'h3E; #100;
A = 8'h8; B = 8'h3F; #100;
A = 8'h8; B = 8'h40; #100;
A = 8'h8; B = 8'h41; #100;
A = 8'h8; B = 8'h42; #100;
A = 8'h8; B = 8'h43; #100;
A = 8'h8; B = 8'h44; #100;
A = 8'h8; B = 8'h45; #100;
A = 8'h8; B = 8'h46; #100;
A = 8'h8; B = 8'h47; #100;
A = 8'h8; B = 8'h48; #100;
A = 8'h8; B = 8'h49; #100;
A = 8'h8; B = 8'h4A; #100;
A = 8'h8; B = 8'h4B; #100;
A = 8'h8; B = 8'h4C; #100;
A = 8'h8; B = 8'h4D; #100;
A = 8'h8; B = 8'h4E; #100;
A = 8'h8; B = 8'h4F; #100;
A = 8'h8; B = 8'h50; #100;
A = 8'h8; B = 8'h51; #100;
A = 8'h8; B = 8'h52; #100;
A = 8'h8; B = 8'h53; #100;
A = 8'h8; B = 8'h54; #100;
A = 8'h8; B = 8'h55; #100;
A = 8'h8; B = 8'h56; #100;
A = 8'h8; B = 8'h57; #100;
A = 8'h8; B = 8'h58; #100;
A = 8'h8; B = 8'h59; #100;
A = 8'h8; B = 8'h5A; #100;
A = 8'h8; B = 8'h5B; #100;
A = 8'h8; B = 8'h5C; #100;
A = 8'h8; B = 8'h5D; #100;
A = 8'h8; B = 8'h5E; #100;
A = 8'h8; B = 8'h5F; #100;
A = 8'h8; B = 8'h60; #100;
A = 8'h8; B = 8'h61; #100;
A = 8'h8; B = 8'h62; #100;
A = 8'h8; B = 8'h63; #100;
A = 8'h8; B = 8'h64; #100;
A = 8'h8; B = 8'h65; #100;
A = 8'h8; B = 8'h66; #100;
A = 8'h8; B = 8'h67; #100;
A = 8'h8; B = 8'h68; #100;
A = 8'h8; B = 8'h69; #100;
A = 8'h8; B = 8'h6A; #100;
A = 8'h8; B = 8'h6B; #100;
A = 8'h8; B = 8'h6C; #100;
A = 8'h8; B = 8'h6D; #100;
A = 8'h8; B = 8'h6E; #100;
A = 8'h8; B = 8'h6F; #100;
A = 8'h8; B = 8'h70; #100;
A = 8'h8; B = 8'h71; #100;
A = 8'h8; B = 8'h72; #100;
A = 8'h8; B = 8'h73; #100;
A = 8'h8; B = 8'h74; #100;
A = 8'h8; B = 8'h75; #100;
A = 8'h8; B = 8'h76; #100;
A = 8'h8; B = 8'h77; #100;
A = 8'h8; B = 8'h78; #100;
A = 8'h8; B = 8'h79; #100;
A = 8'h8; B = 8'h7A; #100;
A = 8'h8; B = 8'h7B; #100;
A = 8'h8; B = 8'h7C; #100;
A = 8'h8; B = 8'h7D; #100;
A = 8'h8; B = 8'h7E; #100;
A = 8'h8; B = 8'h7F; #100;
A = 8'h8; B = 8'h80; #100;
A = 8'h8; B = 8'h81; #100;
A = 8'h8; B = 8'h82; #100;
A = 8'h8; B = 8'h83; #100;
A = 8'h8; B = 8'h84; #100;
A = 8'h8; B = 8'h85; #100;
A = 8'h8; B = 8'h86; #100;
A = 8'h8; B = 8'h87; #100;
A = 8'h8; B = 8'h88; #100;
A = 8'h8; B = 8'h89; #100;
A = 8'h8; B = 8'h8A; #100;
A = 8'h8; B = 8'h8B; #100;
A = 8'h8; B = 8'h8C; #100;
A = 8'h8; B = 8'h8D; #100;
A = 8'h8; B = 8'h8E; #100;
A = 8'h8; B = 8'h8F; #100;
A = 8'h8; B = 8'h90; #100;
A = 8'h8; B = 8'h91; #100;
A = 8'h8; B = 8'h92; #100;
A = 8'h8; B = 8'h93; #100;
A = 8'h8; B = 8'h94; #100;
A = 8'h8; B = 8'h95; #100;
A = 8'h8; B = 8'h96; #100;
A = 8'h8; B = 8'h97; #100;
A = 8'h8; B = 8'h98; #100;
A = 8'h8; B = 8'h99; #100;
A = 8'h8; B = 8'h9A; #100;
A = 8'h8; B = 8'h9B; #100;
A = 8'h8; B = 8'h9C; #100;
A = 8'h8; B = 8'h9D; #100;
A = 8'h8; B = 8'h9E; #100;
A = 8'h8; B = 8'h9F; #100;
A = 8'h8; B = 8'hA0; #100;
A = 8'h8; B = 8'hA1; #100;
A = 8'h8; B = 8'hA2; #100;
A = 8'h8; B = 8'hA3; #100;
A = 8'h8; B = 8'hA4; #100;
A = 8'h8; B = 8'hA5; #100;
A = 8'h8; B = 8'hA6; #100;
A = 8'h8; B = 8'hA7; #100;
A = 8'h8; B = 8'hA8; #100;
A = 8'h8; B = 8'hA9; #100;
A = 8'h8; B = 8'hAA; #100;
A = 8'h8; B = 8'hAB; #100;
A = 8'h8; B = 8'hAC; #100;
A = 8'h8; B = 8'hAD; #100;
A = 8'h8; B = 8'hAE; #100;
A = 8'h8; B = 8'hAF; #100;
A = 8'h8; B = 8'hB0; #100;
A = 8'h8; B = 8'hB1; #100;
A = 8'h8; B = 8'hB2; #100;
A = 8'h8; B = 8'hB3; #100;
A = 8'h8; B = 8'hB4; #100;
A = 8'h8; B = 8'hB5; #100;
A = 8'h8; B = 8'hB6; #100;
A = 8'h8; B = 8'hB7; #100;
A = 8'h8; B = 8'hB8; #100;
A = 8'h8; B = 8'hB9; #100;
A = 8'h8; B = 8'hBA; #100;
A = 8'h8; B = 8'hBB; #100;
A = 8'h8; B = 8'hBC; #100;
A = 8'h8; B = 8'hBD; #100;
A = 8'h8; B = 8'hBE; #100;
A = 8'h8; B = 8'hBF; #100;
A = 8'h8; B = 8'hC0; #100;
A = 8'h8; B = 8'hC1; #100;
A = 8'h8; B = 8'hC2; #100;
A = 8'h8; B = 8'hC3; #100;
A = 8'h8; B = 8'hC4; #100;
A = 8'h8; B = 8'hC5; #100;
A = 8'h8; B = 8'hC6; #100;
A = 8'h8; B = 8'hC7; #100;
A = 8'h8; B = 8'hC8; #100;
A = 8'h8; B = 8'hC9; #100;
A = 8'h8; B = 8'hCA; #100;
A = 8'h8; B = 8'hCB; #100;
A = 8'h8; B = 8'hCC; #100;
A = 8'h8; B = 8'hCD; #100;
A = 8'h8; B = 8'hCE; #100;
A = 8'h8; B = 8'hCF; #100;
A = 8'h8; B = 8'hD0; #100;
A = 8'h8; B = 8'hD1; #100;
A = 8'h8; B = 8'hD2; #100;
A = 8'h8; B = 8'hD3; #100;
A = 8'h8; B = 8'hD4; #100;
A = 8'h8; B = 8'hD5; #100;
A = 8'h8; B = 8'hD6; #100;
A = 8'h8; B = 8'hD7; #100;
A = 8'h8; B = 8'hD8; #100;
A = 8'h8; B = 8'hD9; #100;
A = 8'h8; B = 8'hDA; #100;
A = 8'h8; B = 8'hDB; #100;
A = 8'h8; B = 8'hDC; #100;
A = 8'h8; B = 8'hDD; #100;
A = 8'h8; B = 8'hDE; #100;
A = 8'h8; B = 8'hDF; #100;
A = 8'h8; B = 8'hE0; #100;
A = 8'h8; B = 8'hE1; #100;
A = 8'h8; B = 8'hE2; #100;
A = 8'h8; B = 8'hE3; #100;
A = 8'h8; B = 8'hE4; #100;
A = 8'h8; B = 8'hE5; #100;
A = 8'h8; B = 8'hE6; #100;
A = 8'h8; B = 8'hE7; #100;
A = 8'h8; B = 8'hE8; #100;
A = 8'h8; B = 8'hE9; #100;
A = 8'h8; B = 8'hEA; #100;
A = 8'h8; B = 8'hEB; #100;
A = 8'h8; B = 8'hEC; #100;
A = 8'h8; B = 8'hED; #100;
A = 8'h8; B = 8'hEE; #100;
A = 8'h8; B = 8'hEF; #100;
A = 8'h8; B = 8'hF0; #100;
A = 8'h8; B = 8'hF1; #100;
A = 8'h8; B = 8'hF2; #100;
A = 8'h8; B = 8'hF3; #100;
A = 8'h8; B = 8'hF4; #100;
A = 8'h8; B = 8'hF5; #100;
A = 8'h8; B = 8'hF6; #100;
A = 8'h8; B = 8'hF7; #100;
A = 8'h8; B = 8'hF8; #100;
A = 8'h8; B = 8'hF9; #100;
A = 8'h8; B = 8'hFA; #100;
A = 8'h8; B = 8'hFB; #100;
A = 8'h8; B = 8'hFC; #100;
A = 8'h8; B = 8'hFD; #100;
A = 8'h8; B = 8'hFE; #100;
A = 8'h8; B = 8'hFF; #100;
A = 8'h9; B = 8'h0; #100;
A = 8'h9; B = 8'h1; #100;
A = 8'h9; B = 8'h2; #100;
A = 8'h9; B = 8'h3; #100;
A = 8'h9; B = 8'h4; #100;
A = 8'h9; B = 8'h5; #100;
A = 8'h9; B = 8'h6; #100;
A = 8'h9; B = 8'h7; #100;
A = 8'h9; B = 8'h8; #100;
A = 8'h9; B = 8'h9; #100;
A = 8'h9; B = 8'hA; #100;
A = 8'h9; B = 8'hB; #100;
A = 8'h9; B = 8'hC; #100;
A = 8'h9; B = 8'hD; #100;
A = 8'h9; B = 8'hE; #100;
A = 8'h9; B = 8'hF; #100;
A = 8'h9; B = 8'h10; #100;
A = 8'h9; B = 8'h11; #100;
A = 8'h9; B = 8'h12; #100;
A = 8'h9; B = 8'h13; #100;
A = 8'h9; B = 8'h14; #100;
A = 8'h9; B = 8'h15; #100;
A = 8'h9; B = 8'h16; #100;
A = 8'h9; B = 8'h17; #100;
A = 8'h9; B = 8'h18; #100;
A = 8'h9; B = 8'h19; #100;
A = 8'h9; B = 8'h1A; #100;
A = 8'h9; B = 8'h1B; #100;
A = 8'h9; B = 8'h1C; #100;
A = 8'h9; B = 8'h1D; #100;
A = 8'h9; B = 8'h1E; #100;
A = 8'h9; B = 8'h1F; #100;
A = 8'h9; B = 8'h20; #100;
A = 8'h9; B = 8'h21; #100;
A = 8'h9; B = 8'h22; #100;
A = 8'h9; B = 8'h23; #100;
A = 8'h9; B = 8'h24; #100;
A = 8'h9; B = 8'h25; #100;
A = 8'h9; B = 8'h26; #100;
A = 8'h9; B = 8'h27; #100;
A = 8'h9; B = 8'h28; #100;
A = 8'h9; B = 8'h29; #100;
A = 8'h9; B = 8'h2A; #100;
A = 8'h9; B = 8'h2B; #100;
A = 8'h9; B = 8'h2C; #100;
A = 8'h9; B = 8'h2D; #100;
A = 8'h9; B = 8'h2E; #100;
A = 8'h9; B = 8'h2F; #100;
A = 8'h9; B = 8'h30; #100;
A = 8'h9; B = 8'h31; #100;
A = 8'h9; B = 8'h32; #100;
A = 8'h9; B = 8'h33; #100;
A = 8'h9; B = 8'h34; #100;
A = 8'h9; B = 8'h35; #100;
A = 8'h9; B = 8'h36; #100;
A = 8'h9; B = 8'h37; #100;
A = 8'h9; B = 8'h38; #100;
A = 8'h9; B = 8'h39; #100;
A = 8'h9; B = 8'h3A; #100;
A = 8'h9; B = 8'h3B; #100;
A = 8'h9; B = 8'h3C; #100;
A = 8'h9; B = 8'h3D; #100;
A = 8'h9; B = 8'h3E; #100;
A = 8'h9; B = 8'h3F; #100;
A = 8'h9; B = 8'h40; #100;
A = 8'h9; B = 8'h41; #100;
A = 8'h9; B = 8'h42; #100;
A = 8'h9; B = 8'h43; #100;
A = 8'h9; B = 8'h44; #100;
A = 8'h9; B = 8'h45; #100;
A = 8'h9; B = 8'h46; #100;
A = 8'h9; B = 8'h47; #100;
A = 8'h9; B = 8'h48; #100;
A = 8'h9; B = 8'h49; #100;
A = 8'h9; B = 8'h4A; #100;
A = 8'h9; B = 8'h4B; #100;
A = 8'h9; B = 8'h4C; #100;
A = 8'h9; B = 8'h4D; #100;
A = 8'h9; B = 8'h4E; #100;
A = 8'h9; B = 8'h4F; #100;
A = 8'h9; B = 8'h50; #100;
A = 8'h9; B = 8'h51; #100;
A = 8'h9; B = 8'h52; #100;
A = 8'h9; B = 8'h53; #100;
A = 8'h9; B = 8'h54; #100;
A = 8'h9; B = 8'h55; #100;
A = 8'h9; B = 8'h56; #100;
A = 8'h9; B = 8'h57; #100;
A = 8'h9; B = 8'h58; #100;
A = 8'h9; B = 8'h59; #100;
A = 8'h9; B = 8'h5A; #100;
A = 8'h9; B = 8'h5B; #100;
A = 8'h9; B = 8'h5C; #100;
A = 8'h9; B = 8'h5D; #100;
A = 8'h9; B = 8'h5E; #100;
A = 8'h9; B = 8'h5F; #100;
A = 8'h9; B = 8'h60; #100;
A = 8'h9; B = 8'h61; #100;
A = 8'h9; B = 8'h62; #100;
A = 8'h9; B = 8'h63; #100;
A = 8'h9; B = 8'h64; #100;
A = 8'h9; B = 8'h65; #100;
A = 8'h9; B = 8'h66; #100;
A = 8'h9; B = 8'h67; #100;
A = 8'h9; B = 8'h68; #100;
A = 8'h9; B = 8'h69; #100;
A = 8'h9; B = 8'h6A; #100;
A = 8'h9; B = 8'h6B; #100;
A = 8'h9; B = 8'h6C; #100;
A = 8'h9; B = 8'h6D; #100;
A = 8'h9; B = 8'h6E; #100;
A = 8'h9; B = 8'h6F; #100;
A = 8'h9; B = 8'h70; #100;
A = 8'h9; B = 8'h71; #100;
A = 8'h9; B = 8'h72; #100;
A = 8'h9; B = 8'h73; #100;
A = 8'h9; B = 8'h74; #100;
A = 8'h9; B = 8'h75; #100;
A = 8'h9; B = 8'h76; #100;
A = 8'h9; B = 8'h77; #100;
A = 8'h9; B = 8'h78; #100;
A = 8'h9; B = 8'h79; #100;
A = 8'h9; B = 8'h7A; #100;
A = 8'h9; B = 8'h7B; #100;
A = 8'h9; B = 8'h7C; #100;
A = 8'h9; B = 8'h7D; #100;
A = 8'h9; B = 8'h7E; #100;
A = 8'h9; B = 8'h7F; #100;
A = 8'h9; B = 8'h80; #100;
A = 8'h9; B = 8'h81; #100;
A = 8'h9; B = 8'h82; #100;
A = 8'h9; B = 8'h83; #100;
A = 8'h9; B = 8'h84; #100;
A = 8'h9; B = 8'h85; #100;
A = 8'h9; B = 8'h86; #100;
A = 8'h9; B = 8'h87; #100;
A = 8'h9; B = 8'h88; #100;
A = 8'h9; B = 8'h89; #100;
A = 8'h9; B = 8'h8A; #100;
A = 8'h9; B = 8'h8B; #100;
A = 8'h9; B = 8'h8C; #100;
A = 8'h9; B = 8'h8D; #100;
A = 8'h9; B = 8'h8E; #100;
A = 8'h9; B = 8'h8F; #100;
A = 8'h9; B = 8'h90; #100;
A = 8'h9; B = 8'h91; #100;
A = 8'h9; B = 8'h92; #100;
A = 8'h9; B = 8'h93; #100;
A = 8'h9; B = 8'h94; #100;
A = 8'h9; B = 8'h95; #100;
A = 8'h9; B = 8'h96; #100;
A = 8'h9; B = 8'h97; #100;
A = 8'h9; B = 8'h98; #100;
A = 8'h9; B = 8'h99; #100;
A = 8'h9; B = 8'h9A; #100;
A = 8'h9; B = 8'h9B; #100;
A = 8'h9; B = 8'h9C; #100;
A = 8'h9; B = 8'h9D; #100;
A = 8'h9; B = 8'h9E; #100;
A = 8'h9; B = 8'h9F; #100;
A = 8'h9; B = 8'hA0; #100;
A = 8'h9; B = 8'hA1; #100;
A = 8'h9; B = 8'hA2; #100;
A = 8'h9; B = 8'hA3; #100;
A = 8'h9; B = 8'hA4; #100;
A = 8'h9; B = 8'hA5; #100;
A = 8'h9; B = 8'hA6; #100;
A = 8'h9; B = 8'hA7; #100;
A = 8'h9; B = 8'hA8; #100;
A = 8'h9; B = 8'hA9; #100;
A = 8'h9; B = 8'hAA; #100;
A = 8'h9; B = 8'hAB; #100;
A = 8'h9; B = 8'hAC; #100;
A = 8'h9; B = 8'hAD; #100;
A = 8'h9; B = 8'hAE; #100;
A = 8'h9; B = 8'hAF; #100;
A = 8'h9; B = 8'hB0; #100;
A = 8'h9; B = 8'hB1; #100;
A = 8'h9; B = 8'hB2; #100;
A = 8'h9; B = 8'hB3; #100;
A = 8'h9; B = 8'hB4; #100;
A = 8'h9; B = 8'hB5; #100;
A = 8'h9; B = 8'hB6; #100;
A = 8'h9; B = 8'hB7; #100;
A = 8'h9; B = 8'hB8; #100;
A = 8'h9; B = 8'hB9; #100;
A = 8'h9; B = 8'hBA; #100;
A = 8'h9; B = 8'hBB; #100;
A = 8'h9; B = 8'hBC; #100;
A = 8'h9; B = 8'hBD; #100;
A = 8'h9; B = 8'hBE; #100;
A = 8'h9; B = 8'hBF; #100;
A = 8'h9; B = 8'hC0; #100;
A = 8'h9; B = 8'hC1; #100;
A = 8'h9; B = 8'hC2; #100;
A = 8'h9; B = 8'hC3; #100;
A = 8'h9; B = 8'hC4; #100;
A = 8'h9; B = 8'hC5; #100;
A = 8'h9; B = 8'hC6; #100;
A = 8'h9; B = 8'hC7; #100;
A = 8'h9; B = 8'hC8; #100;
A = 8'h9; B = 8'hC9; #100;
A = 8'h9; B = 8'hCA; #100;
A = 8'h9; B = 8'hCB; #100;
A = 8'h9; B = 8'hCC; #100;
A = 8'h9; B = 8'hCD; #100;
A = 8'h9; B = 8'hCE; #100;
A = 8'h9; B = 8'hCF; #100;
A = 8'h9; B = 8'hD0; #100;
A = 8'h9; B = 8'hD1; #100;
A = 8'h9; B = 8'hD2; #100;
A = 8'h9; B = 8'hD3; #100;
A = 8'h9; B = 8'hD4; #100;
A = 8'h9; B = 8'hD5; #100;
A = 8'h9; B = 8'hD6; #100;
A = 8'h9; B = 8'hD7; #100;
A = 8'h9; B = 8'hD8; #100;
A = 8'h9; B = 8'hD9; #100;
A = 8'h9; B = 8'hDA; #100;
A = 8'h9; B = 8'hDB; #100;
A = 8'h9; B = 8'hDC; #100;
A = 8'h9; B = 8'hDD; #100;
A = 8'h9; B = 8'hDE; #100;
A = 8'h9; B = 8'hDF; #100;
A = 8'h9; B = 8'hE0; #100;
A = 8'h9; B = 8'hE1; #100;
A = 8'h9; B = 8'hE2; #100;
A = 8'h9; B = 8'hE3; #100;
A = 8'h9; B = 8'hE4; #100;
A = 8'h9; B = 8'hE5; #100;
A = 8'h9; B = 8'hE6; #100;
A = 8'h9; B = 8'hE7; #100;
A = 8'h9; B = 8'hE8; #100;
A = 8'h9; B = 8'hE9; #100;
A = 8'h9; B = 8'hEA; #100;
A = 8'h9; B = 8'hEB; #100;
A = 8'h9; B = 8'hEC; #100;
A = 8'h9; B = 8'hED; #100;
A = 8'h9; B = 8'hEE; #100;
A = 8'h9; B = 8'hEF; #100;
A = 8'h9; B = 8'hF0; #100;
A = 8'h9; B = 8'hF1; #100;
A = 8'h9; B = 8'hF2; #100;
A = 8'h9; B = 8'hF3; #100;
A = 8'h9; B = 8'hF4; #100;
A = 8'h9; B = 8'hF5; #100;
A = 8'h9; B = 8'hF6; #100;
A = 8'h9; B = 8'hF7; #100;
A = 8'h9; B = 8'hF8; #100;
A = 8'h9; B = 8'hF9; #100;
A = 8'h9; B = 8'hFA; #100;
A = 8'h9; B = 8'hFB; #100;
A = 8'h9; B = 8'hFC; #100;
A = 8'h9; B = 8'hFD; #100;
A = 8'h9; B = 8'hFE; #100;
A = 8'h9; B = 8'hFF; #100;
A = 8'hA; B = 8'h0; #100;
A = 8'hA; B = 8'h1; #100;
A = 8'hA; B = 8'h2; #100;
A = 8'hA; B = 8'h3; #100;
A = 8'hA; B = 8'h4; #100;
A = 8'hA; B = 8'h5; #100;
A = 8'hA; B = 8'h6; #100;
A = 8'hA; B = 8'h7; #100;
A = 8'hA; B = 8'h8; #100;
A = 8'hA; B = 8'h9; #100;
A = 8'hA; B = 8'hA; #100;
A = 8'hA; B = 8'hB; #100;
A = 8'hA; B = 8'hC; #100;
A = 8'hA; B = 8'hD; #100;
A = 8'hA; B = 8'hE; #100;
A = 8'hA; B = 8'hF; #100;
A = 8'hA; B = 8'h10; #100;
A = 8'hA; B = 8'h11; #100;
A = 8'hA; B = 8'h12; #100;
A = 8'hA; B = 8'h13; #100;
A = 8'hA; B = 8'h14; #100;
A = 8'hA; B = 8'h15; #100;
A = 8'hA; B = 8'h16; #100;
A = 8'hA; B = 8'h17; #100;
A = 8'hA; B = 8'h18; #100;
A = 8'hA; B = 8'h19; #100;
A = 8'hA; B = 8'h1A; #100;
A = 8'hA; B = 8'h1B; #100;
A = 8'hA; B = 8'h1C; #100;
A = 8'hA; B = 8'h1D; #100;
A = 8'hA; B = 8'h1E; #100;
A = 8'hA; B = 8'h1F; #100;
A = 8'hA; B = 8'h20; #100;
A = 8'hA; B = 8'h21; #100;
A = 8'hA; B = 8'h22; #100;
A = 8'hA; B = 8'h23; #100;
A = 8'hA; B = 8'h24; #100;
A = 8'hA; B = 8'h25; #100;
A = 8'hA; B = 8'h26; #100;
A = 8'hA; B = 8'h27; #100;
A = 8'hA; B = 8'h28; #100;
A = 8'hA; B = 8'h29; #100;
A = 8'hA; B = 8'h2A; #100;
A = 8'hA; B = 8'h2B; #100;
A = 8'hA; B = 8'h2C; #100;
A = 8'hA; B = 8'h2D; #100;
A = 8'hA; B = 8'h2E; #100;
A = 8'hA; B = 8'h2F; #100;
A = 8'hA; B = 8'h30; #100;
A = 8'hA; B = 8'h31; #100;
A = 8'hA; B = 8'h32; #100;
A = 8'hA; B = 8'h33; #100;
A = 8'hA; B = 8'h34; #100;
A = 8'hA; B = 8'h35; #100;
A = 8'hA; B = 8'h36; #100;
A = 8'hA; B = 8'h37; #100;
A = 8'hA; B = 8'h38; #100;
A = 8'hA; B = 8'h39; #100;
A = 8'hA; B = 8'h3A; #100;
A = 8'hA; B = 8'h3B; #100;
A = 8'hA; B = 8'h3C; #100;
A = 8'hA; B = 8'h3D; #100;
A = 8'hA; B = 8'h3E; #100;
A = 8'hA; B = 8'h3F; #100;
A = 8'hA; B = 8'h40; #100;
A = 8'hA; B = 8'h41; #100;
A = 8'hA; B = 8'h42; #100;
A = 8'hA; B = 8'h43; #100;
A = 8'hA; B = 8'h44; #100;
A = 8'hA; B = 8'h45; #100;
A = 8'hA; B = 8'h46; #100;
A = 8'hA; B = 8'h47; #100;
A = 8'hA; B = 8'h48; #100;
A = 8'hA; B = 8'h49; #100;
A = 8'hA; B = 8'h4A; #100;
A = 8'hA; B = 8'h4B; #100;
A = 8'hA; B = 8'h4C; #100;
A = 8'hA; B = 8'h4D; #100;
A = 8'hA; B = 8'h4E; #100;
A = 8'hA; B = 8'h4F; #100;
A = 8'hA; B = 8'h50; #100;
A = 8'hA; B = 8'h51; #100;
A = 8'hA; B = 8'h52; #100;
A = 8'hA; B = 8'h53; #100;
A = 8'hA; B = 8'h54; #100;
A = 8'hA; B = 8'h55; #100;
A = 8'hA; B = 8'h56; #100;
A = 8'hA; B = 8'h57; #100;
A = 8'hA; B = 8'h58; #100;
A = 8'hA; B = 8'h59; #100;
A = 8'hA; B = 8'h5A; #100;
A = 8'hA; B = 8'h5B; #100;
A = 8'hA; B = 8'h5C; #100;
A = 8'hA; B = 8'h5D; #100;
A = 8'hA; B = 8'h5E; #100;
A = 8'hA; B = 8'h5F; #100;
A = 8'hA; B = 8'h60; #100;
A = 8'hA; B = 8'h61; #100;
A = 8'hA; B = 8'h62; #100;
A = 8'hA; B = 8'h63; #100;
A = 8'hA; B = 8'h64; #100;
A = 8'hA; B = 8'h65; #100;
A = 8'hA; B = 8'h66; #100;
A = 8'hA; B = 8'h67; #100;
A = 8'hA; B = 8'h68; #100;
A = 8'hA; B = 8'h69; #100;
A = 8'hA; B = 8'h6A; #100;
A = 8'hA; B = 8'h6B; #100;
A = 8'hA; B = 8'h6C; #100;
A = 8'hA; B = 8'h6D; #100;
A = 8'hA; B = 8'h6E; #100;
A = 8'hA; B = 8'h6F; #100;
A = 8'hA; B = 8'h70; #100;
A = 8'hA; B = 8'h71; #100;
A = 8'hA; B = 8'h72; #100;
A = 8'hA; B = 8'h73; #100;
A = 8'hA; B = 8'h74; #100;
A = 8'hA; B = 8'h75; #100;
A = 8'hA; B = 8'h76; #100;
A = 8'hA; B = 8'h77; #100;
A = 8'hA; B = 8'h78; #100;
A = 8'hA; B = 8'h79; #100;
A = 8'hA; B = 8'h7A; #100;
A = 8'hA; B = 8'h7B; #100;
A = 8'hA; B = 8'h7C; #100;
A = 8'hA; B = 8'h7D; #100;
A = 8'hA; B = 8'h7E; #100;
A = 8'hA; B = 8'h7F; #100;
A = 8'hA; B = 8'h80; #100;
A = 8'hA; B = 8'h81; #100;
A = 8'hA; B = 8'h82; #100;
A = 8'hA; B = 8'h83; #100;
A = 8'hA; B = 8'h84; #100;
A = 8'hA; B = 8'h85; #100;
A = 8'hA; B = 8'h86; #100;
A = 8'hA; B = 8'h87; #100;
A = 8'hA; B = 8'h88; #100;
A = 8'hA; B = 8'h89; #100;
A = 8'hA; B = 8'h8A; #100;
A = 8'hA; B = 8'h8B; #100;
A = 8'hA; B = 8'h8C; #100;
A = 8'hA; B = 8'h8D; #100;
A = 8'hA; B = 8'h8E; #100;
A = 8'hA; B = 8'h8F; #100;
A = 8'hA; B = 8'h90; #100;
A = 8'hA; B = 8'h91; #100;
A = 8'hA; B = 8'h92; #100;
A = 8'hA; B = 8'h93; #100;
A = 8'hA; B = 8'h94; #100;
A = 8'hA; B = 8'h95; #100;
A = 8'hA; B = 8'h96; #100;
A = 8'hA; B = 8'h97; #100;
A = 8'hA; B = 8'h98; #100;
A = 8'hA; B = 8'h99; #100;
A = 8'hA; B = 8'h9A; #100;
A = 8'hA; B = 8'h9B; #100;
A = 8'hA; B = 8'h9C; #100;
A = 8'hA; B = 8'h9D; #100;
A = 8'hA; B = 8'h9E; #100;
A = 8'hA; B = 8'h9F; #100;
A = 8'hA; B = 8'hA0; #100;
A = 8'hA; B = 8'hA1; #100;
A = 8'hA; B = 8'hA2; #100;
A = 8'hA; B = 8'hA3; #100;
A = 8'hA; B = 8'hA4; #100;
A = 8'hA; B = 8'hA5; #100;
A = 8'hA; B = 8'hA6; #100;
A = 8'hA; B = 8'hA7; #100;
A = 8'hA; B = 8'hA8; #100;
A = 8'hA; B = 8'hA9; #100;
A = 8'hA; B = 8'hAA; #100;
A = 8'hA; B = 8'hAB; #100;
A = 8'hA; B = 8'hAC; #100;
A = 8'hA; B = 8'hAD; #100;
A = 8'hA; B = 8'hAE; #100;
A = 8'hA; B = 8'hAF; #100;
A = 8'hA; B = 8'hB0; #100;
A = 8'hA; B = 8'hB1; #100;
A = 8'hA; B = 8'hB2; #100;
A = 8'hA; B = 8'hB3; #100;
A = 8'hA; B = 8'hB4; #100;
A = 8'hA; B = 8'hB5; #100;
A = 8'hA; B = 8'hB6; #100;
A = 8'hA; B = 8'hB7; #100;
A = 8'hA; B = 8'hB8; #100;
A = 8'hA; B = 8'hB9; #100;
A = 8'hA; B = 8'hBA; #100;
A = 8'hA; B = 8'hBB; #100;
A = 8'hA; B = 8'hBC; #100;
A = 8'hA; B = 8'hBD; #100;
A = 8'hA; B = 8'hBE; #100;
A = 8'hA; B = 8'hBF; #100;
A = 8'hA; B = 8'hC0; #100;
A = 8'hA; B = 8'hC1; #100;
A = 8'hA; B = 8'hC2; #100;
A = 8'hA; B = 8'hC3; #100;
A = 8'hA; B = 8'hC4; #100;
A = 8'hA; B = 8'hC5; #100;
A = 8'hA; B = 8'hC6; #100;
A = 8'hA; B = 8'hC7; #100;
A = 8'hA; B = 8'hC8; #100;
A = 8'hA; B = 8'hC9; #100;
A = 8'hA; B = 8'hCA; #100;
A = 8'hA; B = 8'hCB; #100;
A = 8'hA; B = 8'hCC; #100;
A = 8'hA; B = 8'hCD; #100;
A = 8'hA; B = 8'hCE; #100;
A = 8'hA; B = 8'hCF; #100;
A = 8'hA; B = 8'hD0; #100;
A = 8'hA; B = 8'hD1; #100;
A = 8'hA; B = 8'hD2; #100;
A = 8'hA; B = 8'hD3; #100;
A = 8'hA; B = 8'hD4; #100;
A = 8'hA; B = 8'hD5; #100;
A = 8'hA; B = 8'hD6; #100;
A = 8'hA; B = 8'hD7; #100;
A = 8'hA; B = 8'hD8; #100;
A = 8'hA; B = 8'hD9; #100;
A = 8'hA; B = 8'hDA; #100;
A = 8'hA; B = 8'hDB; #100;
A = 8'hA; B = 8'hDC; #100;
A = 8'hA; B = 8'hDD; #100;
A = 8'hA; B = 8'hDE; #100;
A = 8'hA; B = 8'hDF; #100;
A = 8'hA; B = 8'hE0; #100;
A = 8'hA; B = 8'hE1; #100;
A = 8'hA; B = 8'hE2; #100;
A = 8'hA; B = 8'hE3; #100;
A = 8'hA; B = 8'hE4; #100;
A = 8'hA; B = 8'hE5; #100;
A = 8'hA; B = 8'hE6; #100;
A = 8'hA; B = 8'hE7; #100;
A = 8'hA; B = 8'hE8; #100;
A = 8'hA; B = 8'hE9; #100;
A = 8'hA; B = 8'hEA; #100;
A = 8'hA; B = 8'hEB; #100;
A = 8'hA; B = 8'hEC; #100;
A = 8'hA; B = 8'hED; #100;
A = 8'hA; B = 8'hEE; #100;
A = 8'hA; B = 8'hEF; #100;
A = 8'hA; B = 8'hF0; #100;
A = 8'hA; B = 8'hF1; #100;
A = 8'hA; B = 8'hF2; #100;
A = 8'hA; B = 8'hF3; #100;
A = 8'hA; B = 8'hF4; #100;
A = 8'hA; B = 8'hF5; #100;
A = 8'hA; B = 8'hF6; #100;
A = 8'hA; B = 8'hF7; #100;
A = 8'hA; B = 8'hF8; #100;
A = 8'hA; B = 8'hF9; #100;
A = 8'hA; B = 8'hFA; #100;
A = 8'hA; B = 8'hFB; #100;
A = 8'hA; B = 8'hFC; #100;
A = 8'hA; B = 8'hFD; #100;
A = 8'hA; B = 8'hFE; #100;
A = 8'hA; B = 8'hFF; #100;
A = 8'hB; B = 8'h0; #100;
A = 8'hB; B = 8'h1; #100;
A = 8'hB; B = 8'h2; #100;
A = 8'hB; B = 8'h3; #100;
A = 8'hB; B = 8'h4; #100;
A = 8'hB; B = 8'h5; #100;
A = 8'hB; B = 8'h6; #100;
A = 8'hB; B = 8'h7; #100;
A = 8'hB; B = 8'h8; #100;
A = 8'hB; B = 8'h9; #100;
A = 8'hB; B = 8'hA; #100;
A = 8'hB; B = 8'hB; #100;
A = 8'hB; B = 8'hC; #100;
A = 8'hB; B = 8'hD; #100;
A = 8'hB; B = 8'hE; #100;
A = 8'hB; B = 8'hF; #100;
A = 8'hB; B = 8'h10; #100;
A = 8'hB; B = 8'h11; #100;
A = 8'hB; B = 8'h12; #100;
A = 8'hB; B = 8'h13; #100;
A = 8'hB; B = 8'h14; #100;
A = 8'hB; B = 8'h15; #100;
A = 8'hB; B = 8'h16; #100;
A = 8'hB; B = 8'h17; #100;
A = 8'hB; B = 8'h18; #100;
A = 8'hB; B = 8'h19; #100;
A = 8'hB; B = 8'h1A; #100;
A = 8'hB; B = 8'h1B; #100;
A = 8'hB; B = 8'h1C; #100;
A = 8'hB; B = 8'h1D; #100;
A = 8'hB; B = 8'h1E; #100;
A = 8'hB; B = 8'h1F; #100;
A = 8'hB; B = 8'h20; #100;
A = 8'hB; B = 8'h21; #100;
A = 8'hB; B = 8'h22; #100;
A = 8'hB; B = 8'h23; #100;
A = 8'hB; B = 8'h24; #100;
A = 8'hB; B = 8'h25; #100;
A = 8'hB; B = 8'h26; #100;
A = 8'hB; B = 8'h27; #100;
A = 8'hB; B = 8'h28; #100;
A = 8'hB; B = 8'h29; #100;
A = 8'hB; B = 8'h2A; #100;
A = 8'hB; B = 8'h2B; #100;
A = 8'hB; B = 8'h2C; #100;
A = 8'hB; B = 8'h2D; #100;
A = 8'hB; B = 8'h2E; #100;
A = 8'hB; B = 8'h2F; #100;
A = 8'hB; B = 8'h30; #100;
A = 8'hB; B = 8'h31; #100;
A = 8'hB; B = 8'h32; #100;
A = 8'hB; B = 8'h33; #100;
A = 8'hB; B = 8'h34; #100;
A = 8'hB; B = 8'h35; #100;
A = 8'hB; B = 8'h36; #100;
A = 8'hB; B = 8'h37; #100;
A = 8'hB; B = 8'h38; #100;
A = 8'hB; B = 8'h39; #100;
A = 8'hB; B = 8'h3A; #100;
A = 8'hB; B = 8'h3B; #100;
A = 8'hB; B = 8'h3C; #100;
A = 8'hB; B = 8'h3D; #100;
A = 8'hB; B = 8'h3E; #100;
A = 8'hB; B = 8'h3F; #100;
A = 8'hB; B = 8'h40; #100;
A = 8'hB; B = 8'h41; #100;
A = 8'hB; B = 8'h42; #100;
A = 8'hB; B = 8'h43; #100;
A = 8'hB; B = 8'h44; #100;
A = 8'hB; B = 8'h45; #100;
A = 8'hB; B = 8'h46; #100;
A = 8'hB; B = 8'h47; #100;
A = 8'hB; B = 8'h48; #100;
A = 8'hB; B = 8'h49; #100;
A = 8'hB; B = 8'h4A; #100;
A = 8'hB; B = 8'h4B; #100;
A = 8'hB; B = 8'h4C; #100;
A = 8'hB; B = 8'h4D; #100;
A = 8'hB; B = 8'h4E; #100;
A = 8'hB; B = 8'h4F; #100;
A = 8'hB; B = 8'h50; #100;
A = 8'hB; B = 8'h51; #100;
A = 8'hB; B = 8'h52; #100;
A = 8'hB; B = 8'h53; #100;
A = 8'hB; B = 8'h54; #100;
A = 8'hB; B = 8'h55; #100;
A = 8'hB; B = 8'h56; #100;
A = 8'hB; B = 8'h57; #100;
A = 8'hB; B = 8'h58; #100;
A = 8'hB; B = 8'h59; #100;
A = 8'hB; B = 8'h5A; #100;
A = 8'hB; B = 8'h5B; #100;
A = 8'hB; B = 8'h5C; #100;
A = 8'hB; B = 8'h5D; #100;
A = 8'hB; B = 8'h5E; #100;
A = 8'hB; B = 8'h5F; #100;
A = 8'hB; B = 8'h60; #100;
A = 8'hB; B = 8'h61; #100;
A = 8'hB; B = 8'h62; #100;
A = 8'hB; B = 8'h63; #100;
A = 8'hB; B = 8'h64; #100;
A = 8'hB; B = 8'h65; #100;
A = 8'hB; B = 8'h66; #100;
A = 8'hB; B = 8'h67; #100;
A = 8'hB; B = 8'h68; #100;
A = 8'hB; B = 8'h69; #100;
A = 8'hB; B = 8'h6A; #100;
A = 8'hB; B = 8'h6B; #100;
A = 8'hB; B = 8'h6C; #100;
A = 8'hB; B = 8'h6D; #100;
A = 8'hB; B = 8'h6E; #100;
A = 8'hB; B = 8'h6F; #100;
A = 8'hB; B = 8'h70; #100;
A = 8'hB; B = 8'h71; #100;
A = 8'hB; B = 8'h72; #100;
A = 8'hB; B = 8'h73; #100;
A = 8'hB; B = 8'h74; #100;
A = 8'hB; B = 8'h75; #100;
A = 8'hB; B = 8'h76; #100;
A = 8'hB; B = 8'h77; #100;
A = 8'hB; B = 8'h78; #100;
A = 8'hB; B = 8'h79; #100;
A = 8'hB; B = 8'h7A; #100;
A = 8'hB; B = 8'h7B; #100;
A = 8'hB; B = 8'h7C; #100;
A = 8'hB; B = 8'h7D; #100;
A = 8'hB; B = 8'h7E; #100;
A = 8'hB; B = 8'h7F; #100;
A = 8'hB; B = 8'h80; #100;
A = 8'hB; B = 8'h81; #100;
A = 8'hB; B = 8'h82; #100;
A = 8'hB; B = 8'h83; #100;
A = 8'hB; B = 8'h84; #100;
A = 8'hB; B = 8'h85; #100;
A = 8'hB; B = 8'h86; #100;
A = 8'hB; B = 8'h87; #100;
A = 8'hB; B = 8'h88; #100;
A = 8'hB; B = 8'h89; #100;
A = 8'hB; B = 8'h8A; #100;
A = 8'hB; B = 8'h8B; #100;
A = 8'hB; B = 8'h8C; #100;
A = 8'hB; B = 8'h8D; #100;
A = 8'hB; B = 8'h8E; #100;
A = 8'hB; B = 8'h8F; #100;
A = 8'hB; B = 8'h90; #100;
A = 8'hB; B = 8'h91; #100;
A = 8'hB; B = 8'h92; #100;
A = 8'hB; B = 8'h93; #100;
A = 8'hB; B = 8'h94; #100;
A = 8'hB; B = 8'h95; #100;
A = 8'hB; B = 8'h96; #100;
A = 8'hB; B = 8'h97; #100;
A = 8'hB; B = 8'h98; #100;
A = 8'hB; B = 8'h99; #100;
A = 8'hB; B = 8'h9A; #100;
A = 8'hB; B = 8'h9B; #100;
A = 8'hB; B = 8'h9C; #100;
A = 8'hB; B = 8'h9D; #100;
A = 8'hB; B = 8'h9E; #100;
A = 8'hB; B = 8'h9F; #100;
A = 8'hB; B = 8'hA0; #100;
A = 8'hB; B = 8'hA1; #100;
A = 8'hB; B = 8'hA2; #100;
A = 8'hB; B = 8'hA3; #100;
A = 8'hB; B = 8'hA4; #100;
A = 8'hB; B = 8'hA5; #100;
A = 8'hB; B = 8'hA6; #100;
A = 8'hB; B = 8'hA7; #100;
A = 8'hB; B = 8'hA8; #100;
A = 8'hB; B = 8'hA9; #100;
A = 8'hB; B = 8'hAA; #100;
A = 8'hB; B = 8'hAB; #100;
A = 8'hB; B = 8'hAC; #100;
A = 8'hB; B = 8'hAD; #100;
A = 8'hB; B = 8'hAE; #100;
A = 8'hB; B = 8'hAF; #100;
A = 8'hB; B = 8'hB0; #100;
A = 8'hB; B = 8'hB1; #100;
A = 8'hB; B = 8'hB2; #100;
A = 8'hB; B = 8'hB3; #100;
A = 8'hB; B = 8'hB4; #100;
A = 8'hB; B = 8'hB5; #100;
A = 8'hB; B = 8'hB6; #100;
A = 8'hB; B = 8'hB7; #100;
A = 8'hB; B = 8'hB8; #100;
A = 8'hB; B = 8'hB9; #100;
A = 8'hB; B = 8'hBA; #100;
A = 8'hB; B = 8'hBB; #100;
A = 8'hB; B = 8'hBC; #100;
A = 8'hB; B = 8'hBD; #100;
A = 8'hB; B = 8'hBE; #100;
A = 8'hB; B = 8'hBF; #100;
A = 8'hB; B = 8'hC0; #100;
A = 8'hB; B = 8'hC1; #100;
A = 8'hB; B = 8'hC2; #100;
A = 8'hB; B = 8'hC3; #100;
A = 8'hB; B = 8'hC4; #100;
A = 8'hB; B = 8'hC5; #100;
A = 8'hB; B = 8'hC6; #100;
A = 8'hB; B = 8'hC7; #100;
A = 8'hB; B = 8'hC8; #100;
A = 8'hB; B = 8'hC9; #100;
A = 8'hB; B = 8'hCA; #100;
A = 8'hB; B = 8'hCB; #100;
A = 8'hB; B = 8'hCC; #100;
A = 8'hB; B = 8'hCD; #100;
A = 8'hB; B = 8'hCE; #100;
A = 8'hB; B = 8'hCF; #100;
A = 8'hB; B = 8'hD0; #100;
A = 8'hB; B = 8'hD1; #100;
A = 8'hB; B = 8'hD2; #100;
A = 8'hB; B = 8'hD3; #100;
A = 8'hB; B = 8'hD4; #100;
A = 8'hB; B = 8'hD5; #100;
A = 8'hB; B = 8'hD6; #100;
A = 8'hB; B = 8'hD7; #100;
A = 8'hB; B = 8'hD8; #100;
A = 8'hB; B = 8'hD9; #100;
A = 8'hB; B = 8'hDA; #100;
A = 8'hB; B = 8'hDB; #100;
A = 8'hB; B = 8'hDC; #100;
A = 8'hB; B = 8'hDD; #100;
A = 8'hB; B = 8'hDE; #100;
A = 8'hB; B = 8'hDF; #100;
A = 8'hB; B = 8'hE0; #100;
A = 8'hB; B = 8'hE1; #100;
A = 8'hB; B = 8'hE2; #100;
A = 8'hB; B = 8'hE3; #100;
A = 8'hB; B = 8'hE4; #100;
A = 8'hB; B = 8'hE5; #100;
A = 8'hB; B = 8'hE6; #100;
A = 8'hB; B = 8'hE7; #100;
A = 8'hB; B = 8'hE8; #100;
A = 8'hB; B = 8'hE9; #100;
A = 8'hB; B = 8'hEA; #100;
A = 8'hB; B = 8'hEB; #100;
A = 8'hB; B = 8'hEC; #100;
A = 8'hB; B = 8'hED; #100;
A = 8'hB; B = 8'hEE; #100;
A = 8'hB; B = 8'hEF; #100;
A = 8'hB; B = 8'hF0; #100;
A = 8'hB; B = 8'hF1; #100;
A = 8'hB; B = 8'hF2; #100;
A = 8'hB; B = 8'hF3; #100;
A = 8'hB; B = 8'hF4; #100;
A = 8'hB; B = 8'hF5; #100;
A = 8'hB; B = 8'hF6; #100;
A = 8'hB; B = 8'hF7; #100;
A = 8'hB; B = 8'hF8; #100;
A = 8'hB; B = 8'hF9; #100;
A = 8'hB; B = 8'hFA; #100;
A = 8'hB; B = 8'hFB; #100;
A = 8'hB; B = 8'hFC; #100;
A = 8'hB; B = 8'hFD; #100;
A = 8'hB; B = 8'hFE; #100;
A = 8'hB; B = 8'hFF; #100;
A = 8'hC; B = 8'h0; #100;
A = 8'hC; B = 8'h1; #100;
A = 8'hC; B = 8'h2; #100;
A = 8'hC; B = 8'h3; #100;
A = 8'hC; B = 8'h4; #100;
A = 8'hC; B = 8'h5; #100;
A = 8'hC; B = 8'h6; #100;
A = 8'hC; B = 8'h7; #100;
A = 8'hC; B = 8'h8; #100;
A = 8'hC; B = 8'h9; #100;
A = 8'hC; B = 8'hA; #100;
A = 8'hC; B = 8'hB; #100;
A = 8'hC; B = 8'hC; #100;
A = 8'hC; B = 8'hD; #100;
A = 8'hC; B = 8'hE; #100;
A = 8'hC; B = 8'hF; #100;
A = 8'hC; B = 8'h10; #100;
A = 8'hC; B = 8'h11; #100;
A = 8'hC; B = 8'h12; #100;
A = 8'hC; B = 8'h13; #100;
A = 8'hC; B = 8'h14; #100;
A = 8'hC; B = 8'h15; #100;
A = 8'hC; B = 8'h16; #100;
A = 8'hC; B = 8'h17; #100;
A = 8'hC; B = 8'h18; #100;
A = 8'hC; B = 8'h19; #100;
A = 8'hC; B = 8'h1A; #100;
A = 8'hC; B = 8'h1B; #100;
A = 8'hC; B = 8'h1C; #100;
A = 8'hC; B = 8'h1D; #100;
A = 8'hC; B = 8'h1E; #100;
A = 8'hC; B = 8'h1F; #100;
A = 8'hC; B = 8'h20; #100;
A = 8'hC; B = 8'h21; #100;
A = 8'hC; B = 8'h22; #100;
A = 8'hC; B = 8'h23; #100;
A = 8'hC; B = 8'h24; #100;
A = 8'hC; B = 8'h25; #100;
A = 8'hC; B = 8'h26; #100;
A = 8'hC; B = 8'h27; #100;
A = 8'hC; B = 8'h28; #100;
A = 8'hC; B = 8'h29; #100;
A = 8'hC; B = 8'h2A; #100;
A = 8'hC; B = 8'h2B; #100;
A = 8'hC; B = 8'h2C; #100;
A = 8'hC; B = 8'h2D; #100;
A = 8'hC; B = 8'h2E; #100;
A = 8'hC; B = 8'h2F; #100;
A = 8'hC; B = 8'h30; #100;
A = 8'hC; B = 8'h31; #100;
A = 8'hC; B = 8'h32; #100;
A = 8'hC; B = 8'h33; #100;
A = 8'hC; B = 8'h34; #100;
A = 8'hC; B = 8'h35; #100;
A = 8'hC; B = 8'h36; #100;
A = 8'hC; B = 8'h37; #100;
A = 8'hC; B = 8'h38; #100;
A = 8'hC; B = 8'h39; #100;
A = 8'hC; B = 8'h3A; #100;
A = 8'hC; B = 8'h3B; #100;
A = 8'hC; B = 8'h3C; #100;
A = 8'hC; B = 8'h3D; #100;
A = 8'hC; B = 8'h3E; #100;
A = 8'hC; B = 8'h3F; #100;
A = 8'hC; B = 8'h40; #100;
A = 8'hC; B = 8'h41; #100;
A = 8'hC; B = 8'h42; #100;
A = 8'hC; B = 8'h43; #100;
A = 8'hC; B = 8'h44; #100;
A = 8'hC; B = 8'h45; #100;
A = 8'hC; B = 8'h46; #100;
A = 8'hC; B = 8'h47; #100;
A = 8'hC; B = 8'h48; #100;
A = 8'hC; B = 8'h49; #100;
A = 8'hC; B = 8'h4A; #100;
A = 8'hC; B = 8'h4B; #100;
A = 8'hC; B = 8'h4C; #100;
A = 8'hC; B = 8'h4D; #100;
A = 8'hC; B = 8'h4E; #100;
A = 8'hC; B = 8'h4F; #100;
A = 8'hC; B = 8'h50; #100;
A = 8'hC; B = 8'h51; #100;
A = 8'hC; B = 8'h52; #100;
A = 8'hC; B = 8'h53; #100;
A = 8'hC; B = 8'h54; #100;
A = 8'hC; B = 8'h55; #100;
A = 8'hC; B = 8'h56; #100;
A = 8'hC; B = 8'h57; #100;
A = 8'hC; B = 8'h58; #100;
A = 8'hC; B = 8'h59; #100;
A = 8'hC; B = 8'h5A; #100;
A = 8'hC; B = 8'h5B; #100;
A = 8'hC; B = 8'h5C; #100;
A = 8'hC; B = 8'h5D; #100;
A = 8'hC; B = 8'h5E; #100;
A = 8'hC; B = 8'h5F; #100;
A = 8'hC; B = 8'h60; #100;
A = 8'hC; B = 8'h61; #100;
A = 8'hC; B = 8'h62; #100;
A = 8'hC; B = 8'h63; #100;
A = 8'hC; B = 8'h64; #100;
A = 8'hC; B = 8'h65; #100;
A = 8'hC; B = 8'h66; #100;
A = 8'hC; B = 8'h67; #100;
A = 8'hC; B = 8'h68; #100;
A = 8'hC; B = 8'h69; #100;
A = 8'hC; B = 8'h6A; #100;
A = 8'hC; B = 8'h6B; #100;
A = 8'hC; B = 8'h6C; #100;
A = 8'hC; B = 8'h6D; #100;
A = 8'hC; B = 8'h6E; #100;
A = 8'hC; B = 8'h6F; #100;
A = 8'hC; B = 8'h70; #100;
A = 8'hC; B = 8'h71; #100;
A = 8'hC; B = 8'h72; #100;
A = 8'hC; B = 8'h73; #100;
A = 8'hC; B = 8'h74; #100;
A = 8'hC; B = 8'h75; #100;
A = 8'hC; B = 8'h76; #100;
A = 8'hC; B = 8'h77; #100;
A = 8'hC; B = 8'h78; #100;
A = 8'hC; B = 8'h79; #100;
A = 8'hC; B = 8'h7A; #100;
A = 8'hC; B = 8'h7B; #100;
A = 8'hC; B = 8'h7C; #100;
A = 8'hC; B = 8'h7D; #100;
A = 8'hC; B = 8'h7E; #100;
A = 8'hC; B = 8'h7F; #100;
A = 8'hC; B = 8'h80; #100;
A = 8'hC; B = 8'h81; #100;
A = 8'hC; B = 8'h82; #100;
A = 8'hC; B = 8'h83; #100;
A = 8'hC; B = 8'h84; #100;
A = 8'hC; B = 8'h85; #100;
A = 8'hC; B = 8'h86; #100;
A = 8'hC; B = 8'h87; #100;
A = 8'hC; B = 8'h88; #100;
A = 8'hC; B = 8'h89; #100;
A = 8'hC; B = 8'h8A; #100;
A = 8'hC; B = 8'h8B; #100;
A = 8'hC; B = 8'h8C; #100;
A = 8'hC; B = 8'h8D; #100;
A = 8'hC; B = 8'h8E; #100;
A = 8'hC; B = 8'h8F; #100;
A = 8'hC; B = 8'h90; #100;
A = 8'hC; B = 8'h91; #100;
A = 8'hC; B = 8'h92; #100;
A = 8'hC; B = 8'h93; #100;
A = 8'hC; B = 8'h94; #100;
A = 8'hC; B = 8'h95; #100;
A = 8'hC; B = 8'h96; #100;
A = 8'hC; B = 8'h97; #100;
A = 8'hC; B = 8'h98; #100;
A = 8'hC; B = 8'h99; #100;
A = 8'hC; B = 8'h9A; #100;
A = 8'hC; B = 8'h9B; #100;
A = 8'hC; B = 8'h9C; #100;
A = 8'hC; B = 8'h9D; #100;
A = 8'hC; B = 8'h9E; #100;
A = 8'hC; B = 8'h9F; #100;
A = 8'hC; B = 8'hA0; #100;
A = 8'hC; B = 8'hA1; #100;
A = 8'hC; B = 8'hA2; #100;
A = 8'hC; B = 8'hA3; #100;
A = 8'hC; B = 8'hA4; #100;
A = 8'hC; B = 8'hA5; #100;
A = 8'hC; B = 8'hA6; #100;
A = 8'hC; B = 8'hA7; #100;
A = 8'hC; B = 8'hA8; #100;
A = 8'hC; B = 8'hA9; #100;
A = 8'hC; B = 8'hAA; #100;
A = 8'hC; B = 8'hAB; #100;
A = 8'hC; B = 8'hAC; #100;
A = 8'hC; B = 8'hAD; #100;
A = 8'hC; B = 8'hAE; #100;
A = 8'hC; B = 8'hAF; #100;
A = 8'hC; B = 8'hB0; #100;
A = 8'hC; B = 8'hB1; #100;
A = 8'hC; B = 8'hB2; #100;
A = 8'hC; B = 8'hB3; #100;
A = 8'hC; B = 8'hB4; #100;
A = 8'hC; B = 8'hB5; #100;
A = 8'hC; B = 8'hB6; #100;
A = 8'hC; B = 8'hB7; #100;
A = 8'hC; B = 8'hB8; #100;
A = 8'hC; B = 8'hB9; #100;
A = 8'hC; B = 8'hBA; #100;
A = 8'hC; B = 8'hBB; #100;
A = 8'hC; B = 8'hBC; #100;
A = 8'hC; B = 8'hBD; #100;
A = 8'hC; B = 8'hBE; #100;
A = 8'hC; B = 8'hBF; #100;
A = 8'hC; B = 8'hC0; #100;
A = 8'hC; B = 8'hC1; #100;
A = 8'hC; B = 8'hC2; #100;
A = 8'hC; B = 8'hC3; #100;
A = 8'hC; B = 8'hC4; #100;
A = 8'hC; B = 8'hC5; #100;
A = 8'hC; B = 8'hC6; #100;
A = 8'hC; B = 8'hC7; #100;
A = 8'hC; B = 8'hC8; #100;
A = 8'hC; B = 8'hC9; #100;
A = 8'hC; B = 8'hCA; #100;
A = 8'hC; B = 8'hCB; #100;
A = 8'hC; B = 8'hCC; #100;
A = 8'hC; B = 8'hCD; #100;
A = 8'hC; B = 8'hCE; #100;
A = 8'hC; B = 8'hCF; #100;
A = 8'hC; B = 8'hD0; #100;
A = 8'hC; B = 8'hD1; #100;
A = 8'hC; B = 8'hD2; #100;
A = 8'hC; B = 8'hD3; #100;
A = 8'hC; B = 8'hD4; #100;
A = 8'hC; B = 8'hD5; #100;
A = 8'hC; B = 8'hD6; #100;
A = 8'hC; B = 8'hD7; #100;
A = 8'hC; B = 8'hD8; #100;
A = 8'hC; B = 8'hD9; #100;
A = 8'hC; B = 8'hDA; #100;
A = 8'hC; B = 8'hDB; #100;
A = 8'hC; B = 8'hDC; #100;
A = 8'hC; B = 8'hDD; #100;
A = 8'hC; B = 8'hDE; #100;
A = 8'hC; B = 8'hDF; #100;
A = 8'hC; B = 8'hE0; #100;
A = 8'hC; B = 8'hE1; #100;
A = 8'hC; B = 8'hE2; #100;
A = 8'hC; B = 8'hE3; #100;
A = 8'hC; B = 8'hE4; #100;
A = 8'hC; B = 8'hE5; #100;
A = 8'hC; B = 8'hE6; #100;
A = 8'hC; B = 8'hE7; #100;
A = 8'hC; B = 8'hE8; #100;
A = 8'hC; B = 8'hE9; #100;
A = 8'hC; B = 8'hEA; #100;
A = 8'hC; B = 8'hEB; #100;
A = 8'hC; B = 8'hEC; #100;
A = 8'hC; B = 8'hED; #100;
A = 8'hC; B = 8'hEE; #100;
A = 8'hC; B = 8'hEF; #100;
A = 8'hC; B = 8'hF0; #100;
A = 8'hC; B = 8'hF1; #100;
A = 8'hC; B = 8'hF2; #100;
A = 8'hC; B = 8'hF3; #100;
A = 8'hC; B = 8'hF4; #100;
A = 8'hC; B = 8'hF5; #100;
A = 8'hC; B = 8'hF6; #100;
A = 8'hC; B = 8'hF7; #100;
A = 8'hC; B = 8'hF8; #100;
A = 8'hC; B = 8'hF9; #100;
A = 8'hC; B = 8'hFA; #100;
A = 8'hC; B = 8'hFB; #100;
A = 8'hC; B = 8'hFC; #100;
A = 8'hC; B = 8'hFD; #100;
A = 8'hC; B = 8'hFE; #100;
A = 8'hC; B = 8'hFF; #100;
A = 8'hD; B = 8'h0; #100;
A = 8'hD; B = 8'h1; #100;
A = 8'hD; B = 8'h2; #100;
A = 8'hD; B = 8'h3; #100;
A = 8'hD; B = 8'h4; #100;
A = 8'hD; B = 8'h5; #100;
A = 8'hD; B = 8'h6; #100;
A = 8'hD; B = 8'h7; #100;
A = 8'hD; B = 8'h8; #100;
A = 8'hD; B = 8'h9; #100;
A = 8'hD; B = 8'hA; #100;
A = 8'hD; B = 8'hB; #100;
A = 8'hD; B = 8'hC; #100;
A = 8'hD; B = 8'hD; #100;
A = 8'hD; B = 8'hE; #100;
A = 8'hD; B = 8'hF; #100;
A = 8'hD; B = 8'h10; #100;
A = 8'hD; B = 8'h11; #100;
A = 8'hD; B = 8'h12; #100;
A = 8'hD; B = 8'h13; #100;
A = 8'hD; B = 8'h14; #100;
A = 8'hD; B = 8'h15; #100;
A = 8'hD; B = 8'h16; #100;
A = 8'hD; B = 8'h17; #100;
A = 8'hD; B = 8'h18; #100;
A = 8'hD; B = 8'h19; #100;
A = 8'hD; B = 8'h1A; #100;
A = 8'hD; B = 8'h1B; #100;
A = 8'hD; B = 8'h1C; #100;
A = 8'hD; B = 8'h1D; #100;
A = 8'hD; B = 8'h1E; #100;
A = 8'hD; B = 8'h1F; #100;
A = 8'hD; B = 8'h20; #100;
A = 8'hD; B = 8'h21; #100;
A = 8'hD; B = 8'h22; #100;
A = 8'hD; B = 8'h23; #100;
A = 8'hD; B = 8'h24; #100;
A = 8'hD; B = 8'h25; #100;
A = 8'hD; B = 8'h26; #100;
A = 8'hD; B = 8'h27; #100;
A = 8'hD; B = 8'h28; #100;
A = 8'hD; B = 8'h29; #100;
A = 8'hD; B = 8'h2A; #100;
A = 8'hD; B = 8'h2B; #100;
A = 8'hD; B = 8'h2C; #100;
A = 8'hD; B = 8'h2D; #100;
A = 8'hD; B = 8'h2E; #100;
A = 8'hD; B = 8'h2F; #100;
A = 8'hD; B = 8'h30; #100;
A = 8'hD; B = 8'h31; #100;
A = 8'hD; B = 8'h32; #100;
A = 8'hD; B = 8'h33; #100;
A = 8'hD; B = 8'h34; #100;
A = 8'hD; B = 8'h35; #100;
A = 8'hD; B = 8'h36; #100;
A = 8'hD; B = 8'h37; #100;
A = 8'hD; B = 8'h38; #100;
A = 8'hD; B = 8'h39; #100;
A = 8'hD; B = 8'h3A; #100;
A = 8'hD; B = 8'h3B; #100;
A = 8'hD; B = 8'h3C; #100;
A = 8'hD; B = 8'h3D; #100;
A = 8'hD; B = 8'h3E; #100;
A = 8'hD; B = 8'h3F; #100;
A = 8'hD; B = 8'h40; #100;
A = 8'hD; B = 8'h41; #100;
A = 8'hD; B = 8'h42; #100;
A = 8'hD; B = 8'h43; #100;
A = 8'hD; B = 8'h44; #100;
A = 8'hD; B = 8'h45; #100;
A = 8'hD; B = 8'h46; #100;
A = 8'hD; B = 8'h47; #100;
A = 8'hD; B = 8'h48; #100;
A = 8'hD; B = 8'h49; #100;
A = 8'hD; B = 8'h4A; #100;
A = 8'hD; B = 8'h4B; #100;
A = 8'hD; B = 8'h4C; #100;
A = 8'hD; B = 8'h4D; #100;
A = 8'hD; B = 8'h4E; #100;
A = 8'hD; B = 8'h4F; #100;
A = 8'hD; B = 8'h50; #100;
A = 8'hD; B = 8'h51; #100;
A = 8'hD; B = 8'h52; #100;
A = 8'hD; B = 8'h53; #100;
A = 8'hD; B = 8'h54; #100;
A = 8'hD; B = 8'h55; #100;
A = 8'hD; B = 8'h56; #100;
A = 8'hD; B = 8'h57; #100;
A = 8'hD; B = 8'h58; #100;
A = 8'hD; B = 8'h59; #100;
A = 8'hD; B = 8'h5A; #100;
A = 8'hD; B = 8'h5B; #100;
A = 8'hD; B = 8'h5C; #100;
A = 8'hD; B = 8'h5D; #100;
A = 8'hD; B = 8'h5E; #100;
A = 8'hD; B = 8'h5F; #100;
A = 8'hD; B = 8'h60; #100;
A = 8'hD; B = 8'h61; #100;
A = 8'hD; B = 8'h62; #100;
A = 8'hD; B = 8'h63; #100;
A = 8'hD; B = 8'h64; #100;
A = 8'hD; B = 8'h65; #100;
A = 8'hD; B = 8'h66; #100;
A = 8'hD; B = 8'h67; #100;
A = 8'hD; B = 8'h68; #100;
A = 8'hD; B = 8'h69; #100;
A = 8'hD; B = 8'h6A; #100;
A = 8'hD; B = 8'h6B; #100;
A = 8'hD; B = 8'h6C; #100;
A = 8'hD; B = 8'h6D; #100;
A = 8'hD; B = 8'h6E; #100;
A = 8'hD; B = 8'h6F; #100;
A = 8'hD; B = 8'h70; #100;
A = 8'hD; B = 8'h71; #100;
A = 8'hD; B = 8'h72; #100;
A = 8'hD; B = 8'h73; #100;
A = 8'hD; B = 8'h74; #100;
A = 8'hD; B = 8'h75; #100;
A = 8'hD; B = 8'h76; #100;
A = 8'hD; B = 8'h77; #100;
A = 8'hD; B = 8'h78; #100;
A = 8'hD; B = 8'h79; #100;
A = 8'hD; B = 8'h7A; #100;
A = 8'hD; B = 8'h7B; #100;
A = 8'hD; B = 8'h7C; #100;
A = 8'hD; B = 8'h7D; #100;
A = 8'hD; B = 8'h7E; #100;
A = 8'hD; B = 8'h7F; #100;
A = 8'hD; B = 8'h80; #100;
A = 8'hD; B = 8'h81; #100;
A = 8'hD; B = 8'h82; #100;
A = 8'hD; B = 8'h83; #100;
A = 8'hD; B = 8'h84; #100;
A = 8'hD; B = 8'h85; #100;
A = 8'hD; B = 8'h86; #100;
A = 8'hD; B = 8'h87; #100;
A = 8'hD; B = 8'h88; #100;
A = 8'hD; B = 8'h89; #100;
A = 8'hD; B = 8'h8A; #100;
A = 8'hD; B = 8'h8B; #100;
A = 8'hD; B = 8'h8C; #100;
A = 8'hD; B = 8'h8D; #100;
A = 8'hD; B = 8'h8E; #100;
A = 8'hD; B = 8'h8F; #100;
A = 8'hD; B = 8'h90; #100;
A = 8'hD; B = 8'h91; #100;
A = 8'hD; B = 8'h92; #100;
A = 8'hD; B = 8'h93; #100;
A = 8'hD; B = 8'h94; #100;
A = 8'hD; B = 8'h95; #100;
A = 8'hD; B = 8'h96; #100;
A = 8'hD; B = 8'h97; #100;
A = 8'hD; B = 8'h98; #100;
A = 8'hD; B = 8'h99; #100;
A = 8'hD; B = 8'h9A; #100;
A = 8'hD; B = 8'h9B; #100;
A = 8'hD; B = 8'h9C; #100;
A = 8'hD; B = 8'h9D; #100;
A = 8'hD; B = 8'h9E; #100;
A = 8'hD; B = 8'h9F; #100;
A = 8'hD; B = 8'hA0; #100;
A = 8'hD; B = 8'hA1; #100;
A = 8'hD; B = 8'hA2; #100;
A = 8'hD; B = 8'hA3; #100;
A = 8'hD; B = 8'hA4; #100;
A = 8'hD; B = 8'hA5; #100;
A = 8'hD; B = 8'hA6; #100;
A = 8'hD; B = 8'hA7; #100;
A = 8'hD; B = 8'hA8; #100;
A = 8'hD; B = 8'hA9; #100;
A = 8'hD; B = 8'hAA; #100;
A = 8'hD; B = 8'hAB; #100;
A = 8'hD; B = 8'hAC; #100;
A = 8'hD; B = 8'hAD; #100;
A = 8'hD; B = 8'hAE; #100;
A = 8'hD; B = 8'hAF; #100;
A = 8'hD; B = 8'hB0; #100;
A = 8'hD; B = 8'hB1; #100;
A = 8'hD; B = 8'hB2; #100;
A = 8'hD; B = 8'hB3; #100;
A = 8'hD; B = 8'hB4; #100;
A = 8'hD; B = 8'hB5; #100;
A = 8'hD; B = 8'hB6; #100;
A = 8'hD; B = 8'hB7; #100;
A = 8'hD; B = 8'hB8; #100;
A = 8'hD; B = 8'hB9; #100;
A = 8'hD; B = 8'hBA; #100;
A = 8'hD; B = 8'hBB; #100;
A = 8'hD; B = 8'hBC; #100;
A = 8'hD; B = 8'hBD; #100;
A = 8'hD; B = 8'hBE; #100;
A = 8'hD; B = 8'hBF; #100;
A = 8'hD; B = 8'hC0; #100;
A = 8'hD; B = 8'hC1; #100;
A = 8'hD; B = 8'hC2; #100;
A = 8'hD; B = 8'hC3; #100;
A = 8'hD; B = 8'hC4; #100;
A = 8'hD; B = 8'hC5; #100;
A = 8'hD; B = 8'hC6; #100;
A = 8'hD; B = 8'hC7; #100;
A = 8'hD; B = 8'hC8; #100;
A = 8'hD; B = 8'hC9; #100;
A = 8'hD; B = 8'hCA; #100;
A = 8'hD; B = 8'hCB; #100;
A = 8'hD; B = 8'hCC; #100;
A = 8'hD; B = 8'hCD; #100;
A = 8'hD; B = 8'hCE; #100;
A = 8'hD; B = 8'hCF; #100;
A = 8'hD; B = 8'hD0; #100;
A = 8'hD; B = 8'hD1; #100;
A = 8'hD; B = 8'hD2; #100;
A = 8'hD; B = 8'hD3; #100;
A = 8'hD; B = 8'hD4; #100;
A = 8'hD; B = 8'hD5; #100;
A = 8'hD; B = 8'hD6; #100;
A = 8'hD; B = 8'hD7; #100;
A = 8'hD; B = 8'hD8; #100;
A = 8'hD; B = 8'hD9; #100;
A = 8'hD; B = 8'hDA; #100;
A = 8'hD; B = 8'hDB; #100;
A = 8'hD; B = 8'hDC; #100;
A = 8'hD; B = 8'hDD; #100;
A = 8'hD; B = 8'hDE; #100;
A = 8'hD; B = 8'hDF; #100;
A = 8'hD; B = 8'hE0; #100;
A = 8'hD; B = 8'hE1; #100;
A = 8'hD; B = 8'hE2; #100;
A = 8'hD; B = 8'hE3; #100;
A = 8'hD; B = 8'hE4; #100;
A = 8'hD; B = 8'hE5; #100;
A = 8'hD; B = 8'hE6; #100;
A = 8'hD; B = 8'hE7; #100;
A = 8'hD; B = 8'hE8; #100;
A = 8'hD; B = 8'hE9; #100;
A = 8'hD; B = 8'hEA; #100;
A = 8'hD; B = 8'hEB; #100;
A = 8'hD; B = 8'hEC; #100;
A = 8'hD; B = 8'hED; #100;
A = 8'hD; B = 8'hEE; #100;
A = 8'hD; B = 8'hEF; #100;
A = 8'hD; B = 8'hF0; #100;
A = 8'hD; B = 8'hF1; #100;
A = 8'hD; B = 8'hF2; #100;
A = 8'hD; B = 8'hF3; #100;
A = 8'hD; B = 8'hF4; #100;
A = 8'hD; B = 8'hF5; #100;
A = 8'hD; B = 8'hF6; #100;
A = 8'hD; B = 8'hF7; #100;
A = 8'hD; B = 8'hF8; #100;
A = 8'hD; B = 8'hF9; #100;
A = 8'hD; B = 8'hFA; #100;
A = 8'hD; B = 8'hFB; #100;
A = 8'hD; B = 8'hFC; #100;
A = 8'hD; B = 8'hFD; #100;
A = 8'hD; B = 8'hFE; #100;
A = 8'hD; B = 8'hFF; #100;
A = 8'hE; B = 8'h0; #100;
A = 8'hE; B = 8'h1; #100;
A = 8'hE; B = 8'h2; #100;
A = 8'hE; B = 8'h3; #100;
A = 8'hE; B = 8'h4; #100;
A = 8'hE; B = 8'h5; #100;
A = 8'hE; B = 8'h6; #100;
A = 8'hE; B = 8'h7; #100;
A = 8'hE; B = 8'h8; #100;
A = 8'hE; B = 8'h9; #100;
A = 8'hE; B = 8'hA; #100;
A = 8'hE; B = 8'hB; #100;
A = 8'hE; B = 8'hC; #100;
A = 8'hE; B = 8'hD; #100;
A = 8'hE; B = 8'hE; #100;
A = 8'hE; B = 8'hF; #100;
A = 8'hE; B = 8'h10; #100;
A = 8'hE; B = 8'h11; #100;
A = 8'hE; B = 8'h12; #100;
A = 8'hE; B = 8'h13; #100;
A = 8'hE; B = 8'h14; #100;
A = 8'hE; B = 8'h15; #100;
A = 8'hE; B = 8'h16; #100;
A = 8'hE; B = 8'h17; #100;
A = 8'hE; B = 8'h18; #100;
A = 8'hE; B = 8'h19; #100;
A = 8'hE; B = 8'h1A; #100;
A = 8'hE; B = 8'h1B; #100;
A = 8'hE; B = 8'h1C; #100;
A = 8'hE; B = 8'h1D; #100;
A = 8'hE; B = 8'h1E; #100;
A = 8'hE; B = 8'h1F; #100;
A = 8'hE; B = 8'h20; #100;
A = 8'hE; B = 8'h21; #100;
A = 8'hE; B = 8'h22; #100;
A = 8'hE; B = 8'h23; #100;
A = 8'hE; B = 8'h24; #100;
A = 8'hE; B = 8'h25; #100;
A = 8'hE; B = 8'h26; #100;
A = 8'hE; B = 8'h27; #100;
A = 8'hE; B = 8'h28; #100;
A = 8'hE; B = 8'h29; #100;
A = 8'hE; B = 8'h2A; #100;
A = 8'hE; B = 8'h2B; #100;
A = 8'hE; B = 8'h2C; #100;
A = 8'hE; B = 8'h2D; #100;
A = 8'hE; B = 8'h2E; #100;
A = 8'hE; B = 8'h2F; #100;
A = 8'hE; B = 8'h30; #100;
A = 8'hE; B = 8'h31; #100;
A = 8'hE; B = 8'h32; #100;
A = 8'hE; B = 8'h33; #100;
A = 8'hE; B = 8'h34; #100;
A = 8'hE; B = 8'h35; #100;
A = 8'hE; B = 8'h36; #100;
A = 8'hE; B = 8'h37; #100;
A = 8'hE; B = 8'h38; #100;
A = 8'hE; B = 8'h39; #100;
A = 8'hE; B = 8'h3A; #100;
A = 8'hE; B = 8'h3B; #100;
A = 8'hE; B = 8'h3C; #100;
A = 8'hE; B = 8'h3D; #100;
A = 8'hE; B = 8'h3E; #100;
A = 8'hE; B = 8'h3F; #100;
A = 8'hE; B = 8'h40; #100;
A = 8'hE; B = 8'h41; #100;
A = 8'hE; B = 8'h42; #100;
A = 8'hE; B = 8'h43; #100;
A = 8'hE; B = 8'h44; #100;
A = 8'hE; B = 8'h45; #100;
A = 8'hE; B = 8'h46; #100;
A = 8'hE; B = 8'h47; #100;
A = 8'hE; B = 8'h48; #100;
A = 8'hE; B = 8'h49; #100;
A = 8'hE; B = 8'h4A; #100;
A = 8'hE; B = 8'h4B; #100;
A = 8'hE; B = 8'h4C; #100;
A = 8'hE; B = 8'h4D; #100;
A = 8'hE; B = 8'h4E; #100;
A = 8'hE; B = 8'h4F; #100;
A = 8'hE; B = 8'h50; #100;
A = 8'hE; B = 8'h51; #100;
A = 8'hE; B = 8'h52; #100;
A = 8'hE; B = 8'h53; #100;
A = 8'hE; B = 8'h54; #100;
A = 8'hE; B = 8'h55; #100;
A = 8'hE; B = 8'h56; #100;
A = 8'hE; B = 8'h57; #100;
A = 8'hE; B = 8'h58; #100;
A = 8'hE; B = 8'h59; #100;
A = 8'hE; B = 8'h5A; #100;
A = 8'hE; B = 8'h5B; #100;
A = 8'hE; B = 8'h5C; #100;
A = 8'hE; B = 8'h5D; #100;
A = 8'hE; B = 8'h5E; #100;
A = 8'hE; B = 8'h5F; #100;
A = 8'hE; B = 8'h60; #100;
A = 8'hE; B = 8'h61; #100;
A = 8'hE; B = 8'h62; #100;
A = 8'hE; B = 8'h63; #100;
A = 8'hE; B = 8'h64; #100;
A = 8'hE; B = 8'h65; #100;
A = 8'hE; B = 8'h66; #100;
A = 8'hE; B = 8'h67; #100;
A = 8'hE; B = 8'h68; #100;
A = 8'hE; B = 8'h69; #100;
A = 8'hE; B = 8'h6A; #100;
A = 8'hE; B = 8'h6B; #100;
A = 8'hE; B = 8'h6C; #100;
A = 8'hE; B = 8'h6D; #100;
A = 8'hE; B = 8'h6E; #100;
A = 8'hE; B = 8'h6F; #100;
A = 8'hE; B = 8'h70; #100;
A = 8'hE; B = 8'h71; #100;
A = 8'hE; B = 8'h72; #100;
A = 8'hE; B = 8'h73; #100;
A = 8'hE; B = 8'h74; #100;
A = 8'hE; B = 8'h75; #100;
A = 8'hE; B = 8'h76; #100;
A = 8'hE; B = 8'h77; #100;
A = 8'hE; B = 8'h78; #100;
A = 8'hE; B = 8'h79; #100;
A = 8'hE; B = 8'h7A; #100;
A = 8'hE; B = 8'h7B; #100;
A = 8'hE; B = 8'h7C; #100;
A = 8'hE; B = 8'h7D; #100;
A = 8'hE; B = 8'h7E; #100;
A = 8'hE; B = 8'h7F; #100;
A = 8'hE; B = 8'h80; #100;
A = 8'hE; B = 8'h81; #100;
A = 8'hE; B = 8'h82; #100;
A = 8'hE; B = 8'h83; #100;
A = 8'hE; B = 8'h84; #100;
A = 8'hE; B = 8'h85; #100;
A = 8'hE; B = 8'h86; #100;
A = 8'hE; B = 8'h87; #100;
A = 8'hE; B = 8'h88; #100;
A = 8'hE; B = 8'h89; #100;
A = 8'hE; B = 8'h8A; #100;
A = 8'hE; B = 8'h8B; #100;
A = 8'hE; B = 8'h8C; #100;
A = 8'hE; B = 8'h8D; #100;
A = 8'hE; B = 8'h8E; #100;
A = 8'hE; B = 8'h8F; #100;
A = 8'hE; B = 8'h90; #100;
A = 8'hE; B = 8'h91; #100;
A = 8'hE; B = 8'h92; #100;
A = 8'hE; B = 8'h93; #100;
A = 8'hE; B = 8'h94; #100;
A = 8'hE; B = 8'h95; #100;
A = 8'hE; B = 8'h96; #100;
A = 8'hE; B = 8'h97; #100;
A = 8'hE; B = 8'h98; #100;
A = 8'hE; B = 8'h99; #100;
A = 8'hE; B = 8'h9A; #100;
A = 8'hE; B = 8'h9B; #100;
A = 8'hE; B = 8'h9C; #100;
A = 8'hE; B = 8'h9D; #100;
A = 8'hE; B = 8'h9E; #100;
A = 8'hE; B = 8'h9F; #100;
A = 8'hE; B = 8'hA0; #100;
A = 8'hE; B = 8'hA1; #100;
A = 8'hE; B = 8'hA2; #100;
A = 8'hE; B = 8'hA3; #100;
A = 8'hE; B = 8'hA4; #100;
A = 8'hE; B = 8'hA5; #100;
A = 8'hE; B = 8'hA6; #100;
A = 8'hE; B = 8'hA7; #100;
A = 8'hE; B = 8'hA8; #100;
A = 8'hE; B = 8'hA9; #100;
A = 8'hE; B = 8'hAA; #100;
A = 8'hE; B = 8'hAB; #100;
A = 8'hE; B = 8'hAC; #100;
A = 8'hE; B = 8'hAD; #100;
A = 8'hE; B = 8'hAE; #100;
A = 8'hE; B = 8'hAF; #100;
A = 8'hE; B = 8'hB0; #100;
A = 8'hE; B = 8'hB1; #100;
A = 8'hE; B = 8'hB2; #100;
A = 8'hE; B = 8'hB3; #100;
A = 8'hE; B = 8'hB4; #100;
A = 8'hE; B = 8'hB5; #100;
A = 8'hE; B = 8'hB6; #100;
A = 8'hE; B = 8'hB7; #100;
A = 8'hE; B = 8'hB8; #100;
A = 8'hE; B = 8'hB9; #100;
A = 8'hE; B = 8'hBA; #100;
A = 8'hE; B = 8'hBB; #100;
A = 8'hE; B = 8'hBC; #100;
A = 8'hE; B = 8'hBD; #100;
A = 8'hE; B = 8'hBE; #100;
A = 8'hE; B = 8'hBF; #100;
A = 8'hE; B = 8'hC0; #100;
A = 8'hE; B = 8'hC1; #100;
A = 8'hE; B = 8'hC2; #100;
A = 8'hE; B = 8'hC3; #100;
A = 8'hE; B = 8'hC4; #100;
A = 8'hE; B = 8'hC5; #100;
A = 8'hE; B = 8'hC6; #100;
A = 8'hE; B = 8'hC7; #100;
A = 8'hE; B = 8'hC8; #100;
A = 8'hE; B = 8'hC9; #100;
A = 8'hE; B = 8'hCA; #100;
A = 8'hE; B = 8'hCB; #100;
A = 8'hE; B = 8'hCC; #100;
A = 8'hE; B = 8'hCD; #100;
A = 8'hE; B = 8'hCE; #100;
A = 8'hE; B = 8'hCF; #100;
A = 8'hE; B = 8'hD0; #100;
A = 8'hE; B = 8'hD1; #100;
A = 8'hE; B = 8'hD2; #100;
A = 8'hE; B = 8'hD3; #100;
A = 8'hE; B = 8'hD4; #100;
A = 8'hE; B = 8'hD5; #100;
A = 8'hE; B = 8'hD6; #100;
A = 8'hE; B = 8'hD7; #100;
A = 8'hE; B = 8'hD8; #100;
A = 8'hE; B = 8'hD9; #100;
A = 8'hE; B = 8'hDA; #100;
A = 8'hE; B = 8'hDB; #100;
A = 8'hE; B = 8'hDC; #100;
A = 8'hE; B = 8'hDD; #100;
A = 8'hE; B = 8'hDE; #100;
A = 8'hE; B = 8'hDF; #100;
A = 8'hE; B = 8'hE0; #100;
A = 8'hE; B = 8'hE1; #100;
A = 8'hE; B = 8'hE2; #100;
A = 8'hE; B = 8'hE3; #100;
A = 8'hE; B = 8'hE4; #100;
A = 8'hE; B = 8'hE5; #100;
A = 8'hE; B = 8'hE6; #100;
A = 8'hE; B = 8'hE7; #100;
A = 8'hE; B = 8'hE8; #100;
A = 8'hE; B = 8'hE9; #100;
A = 8'hE; B = 8'hEA; #100;
A = 8'hE; B = 8'hEB; #100;
A = 8'hE; B = 8'hEC; #100;
A = 8'hE; B = 8'hED; #100;
A = 8'hE; B = 8'hEE; #100;
A = 8'hE; B = 8'hEF; #100;
A = 8'hE; B = 8'hF0; #100;
A = 8'hE; B = 8'hF1; #100;
A = 8'hE; B = 8'hF2; #100;
A = 8'hE; B = 8'hF3; #100;
A = 8'hE; B = 8'hF4; #100;
A = 8'hE; B = 8'hF5; #100;
A = 8'hE; B = 8'hF6; #100;
A = 8'hE; B = 8'hF7; #100;
A = 8'hE; B = 8'hF8; #100;
A = 8'hE; B = 8'hF9; #100;
A = 8'hE; B = 8'hFA; #100;
A = 8'hE; B = 8'hFB; #100;
A = 8'hE; B = 8'hFC; #100;
A = 8'hE; B = 8'hFD; #100;
A = 8'hE; B = 8'hFE; #100;
A = 8'hE; B = 8'hFF; #100;
A = 8'hF; B = 8'h0; #100;
A = 8'hF; B = 8'h1; #100;
A = 8'hF; B = 8'h2; #100;
A = 8'hF; B = 8'h3; #100;
A = 8'hF; B = 8'h4; #100;
A = 8'hF; B = 8'h5; #100;
A = 8'hF; B = 8'h6; #100;
A = 8'hF; B = 8'h7; #100;
A = 8'hF; B = 8'h8; #100;
A = 8'hF; B = 8'h9; #100;
A = 8'hF; B = 8'hA; #100;
A = 8'hF; B = 8'hB; #100;
A = 8'hF; B = 8'hC; #100;
A = 8'hF; B = 8'hD; #100;
A = 8'hF; B = 8'hE; #100;
A = 8'hF; B = 8'hF; #100;
A = 8'hF; B = 8'h10; #100;
A = 8'hF; B = 8'h11; #100;
A = 8'hF; B = 8'h12; #100;
A = 8'hF; B = 8'h13; #100;
A = 8'hF; B = 8'h14; #100;
A = 8'hF; B = 8'h15; #100;
A = 8'hF; B = 8'h16; #100;
A = 8'hF; B = 8'h17; #100;
A = 8'hF; B = 8'h18; #100;
A = 8'hF; B = 8'h19; #100;
A = 8'hF; B = 8'h1A; #100;
A = 8'hF; B = 8'h1B; #100;
A = 8'hF; B = 8'h1C; #100;
A = 8'hF; B = 8'h1D; #100;
A = 8'hF; B = 8'h1E; #100;
A = 8'hF; B = 8'h1F; #100;
A = 8'hF; B = 8'h20; #100;
A = 8'hF; B = 8'h21; #100;
A = 8'hF; B = 8'h22; #100;
A = 8'hF; B = 8'h23; #100;
A = 8'hF; B = 8'h24; #100;
A = 8'hF; B = 8'h25; #100;
A = 8'hF; B = 8'h26; #100;
A = 8'hF; B = 8'h27; #100;
A = 8'hF; B = 8'h28; #100;
A = 8'hF; B = 8'h29; #100;
A = 8'hF; B = 8'h2A; #100;
A = 8'hF; B = 8'h2B; #100;
A = 8'hF; B = 8'h2C; #100;
A = 8'hF; B = 8'h2D; #100;
A = 8'hF; B = 8'h2E; #100;
A = 8'hF; B = 8'h2F; #100;
A = 8'hF; B = 8'h30; #100;
A = 8'hF; B = 8'h31; #100;
A = 8'hF; B = 8'h32; #100;
A = 8'hF; B = 8'h33; #100;
A = 8'hF; B = 8'h34; #100;
A = 8'hF; B = 8'h35; #100;
A = 8'hF; B = 8'h36; #100;
A = 8'hF; B = 8'h37; #100;
A = 8'hF; B = 8'h38; #100;
A = 8'hF; B = 8'h39; #100;
A = 8'hF; B = 8'h3A; #100;
A = 8'hF; B = 8'h3B; #100;
A = 8'hF; B = 8'h3C; #100;
A = 8'hF; B = 8'h3D; #100;
A = 8'hF; B = 8'h3E; #100;
A = 8'hF; B = 8'h3F; #100;
A = 8'hF; B = 8'h40; #100;
A = 8'hF; B = 8'h41; #100;
A = 8'hF; B = 8'h42; #100;
A = 8'hF; B = 8'h43; #100;
A = 8'hF; B = 8'h44; #100;
A = 8'hF; B = 8'h45; #100;
A = 8'hF; B = 8'h46; #100;
A = 8'hF; B = 8'h47; #100;
A = 8'hF; B = 8'h48; #100;
A = 8'hF; B = 8'h49; #100;
A = 8'hF; B = 8'h4A; #100;
A = 8'hF; B = 8'h4B; #100;
A = 8'hF; B = 8'h4C; #100;
A = 8'hF; B = 8'h4D; #100;
A = 8'hF; B = 8'h4E; #100;
A = 8'hF; B = 8'h4F; #100;
A = 8'hF; B = 8'h50; #100;
A = 8'hF; B = 8'h51; #100;
A = 8'hF; B = 8'h52; #100;
A = 8'hF; B = 8'h53; #100;
A = 8'hF; B = 8'h54; #100;
A = 8'hF; B = 8'h55; #100;
A = 8'hF; B = 8'h56; #100;
A = 8'hF; B = 8'h57; #100;
A = 8'hF; B = 8'h58; #100;
A = 8'hF; B = 8'h59; #100;
A = 8'hF; B = 8'h5A; #100;
A = 8'hF; B = 8'h5B; #100;
A = 8'hF; B = 8'h5C; #100;
A = 8'hF; B = 8'h5D; #100;
A = 8'hF; B = 8'h5E; #100;
A = 8'hF; B = 8'h5F; #100;
A = 8'hF; B = 8'h60; #100;
A = 8'hF; B = 8'h61; #100;
A = 8'hF; B = 8'h62; #100;
A = 8'hF; B = 8'h63; #100;
A = 8'hF; B = 8'h64; #100;
A = 8'hF; B = 8'h65; #100;
A = 8'hF; B = 8'h66; #100;
A = 8'hF; B = 8'h67; #100;
A = 8'hF; B = 8'h68; #100;
A = 8'hF; B = 8'h69; #100;
A = 8'hF; B = 8'h6A; #100;
A = 8'hF; B = 8'h6B; #100;
A = 8'hF; B = 8'h6C; #100;
A = 8'hF; B = 8'h6D; #100;
A = 8'hF; B = 8'h6E; #100;
A = 8'hF; B = 8'h6F; #100;
A = 8'hF; B = 8'h70; #100;
A = 8'hF; B = 8'h71; #100;
A = 8'hF; B = 8'h72; #100;
A = 8'hF; B = 8'h73; #100;
A = 8'hF; B = 8'h74; #100;
A = 8'hF; B = 8'h75; #100;
A = 8'hF; B = 8'h76; #100;
A = 8'hF; B = 8'h77; #100;
A = 8'hF; B = 8'h78; #100;
A = 8'hF; B = 8'h79; #100;
A = 8'hF; B = 8'h7A; #100;
A = 8'hF; B = 8'h7B; #100;
A = 8'hF; B = 8'h7C; #100;
A = 8'hF; B = 8'h7D; #100;
A = 8'hF; B = 8'h7E; #100;
A = 8'hF; B = 8'h7F; #100;
A = 8'hF; B = 8'h80; #100;
A = 8'hF; B = 8'h81; #100;
A = 8'hF; B = 8'h82; #100;
A = 8'hF; B = 8'h83; #100;
A = 8'hF; B = 8'h84; #100;
A = 8'hF; B = 8'h85; #100;
A = 8'hF; B = 8'h86; #100;
A = 8'hF; B = 8'h87; #100;
A = 8'hF; B = 8'h88; #100;
A = 8'hF; B = 8'h89; #100;
A = 8'hF; B = 8'h8A; #100;
A = 8'hF; B = 8'h8B; #100;
A = 8'hF; B = 8'h8C; #100;
A = 8'hF; B = 8'h8D; #100;
A = 8'hF; B = 8'h8E; #100;
A = 8'hF; B = 8'h8F; #100;
A = 8'hF; B = 8'h90; #100;
A = 8'hF; B = 8'h91; #100;
A = 8'hF; B = 8'h92; #100;
A = 8'hF; B = 8'h93; #100;
A = 8'hF; B = 8'h94; #100;
A = 8'hF; B = 8'h95; #100;
A = 8'hF; B = 8'h96; #100;
A = 8'hF; B = 8'h97; #100;
A = 8'hF; B = 8'h98; #100;
A = 8'hF; B = 8'h99; #100;
A = 8'hF; B = 8'h9A; #100;
A = 8'hF; B = 8'h9B; #100;
A = 8'hF; B = 8'h9C; #100;
A = 8'hF; B = 8'h9D; #100;
A = 8'hF; B = 8'h9E; #100;
A = 8'hF; B = 8'h9F; #100;
A = 8'hF; B = 8'hA0; #100;
A = 8'hF; B = 8'hA1; #100;
A = 8'hF; B = 8'hA2; #100;
A = 8'hF; B = 8'hA3; #100;
A = 8'hF; B = 8'hA4; #100;
A = 8'hF; B = 8'hA5; #100;
A = 8'hF; B = 8'hA6; #100;
A = 8'hF; B = 8'hA7; #100;
A = 8'hF; B = 8'hA8; #100;
A = 8'hF; B = 8'hA9; #100;
A = 8'hF; B = 8'hAA; #100;
A = 8'hF; B = 8'hAB; #100;
A = 8'hF; B = 8'hAC; #100;
A = 8'hF; B = 8'hAD; #100;
A = 8'hF; B = 8'hAE; #100;
A = 8'hF; B = 8'hAF; #100;
A = 8'hF; B = 8'hB0; #100;
A = 8'hF; B = 8'hB1; #100;
A = 8'hF; B = 8'hB2; #100;
A = 8'hF; B = 8'hB3; #100;
A = 8'hF; B = 8'hB4; #100;
A = 8'hF; B = 8'hB5; #100;
A = 8'hF; B = 8'hB6; #100;
A = 8'hF; B = 8'hB7; #100;
A = 8'hF; B = 8'hB8; #100;
A = 8'hF; B = 8'hB9; #100;
A = 8'hF; B = 8'hBA; #100;
A = 8'hF; B = 8'hBB; #100;
A = 8'hF; B = 8'hBC; #100;
A = 8'hF; B = 8'hBD; #100;
A = 8'hF; B = 8'hBE; #100;
A = 8'hF; B = 8'hBF; #100;
A = 8'hF; B = 8'hC0; #100;
A = 8'hF; B = 8'hC1; #100;
A = 8'hF; B = 8'hC2; #100;
A = 8'hF; B = 8'hC3; #100;
A = 8'hF; B = 8'hC4; #100;
A = 8'hF; B = 8'hC5; #100;
A = 8'hF; B = 8'hC6; #100;
A = 8'hF; B = 8'hC7; #100;
A = 8'hF; B = 8'hC8; #100;
A = 8'hF; B = 8'hC9; #100;
A = 8'hF; B = 8'hCA; #100;
A = 8'hF; B = 8'hCB; #100;
A = 8'hF; B = 8'hCC; #100;
A = 8'hF; B = 8'hCD; #100;
A = 8'hF; B = 8'hCE; #100;
A = 8'hF; B = 8'hCF; #100;
A = 8'hF; B = 8'hD0; #100;
A = 8'hF; B = 8'hD1; #100;
A = 8'hF; B = 8'hD2; #100;
A = 8'hF; B = 8'hD3; #100;
A = 8'hF; B = 8'hD4; #100;
A = 8'hF; B = 8'hD5; #100;
A = 8'hF; B = 8'hD6; #100;
A = 8'hF; B = 8'hD7; #100;
A = 8'hF; B = 8'hD8; #100;
A = 8'hF; B = 8'hD9; #100;
A = 8'hF; B = 8'hDA; #100;
A = 8'hF; B = 8'hDB; #100;
A = 8'hF; B = 8'hDC; #100;
A = 8'hF; B = 8'hDD; #100;
A = 8'hF; B = 8'hDE; #100;
A = 8'hF; B = 8'hDF; #100;
A = 8'hF; B = 8'hE0; #100;
A = 8'hF; B = 8'hE1; #100;
A = 8'hF; B = 8'hE2; #100;
A = 8'hF; B = 8'hE3; #100;
A = 8'hF; B = 8'hE4; #100;
A = 8'hF; B = 8'hE5; #100;
A = 8'hF; B = 8'hE6; #100;
A = 8'hF; B = 8'hE7; #100;
A = 8'hF; B = 8'hE8; #100;
A = 8'hF; B = 8'hE9; #100;
A = 8'hF; B = 8'hEA; #100;
A = 8'hF; B = 8'hEB; #100;
A = 8'hF; B = 8'hEC; #100;
A = 8'hF; B = 8'hED; #100;
A = 8'hF; B = 8'hEE; #100;
A = 8'hF; B = 8'hEF; #100;
A = 8'hF; B = 8'hF0; #100;
A = 8'hF; B = 8'hF1; #100;
A = 8'hF; B = 8'hF2; #100;
A = 8'hF; B = 8'hF3; #100;
A = 8'hF; B = 8'hF4; #100;
A = 8'hF; B = 8'hF5; #100;
A = 8'hF; B = 8'hF6; #100;
A = 8'hF; B = 8'hF7; #100;
A = 8'hF; B = 8'hF8; #100;
A = 8'hF; B = 8'hF9; #100;
A = 8'hF; B = 8'hFA; #100;
A = 8'hF; B = 8'hFB; #100;
A = 8'hF; B = 8'hFC; #100;
A = 8'hF; B = 8'hFD; #100;
A = 8'hF; B = 8'hFE; #100;
A = 8'hF; B = 8'hFF; #100;
A = 8'h10; B = 8'h0; #100;
A = 8'h10; B = 8'h1; #100;
A = 8'h10; B = 8'h2; #100;
A = 8'h10; B = 8'h3; #100;
A = 8'h10; B = 8'h4; #100;
A = 8'h10; B = 8'h5; #100;
A = 8'h10; B = 8'h6; #100;
A = 8'h10; B = 8'h7; #100;
A = 8'h10; B = 8'h8; #100;
A = 8'h10; B = 8'h9; #100;
A = 8'h10; B = 8'hA; #100;
A = 8'h10; B = 8'hB; #100;
A = 8'h10; B = 8'hC; #100;
A = 8'h10; B = 8'hD; #100;
A = 8'h10; B = 8'hE; #100;
A = 8'h10; B = 8'hF; #100;
A = 8'h10; B = 8'h10; #100;
A = 8'h10; B = 8'h11; #100;
A = 8'h10; B = 8'h12; #100;
A = 8'h10; B = 8'h13; #100;
A = 8'h10; B = 8'h14; #100;
A = 8'h10; B = 8'h15; #100;
A = 8'h10; B = 8'h16; #100;
A = 8'h10; B = 8'h17; #100;
A = 8'h10; B = 8'h18; #100;
A = 8'h10; B = 8'h19; #100;
A = 8'h10; B = 8'h1A; #100;
A = 8'h10; B = 8'h1B; #100;
A = 8'h10; B = 8'h1C; #100;
A = 8'h10; B = 8'h1D; #100;
A = 8'h10; B = 8'h1E; #100;
A = 8'h10; B = 8'h1F; #100;
A = 8'h10; B = 8'h20; #100;
A = 8'h10; B = 8'h21; #100;
A = 8'h10; B = 8'h22; #100;
A = 8'h10; B = 8'h23; #100;
A = 8'h10; B = 8'h24; #100;
A = 8'h10; B = 8'h25; #100;
A = 8'h10; B = 8'h26; #100;
A = 8'h10; B = 8'h27; #100;
A = 8'h10; B = 8'h28; #100;
A = 8'h10; B = 8'h29; #100;
A = 8'h10; B = 8'h2A; #100;
A = 8'h10; B = 8'h2B; #100;
A = 8'h10; B = 8'h2C; #100;
A = 8'h10; B = 8'h2D; #100;
A = 8'h10; B = 8'h2E; #100;
A = 8'h10; B = 8'h2F; #100;
A = 8'h10; B = 8'h30; #100;
A = 8'h10; B = 8'h31; #100;
A = 8'h10; B = 8'h32; #100;
A = 8'h10; B = 8'h33; #100;
A = 8'h10; B = 8'h34; #100;
A = 8'h10; B = 8'h35; #100;
A = 8'h10; B = 8'h36; #100;
A = 8'h10; B = 8'h37; #100;
A = 8'h10; B = 8'h38; #100;
A = 8'h10; B = 8'h39; #100;
A = 8'h10; B = 8'h3A; #100;
A = 8'h10; B = 8'h3B; #100;
A = 8'h10; B = 8'h3C; #100;
A = 8'h10; B = 8'h3D; #100;
A = 8'h10; B = 8'h3E; #100;
A = 8'h10; B = 8'h3F; #100;
A = 8'h10; B = 8'h40; #100;
A = 8'h10; B = 8'h41; #100;
A = 8'h10; B = 8'h42; #100;
A = 8'h10; B = 8'h43; #100;
A = 8'h10; B = 8'h44; #100;
A = 8'h10; B = 8'h45; #100;
A = 8'h10; B = 8'h46; #100;
A = 8'h10; B = 8'h47; #100;
A = 8'h10; B = 8'h48; #100;
A = 8'h10; B = 8'h49; #100;
A = 8'h10; B = 8'h4A; #100;
A = 8'h10; B = 8'h4B; #100;
A = 8'h10; B = 8'h4C; #100;
A = 8'h10; B = 8'h4D; #100;
A = 8'h10; B = 8'h4E; #100;
A = 8'h10; B = 8'h4F; #100;
A = 8'h10; B = 8'h50; #100;
A = 8'h10; B = 8'h51; #100;
A = 8'h10; B = 8'h52; #100;
A = 8'h10; B = 8'h53; #100;
A = 8'h10; B = 8'h54; #100;
A = 8'h10; B = 8'h55; #100;
A = 8'h10; B = 8'h56; #100;
A = 8'h10; B = 8'h57; #100;
A = 8'h10; B = 8'h58; #100;
A = 8'h10; B = 8'h59; #100;
A = 8'h10; B = 8'h5A; #100;
A = 8'h10; B = 8'h5B; #100;
A = 8'h10; B = 8'h5C; #100;
A = 8'h10; B = 8'h5D; #100;
A = 8'h10; B = 8'h5E; #100;
A = 8'h10; B = 8'h5F; #100;
A = 8'h10; B = 8'h60; #100;
A = 8'h10; B = 8'h61; #100;
A = 8'h10; B = 8'h62; #100;
A = 8'h10; B = 8'h63; #100;
A = 8'h10; B = 8'h64; #100;
A = 8'h10; B = 8'h65; #100;
A = 8'h10; B = 8'h66; #100;
A = 8'h10; B = 8'h67; #100;
A = 8'h10; B = 8'h68; #100;
A = 8'h10; B = 8'h69; #100;
A = 8'h10; B = 8'h6A; #100;
A = 8'h10; B = 8'h6B; #100;
A = 8'h10; B = 8'h6C; #100;
A = 8'h10; B = 8'h6D; #100;
A = 8'h10; B = 8'h6E; #100;
A = 8'h10; B = 8'h6F; #100;
A = 8'h10; B = 8'h70; #100;
A = 8'h10; B = 8'h71; #100;
A = 8'h10; B = 8'h72; #100;
A = 8'h10; B = 8'h73; #100;
A = 8'h10; B = 8'h74; #100;
A = 8'h10; B = 8'h75; #100;
A = 8'h10; B = 8'h76; #100;
A = 8'h10; B = 8'h77; #100;
A = 8'h10; B = 8'h78; #100;
A = 8'h10; B = 8'h79; #100;
A = 8'h10; B = 8'h7A; #100;
A = 8'h10; B = 8'h7B; #100;
A = 8'h10; B = 8'h7C; #100;
A = 8'h10; B = 8'h7D; #100;
A = 8'h10; B = 8'h7E; #100;
A = 8'h10; B = 8'h7F; #100;
A = 8'h10; B = 8'h80; #100;
A = 8'h10; B = 8'h81; #100;
A = 8'h10; B = 8'h82; #100;
A = 8'h10; B = 8'h83; #100;
A = 8'h10; B = 8'h84; #100;
A = 8'h10; B = 8'h85; #100;
A = 8'h10; B = 8'h86; #100;
A = 8'h10; B = 8'h87; #100;
A = 8'h10; B = 8'h88; #100;
A = 8'h10; B = 8'h89; #100;
A = 8'h10; B = 8'h8A; #100;
A = 8'h10; B = 8'h8B; #100;
A = 8'h10; B = 8'h8C; #100;
A = 8'h10; B = 8'h8D; #100;
A = 8'h10; B = 8'h8E; #100;
A = 8'h10; B = 8'h8F; #100;
A = 8'h10; B = 8'h90; #100;
A = 8'h10; B = 8'h91; #100;
A = 8'h10; B = 8'h92; #100;
A = 8'h10; B = 8'h93; #100;
A = 8'h10; B = 8'h94; #100;
A = 8'h10; B = 8'h95; #100;
A = 8'h10; B = 8'h96; #100;
A = 8'h10; B = 8'h97; #100;
A = 8'h10; B = 8'h98; #100;
A = 8'h10; B = 8'h99; #100;
A = 8'h10; B = 8'h9A; #100;
A = 8'h10; B = 8'h9B; #100;
A = 8'h10; B = 8'h9C; #100;
A = 8'h10; B = 8'h9D; #100;
A = 8'h10; B = 8'h9E; #100;
A = 8'h10; B = 8'h9F; #100;
A = 8'h10; B = 8'hA0; #100;
A = 8'h10; B = 8'hA1; #100;
A = 8'h10; B = 8'hA2; #100;
A = 8'h10; B = 8'hA3; #100;
A = 8'h10; B = 8'hA4; #100;
A = 8'h10; B = 8'hA5; #100;
A = 8'h10; B = 8'hA6; #100;
A = 8'h10; B = 8'hA7; #100;
A = 8'h10; B = 8'hA8; #100;
A = 8'h10; B = 8'hA9; #100;
A = 8'h10; B = 8'hAA; #100;
A = 8'h10; B = 8'hAB; #100;
A = 8'h10; B = 8'hAC; #100;
A = 8'h10; B = 8'hAD; #100;
A = 8'h10; B = 8'hAE; #100;
A = 8'h10; B = 8'hAF; #100;
A = 8'h10; B = 8'hB0; #100;
A = 8'h10; B = 8'hB1; #100;
A = 8'h10; B = 8'hB2; #100;
A = 8'h10; B = 8'hB3; #100;
A = 8'h10; B = 8'hB4; #100;
A = 8'h10; B = 8'hB5; #100;
A = 8'h10; B = 8'hB6; #100;
A = 8'h10; B = 8'hB7; #100;
A = 8'h10; B = 8'hB8; #100;
A = 8'h10; B = 8'hB9; #100;
A = 8'h10; B = 8'hBA; #100;
A = 8'h10; B = 8'hBB; #100;
A = 8'h10; B = 8'hBC; #100;
A = 8'h10; B = 8'hBD; #100;
A = 8'h10; B = 8'hBE; #100;
A = 8'h10; B = 8'hBF; #100;
A = 8'h10; B = 8'hC0; #100;
A = 8'h10; B = 8'hC1; #100;
A = 8'h10; B = 8'hC2; #100;
A = 8'h10; B = 8'hC3; #100;
A = 8'h10; B = 8'hC4; #100;
A = 8'h10; B = 8'hC5; #100;
A = 8'h10; B = 8'hC6; #100;
A = 8'h10; B = 8'hC7; #100;
A = 8'h10; B = 8'hC8; #100;
A = 8'h10; B = 8'hC9; #100;
A = 8'h10; B = 8'hCA; #100;
A = 8'h10; B = 8'hCB; #100;
A = 8'h10; B = 8'hCC; #100;
A = 8'h10; B = 8'hCD; #100;
A = 8'h10; B = 8'hCE; #100;
A = 8'h10; B = 8'hCF; #100;
A = 8'h10; B = 8'hD0; #100;
A = 8'h10; B = 8'hD1; #100;
A = 8'h10; B = 8'hD2; #100;
A = 8'h10; B = 8'hD3; #100;
A = 8'h10; B = 8'hD4; #100;
A = 8'h10; B = 8'hD5; #100;
A = 8'h10; B = 8'hD6; #100;
A = 8'h10; B = 8'hD7; #100;
A = 8'h10; B = 8'hD8; #100;
A = 8'h10; B = 8'hD9; #100;
A = 8'h10; B = 8'hDA; #100;
A = 8'h10; B = 8'hDB; #100;
A = 8'h10; B = 8'hDC; #100;
A = 8'h10; B = 8'hDD; #100;
A = 8'h10; B = 8'hDE; #100;
A = 8'h10; B = 8'hDF; #100;
A = 8'h10; B = 8'hE0; #100;
A = 8'h10; B = 8'hE1; #100;
A = 8'h10; B = 8'hE2; #100;
A = 8'h10; B = 8'hE3; #100;
A = 8'h10; B = 8'hE4; #100;
A = 8'h10; B = 8'hE5; #100;
A = 8'h10; B = 8'hE6; #100;
A = 8'h10; B = 8'hE7; #100;
A = 8'h10; B = 8'hE8; #100;
A = 8'h10; B = 8'hE9; #100;
A = 8'h10; B = 8'hEA; #100;
A = 8'h10; B = 8'hEB; #100;
A = 8'h10; B = 8'hEC; #100;
A = 8'h10; B = 8'hED; #100;
A = 8'h10; B = 8'hEE; #100;
A = 8'h10; B = 8'hEF; #100;
A = 8'h10; B = 8'hF0; #100;
A = 8'h10; B = 8'hF1; #100;
A = 8'h10; B = 8'hF2; #100;
A = 8'h10; B = 8'hF3; #100;
A = 8'h10; B = 8'hF4; #100;
A = 8'h10; B = 8'hF5; #100;
A = 8'h10; B = 8'hF6; #100;
A = 8'h10; B = 8'hF7; #100;
A = 8'h10; B = 8'hF8; #100;
A = 8'h10; B = 8'hF9; #100;
A = 8'h10; B = 8'hFA; #100;
A = 8'h10; B = 8'hFB; #100;
A = 8'h10; B = 8'hFC; #100;
A = 8'h10; B = 8'hFD; #100;
A = 8'h10; B = 8'hFE; #100;
A = 8'h10; B = 8'hFF; #100;
A = 8'h11; B = 8'h0; #100;
A = 8'h11; B = 8'h1; #100;
A = 8'h11; B = 8'h2; #100;
A = 8'h11; B = 8'h3; #100;
A = 8'h11; B = 8'h4; #100;
A = 8'h11; B = 8'h5; #100;
A = 8'h11; B = 8'h6; #100;
A = 8'h11; B = 8'h7; #100;
A = 8'h11; B = 8'h8; #100;
A = 8'h11; B = 8'h9; #100;
A = 8'h11; B = 8'hA; #100;
A = 8'h11; B = 8'hB; #100;
A = 8'h11; B = 8'hC; #100;
A = 8'h11; B = 8'hD; #100;
A = 8'h11; B = 8'hE; #100;
A = 8'h11; B = 8'hF; #100;
A = 8'h11; B = 8'h10; #100;
A = 8'h11; B = 8'h11; #100;
A = 8'h11; B = 8'h12; #100;
A = 8'h11; B = 8'h13; #100;
A = 8'h11; B = 8'h14; #100;
A = 8'h11; B = 8'h15; #100;
A = 8'h11; B = 8'h16; #100;
A = 8'h11; B = 8'h17; #100;
A = 8'h11; B = 8'h18; #100;
A = 8'h11; B = 8'h19; #100;
A = 8'h11; B = 8'h1A; #100;
A = 8'h11; B = 8'h1B; #100;
A = 8'h11; B = 8'h1C; #100;
A = 8'h11; B = 8'h1D; #100;
A = 8'h11; B = 8'h1E; #100;
A = 8'h11; B = 8'h1F; #100;
A = 8'h11; B = 8'h20; #100;
A = 8'h11; B = 8'h21; #100;
A = 8'h11; B = 8'h22; #100;
A = 8'h11; B = 8'h23; #100;
A = 8'h11; B = 8'h24; #100;
A = 8'h11; B = 8'h25; #100;
A = 8'h11; B = 8'h26; #100;
A = 8'h11; B = 8'h27; #100;
A = 8'h11; B = 8'h28; #100;
A = 8'h11; B = 8'h29; #100;
A = 8'h11; B = 8'h2A; #100;
A = 8'h11; B = 8'h2B; #100;
A = 8'h11; B = 8'h2C; #100;
A = 8'h11; B = 8'h2D; #100;
A = 8'h11; B = 8'h2E; #100;
A = 8'h11; B = 8'h2F; #100;
A = 8'h11; B = 8'h30; #100;
A = 8'h11; B = 8'h31; #100;
A = 8'h11; B = 8'h32; #100;
A = 8'h11; B = 8'h33; #100;
A = 8'h11; B = 8'h34; #100;
A = 8'h11; B = 8'h35; #100;
A = 8'h11; B = 8'h36; #100;
A = 8'h11; B = 8'h37; #100;
A = 8'h11; B = 8'h38; #100;
A = 8'h11; B = 8'h39; #100;
A = 8'h11; B = 8'h3A; #100;
A = 8'h11; B = 8'h3B; #100;
A = 8'h11; B = 8'h3C; #100;
A = 8'h11; B = 8'h3D; #100;
A = 8'h11; B = 8'h3E; #100;
A = 8'h11; B = 8'h3F; #100;
A = 8'h11; B = 8'h40; #100;
A = 8'h11; B = 8'h41; #100;
A = 8'h11; B = 8'h42; #100;
A = 8'h11; B = 8'h43; #100;
A = 8'h11; B = 8'h44; #100;
A = 8'h11; B = 8'h45; #100;
A = 8'h11; B = 8'h46; #100;
A = 8'h11; B = 8'h47; #100;
A = 8'h11; B = 8'h48; #100;
A = 8'h11; B = 8'h49; #100;
A = 8'h11; B = 8'h4A; #100;
A = 8'h11; B = 8'h4B; #100;
A = 8'h11; B = 8'h4C; #100;
A = 8'h11; B = 8'h4D; #100;
A = 8'h11; B = 8'h4E; #100;
A = 8'h11; B = 8'h4F; #100;
A = 8'h11; B = 8'h50; #100;
A = 8'h11; B = 8'h51; #100;
A = 8'h11; B = 8'h52; #100;
A = 8'h11; B = 8'h53; #100;
A = 8'h11; B = 8'h54; #100;
A = 8'h11; B = 8'h55; #100;
A = 8'h11; B = 8'h56; #100;
A = 8'h11; B = 8'h57; #100;
A = 8'h11; B = 8'h58; #100;
A = 8'h11; B = 8'h59; #100;
A = 8'h11; B = 8'h5A; #100;
A = 8'h11; B = 8'h5B; #100;
A = 8'h11; B = 8'h5C; #100;
A = 8'h11; B = 8'h5D; #100;
A = 8'h11; B = 8'h5E; #100;
A = 8'h11; B = 8'h5F; #100;
A = 8'h11; B = 8'h60; #100;
A = 8'h11; B = 8'h61; #100;
A = 8'h11; B = 8'h62; #100;
A = 8'h11; B = 8'h63; #100;
A = 8'h11; B = 8'h64; #100;
A = 8'h11; B = 8'h65; #100;
A = 8'h11; B = 8'h66; #100;
A = 8'h11; B = 8'h67; #100;
A = 8'h11; B = 8'h68; #100;
A = 8'h11; B = 8'h69; #100;
A = 8'h11; B = 8'h6A; #100;
A = 8'h11; B = 8'h6B; #100;
A = 8'h11; B = 8'h6C; #100;
A = 8'h11; B = 8'h6D; #100;
A = 8'h11; B = 8'h6E; #100;
A = 8'h11; B = 8'h6F; #100;
A = 8'h11; B = 8'h70; #100;
A = 8'h11; B = 8'h71; #100;
A = 8'h11; B = 8'h72; #100;
A = 8'h11; B = 8'h73; #100;
A = 8'h11; B = 8'h74; #100;
A = 8'h11; B = 8'h75; #100;
A = 8'h11; B = 8'h76; #100;
A = 8'h11; B = 8'h77; #100;
A = 8'h11; B = 8'h78; #100;
A = 8'h11; B = 8'h79; #100;
A = 8'h11; B = 8'h7A; #100;
A = 8'h11; B = 8'h7B; #100;
A = 8'h11; B = 8'h7C; #100;
A = 8'h11; B = 8'h7D; #100;
A = 8'h11; B = 8'h7E; #100;
A = 8'h11; B = 8'h7F; #100;
A = 8'h11; B = 8'h80; #100;
A = 8'h11; B = 8'h81; #100;
A = 8'h11; B = 8'h82; #100;
A = 8'h11; B = 8'h83; #100;
A = 8'h11; B = 8'h84; #100;
A = 8'h11; B = 8'h85; #100;
A = 8'h11; B = 8'h86; #100;
A = 8'h11; B = 8'h87; #100;
A = 8'h11; B = 8'h88; #100;
A = 8'h11; B = 8'h89; #100;
A = 8'h11; B = 8'h8A; #100;
A = 8'h11; B = 8'h8B; #100;
A = 8'h11; B = 8'h8C; #100;
A = 8'h11; B = 8'h8D; #100;
A = 8'h11; B = 8'h8E; #100;
A = 8'h11; B = 8'h8F; #100;
A = 8'h11; B = 8'h90; #100;
A = 8'h11; B = 8'h91; #100;
A = 8'h11; B = 8'h92; #100;
A = 8'h11; B = 8'h93; #100;
A = 8'h11; B = 8'h94; #100;
A = 8'h11; B = 8'h95; #100;
A = 8'h11; B = 8'h96; #100;
A = 8'h11; B = 8'h97; #100;
A = 8'h11; B = 8'h98; #100;
A = 8'h11; B = 8'h99; #100;
A = 8'h11; B = 8'h9A; #100;
A = 8'h11; B = 8'h9B; #100;
A = 8'h11; B = 8'h9C; #100;
A = 8'h11; B = 8'h9D; #100;
A = 8'h11; B = 8'h9E; #100;
A = 8'h11; B = 8'h9F; #100;
A = 8'h11; B = 8'hA0; #100;
A = 8'h11; B = 8'hA1; #100;
A = 8'h11; B = 8'hA2; #100;
A = 8'h11; B = 8'hA3; #100;
A = 8'h11; B = 8'hA4; #100;
A = 8'h11; B = 8'hA5; #100;
A = 8'h11; B = 8'hA6; #100;
A = 8'h11; B = 8'hA7; #100;
A = 8'h11; B = 8'hA8; #100;
A = 8'h11; B = 8'hA9; #100;
A = 8'h11; B = 8'hAA; #100;
A = 8'h11; B = 8'hAB; #100;
A = 8'h11; B = 8'hAC; #100;
A = 8'h11; B = 8'hAD; #100;
A = 8'h11; B = 8'hAE; #100;
A = 8'h11; B = 8'hAF; #100;
A = 8'h11; B = 8'hB0; #100;
A = 8'h11; B = 8'hB1; #100;
A = 8'h11; B = 8'hB2; #100;
A = 8'h11; B = 8'hB3; #100;
A = 8'h11; B = 8'hB4; #100;
A = 8'h11; B = 8'hB5; #100;
A = 8'h11; B = 8'hB6; #100;
A = 8'h11; B = 8'hB7; #100;
A = 8'h11; B = 8'hB8; #100;
A = 8'h11; B = 8'hB9; #100;
A = 8'h11; B = 8'hBA; #100;
A = 8'h11; B = 8'hBB; #100;
A = 8'h11; B = 8'hBC; #100;
A = 8'h11; B = 8'hBD; #100;
A = 8'h11; B = 8'hBE; #100;
A = 8'h11; B = 8'hBF; #100;
A = 8'h11; B = 8'hC0; #100;
A = 8'h11; B = 8'hC1; #100;
A = 8'h11; B = 8'hC2; #100;
A = 8'h11; B = 8'hC3; #100;
A = 8'h11; B = 8'hC4; #100;
A = 8'h11; B = 8'hC5; #100;
A = 8'h11; B = 8'hC6; #100;
A = 8'h11; B = 8'hC7; #100;
A = 8'h11; B = 8'hC8; #100;
A = 8'h11; B = 8'hC9; #100;
A = 8'h11; B = 8'hCA; #100;
A = 8'h11; B = 8'hCB; #100;
A = 8'h11; B = 8'hCC; #100;
A = 8'h11; B = 8'hCD; #100;
A = 8'h11; B = 8'hCE; #100;
A = 8'h11; B = 8'hCF; #100;
A = 8'h11; B = 8'hD0; #100;
A = 8'h11; B = 8'hD1; #100;
A = 8'h11; B = 8'hD2; #100;
A = 8'h11; B = 8'hD3; #100;
A = 8'h11; B = 8'hD4; #100;
A = 8'h11; B = 8'hD5; #100;
A = 8'h11; B = 8'hD6; #100;
A = 8'h11; B = 8'hD7; #100;
A = 8'h11; B = 8'hD8; #100;
A = 8'h11; B = 8'hD9; #100;
A = 8'h11; B = 8'hDA; #100;
A = 8'h11; B = 8'hDB; #100;
A = 8'h11; B = 8'hDC; #100;
A = 8'h11; B = 8'hDD; #100;
A = 8'h11; B = 8'hDE; #100;
A = 8'h11; B = 8'hDF; #100;
A = 8'h11; B = 8'hE0; #100;
A = 8'h11; B = 8'hE1; #100;
A = 8'h11; B = 8'hE2; #100;
A = 8'h11; B = 8'hE3; #100;
A = 8'h11; B = 8'hE4; #100;
A = 8'h11; B = 8'hE5; #100;
A = 8'h11; B = 8'hE6; #100;
A = 8'h11; B = 8'hE7; #100;
A = 8'h11; B = 8'hE8; #100;
A = 8'h11; B = 8'hE9; #100;
A = 8'h11; B = 8'hEA; #100;
A = 8'h11; B = 8'hEB; #100;
A = 8'h11; B = 8'hEC; #100;
A = 8'h11; B = 8'hED; #100;
A = 8'h11; B = 8'hEE; #100;
A = 8'h11; B = 8'hEF; #100;
A = 8'h11; B = 8'hF0; #100;
A = 8'h11; B = 8'hF1; #100;
A = 8'h11; B = 8'hF2; #100;
A = 8'h11; B = 8'hF3; #100;
A = 8'h11; B = 8'hF4; #100;
A = 8'h11; B = 8'hF5; #100;
A = 8'h11; B = 8'hF6; #100;
A = 8'h11; B = 8'hF7; #100;
A = 8'h11; B = 8'hF8; #100;
A = 8'h11; B = 8'hF9; #100;
A = 8'h11; B = 8'hFA; #100;
A = 8'h11; B = 8'hFB; #100;
A = 8'h11; B = 8'hFC; #100;
A = 8'h11; B = 8'hFD; #100;
A = 8'h11; B = 8'hFE; #100;
A = 8'h11; B = 8'hFF; #100;
A = 8'h12; B = 8'h0; #100;
A = 8'h12; B = 8'h1; #100;
A = 8'h12; B = 8'h2; #100;
A = 8'h12; B = 8'h3; #100;
A = 8'h12; B = 8'h4; #100;
A = 8'h12; B = 8'h5; #100;
A = 8'h12; B = 8'h6; #100;
A = 8'h12; B = 8'h7; #100;
A = 8'h12; B = 8'h8; #100;
A = 8'h12; B = 8'h9; #100;
A = 8'h12; B = 8'hA; #100;
A = 8'h12; B = 8'hB; #100;
A = 8'h12; B = 8'hC; #100;
A = 8'h12; B = 8'hD; #100;
A = 8'h12; B = 8'hE; #100;
A = 8'h12; B = 8'hF; #100;
A = 8'h12; B = 8'h10; #100;
A = 8'h12; B = 8'h11; #100;
A = 8'h12; B = 8'h12; #100;
A = 8'h12; B = 8'h13; #100;
A = 8'h12; B = 8'h14; #100;
A = 8'h12; B = 8'h15; #100;
A = 8'h12; B = 8'h16; #100;
A = 8'h12; B = 8'h17; #100;
A = 8'h12; B = 8'h18; #100;
A = 8'h12; B = 8'h19; #100;
A = 8'h12; B = 8'h1A; #100;
A = 8'h12; B = 8'h1B; #100;
A = 8'h12; B = 8'h1C; #100;
A = 8'h12; B = 8'h1D; #100;
A = 8'h12; B = 8'h1E; #100;
A = 8'h12; B = 8'h1F; #100;
A = 8'h12; B = 8'h20; #100;
A = 8'h12; B = 8'h21; #100;
A = 8'h12; B = 8'h22; #100;
A = 8'h12; B = 8'h23; #100;
A = 8'h12; B = 8'h24; #100;
A = 8'h12; B = 8'h25; #100;
A = 8'h12; B = 8'h26; #100;
A = 8'h12; B = 8'h27; #100;
A = 8'h12; B = 8'h28; #100;
A = 8'h12; B = 8'h29; #100;
A = 8'h12; B = 8'h2A; #100;
A = 8'h12; B = 8'h2B; #100;
A = 8'h12; B = 8'h2C; #100;
A = 8'h12; B = 8'h2D; #100;
A = 8'h12; B = 8'h2E; #100;
A = 8'h12; B = 8'h2F; #100;
A = 8'h12; B = 8'h30; #100;
A = 8'h12; B = 8'h31; #100;
A = 8'h12; B = 8'h32; #100;
A = 8'h12; B = 8'h33; #100;
A = 8'h12; B = 8'h34; #100;
A = 8'h12; B = 8'h35; #100;
A = 8'h12; B = 8'h36; #100;
A = 8'h12; B = 8'h37; #100;
A = 8'h12; B = 8'h38; #100;
A = 8'h12; B = 8'h39; #100;
A = 8'h12; B = 8'h3A; #100;
A = 8'h12; B = 8'h3B; #100;
A = 8'h12; B = 8'h3C; #100;
A = 8'h12; B = 8'h3D; #100;
A = 8'h12; B = 8'h3E; #100;
A = 8'h12; B = 8'h3F; #100;
A = 8'h12; B = 8'h40; #100;
A = 8'h12; B = 8'h41; #100;
A = 8'h12; B = 8'h42; #100;
A = 8'h12; B = 8'h43; #100;
A = 8'h12; B = 8'h44; #100;
A = 8'h12; B = 8'h45; #100;
A = 8'h12; B = 8'h46; #100;
A = 8'h12; B = 8'h47; #100;
A = 8'h12; B = 8'h48; #100;
A = 8'h12; B = 8'h49; #100;
A = 8'h12; B = 8'h4A; #100;
A = 8'h12; B = 8'h4B; #100;
A = 8'h12; B = 8'h4C; #100;
A = 8'h12; B = 8'h4D; #100;
A = 8'h12; B = 8'h4E; #100;
A = 8'h12; B = 8'h4F; #100;
A = 8'h12; B = 8'h50; #100;
A = 8'h12; B = 8'h51; #100;
A = 8'h12; B = 8'h52; #100;
A = 8'h12; B = 8'h53; #100;
A = 8'h12; B = 8'h54; #100;
A = 8'h12; B = 8'h55; #100;
A = 8'h12; B = 8'h56; #100;
A = 8'h12; B = 8'h57; #100;
A = 8'h12; B = 8'h58; #100;
A = 8'h12; B = 8'h59; #100;
A = 8'h12; B = 8'h5A; #100;
A = 8'h12; B = 8'h5B; #100;
A = 8'h12; B = 8'h5C; #100;
A = 8'h12; B = 8'h5D; #100;
A = 8'h12; B = 8'h5E; #100;
A = 8'h12; B = 8'h5F; #100;
A = 8'h12; B = 8'h60; #100;
A = 8'h12; B = 8'h61; #100;
A = 8'h12; B = 8'h62; #100;
A = 8'h12; B = 8'h63; #100;
A = 8'h12; B = 8'h64; #100;
A = 8'h12; B = 8'h65; #100;
A = 8'h12; B = 8'h66; #100;
A = 8'h12; B = 8'h67; #100;
A = 8'h12; B = 8'h68; #100;
A = 8'h12; B = 8'h69; #100;
A = 8'h12; B = 8'h6A; #100;
A = 8'h12; B = 8'h6B; #100;
A = 8'h12; B = 8'h6C; #100;
A = 8'h12; B = 8'h6D; #100;
A = 8'h12; B = 8'h6E; #100;
A = 8'h12; B = 8'h6F; #100;
A = 8'h12; B = 8'h70; #100;
A = 8'h12; B = 8'h71; #100;
A = 8'h12; B = 8'h72; #100;
A = 8'h12; B = 8'h73; #100;
A = 8'h12; B = 8'h74; #100;
A = 8'h12; B = 8'h75; #100;
A = 8'h12; B = 8'h76; #100;
A = 8'h12; B = 8'h77; #100;
A = 8'h12; B = 8'h78; #100;
A = 8'h12; B = 8'h79; #100;
A = 8'h12; B = 8'h7A; #100;
A = 8'h12; B = 8'h7B; #100;
A = 8'h12; B = 8'h7C; #100;
A = 8'h12; B = 8'h7D; #100;
A = 8'h12; B = 8'h7E; #100;
A = 8'h12; B = 8'h7F; #100;
A = 8'h12; B = 8'h80; #100;
A = 8'h12; B = 8'h81; #100;
A = 8'h12; B = 8'h82; #100;
A = 8'h12; B = 8'h83; #100;
A = 8'h12; B = 8'h84; #100;
A = 8'h12; B = 8'h85; #100;
A = 8'h12; B = 8'h86; #100;
A = 8'h12; B = 8'h87; #100;
A = 8'h12; B = 8'h88; #100;
A = 8'h12; B = 8'h89; #100;
A = 8'h12; B = 8'h8A; #100;
A = 8'h12; B = 8'h8B; #100;
A = 8'h12; B = 8'h8C; #100;
A = 8'h12; B = 8'h8D; #100;
A = 8'h12; B = 8'h8E; #100;
A = 8'h12; B = 8'h8F; #100;
A = 8'h12; B = 8'h90; #100;
A = 8'h12; B = 8'h91; #100;
A = 8'h12; B = 8'h92; #100;
A = 8'h12; B = 8'h93; #100;
A = 8'h12; B = 8'h94; #100;
A = 8'h12; B = 8'h95; #100;
A = 8'h12; B = 8'h96; #100;
A = 8'h12; B = 8'h97; #100;
A = 8'h12; B = 8'h98; #100;
A = 8'h12; B = 8'h99; #100;
A = 8'h12; B = 8'h9A; #100;
A = 8'h12; B = 8'h9B; #100;
A = 8'h12; B = 8'h9C; #100;
A = 8'h12; B = 8'h9D; #100;
A = 8'h12; B = 8'h9E; #100;
A = 8'h12; B = 8'h9F; #100;
A = 8'h12; B = 8'hA0; #100;
A = 8'h12; B = 8'hA1; #100;
A = 8'h12; B = 8'hA2; #100;
A = 8'h12; B = 8'hA3; #100;
A = 8'h12; B = 8'hA4; #100;
A = 8'h12; B = 8'hA5; #100;
A = 8'h12; B = 8'hA6; #100;
A = 8'h12; B = 8'hA7; #100;
A = 8'h12; B = 8'hA8; #100;
A = 8'h12; B = 8'hA9; #100;
A = 8'h12; B = 8'hAA; #100;
A = 8'h12; B = 8'hAB; #100;
A = 8'h12; B = 8'hAC; #100;
A = 8'h12; B = 8'hAD; #100;
A = 8'h12; B = 8'hAE; #100;
A = 8'h12; B = 8'hAF; #100;
A = 8'h12; B = 8'hB0; #100;
A = 8'h12; B = 8'hB1; #100;
A = 8'h12; B = 8'hB2; #100;
A = 8'h12; B = 8'hB3; #100;
A = 8'h12; B = 8'hB4; #100;
A = 8'h12; B = 8'hB5; #100;
A = 8'h12; B = 8'hB6; #100;
A = 8'h12; B = 8'hB7; #100;
A = 8'h12; B = 8'hB8; #100;
A = 8'h12; B = 8'hB9; #100;
A = 8'h12; B = 8'hBA; #100;
A = 8'h12; B = 8'hBB; #100;
A = 8'h12; B = 8'hBC; #100;
A = 8'h12; B = 8'hBD; #100;
A = 8'h12; B = 8'hBE; #100;
A = 8'h12; B = 8'hBF; #100;
A = 8'h12; B = 8'hC0; #100;
A = 8'h12; B = 8'hC1; #100;
A = 8'h12; B = 8'hC2; #100;
A = 8'h12; B = 8'hC3; #100;
A = 8'h12; B = 8'hC4; #100;
A = 8'h12; B = 8'hC5; #100;
A = 8'h12; B = 8'hC6; #100;
A = 8'h12; B = 8'hC7; #100;
A = 8'h12; B = 8'hC8; #100;
A = 8'h12; B = 8'hC9; #100;
A = 8'h12; B = 8'hCA; #100;
A = 8'h12; B = 8'hCB; #100;
A = 8'h12; B = 8'hCC; #100;
A = 8'h12; B = 8'hCD; #100;
A = 8'h12; B = 8'hCE; #100;
A = 8'h12; B = 8'hCF; #100;
A = 8'h12; B = 8'hD0; #100;
A = 8'h12; B = 8'hD1; #100;
A = 8'h12; B = 8'hD2; #100;
A = 8'h12; B = 8'hD3; #100;
A = 8'h12; B = 8'hD4; #100;
A = 8'h12; B = 8'hD5; #100;
A = 8'h12; B = 8'hD6; #100;
A = 8'h12; B = 8'hD7; #100;
A = 8'h12; B = 8'hD8; #100;
A = 8'h12; B = 8'hD9; #100;
A = 8'h12; B = 8'hDA; #100;
A = 8'h12; B = 8'hDB; #100;
A = 8'h12; B = 8'hDC; #100;
A = 8'h12; B = 8'hDD; #100;
A = 8'h12; B = 8'hDE; #100;
A = 8'h12; B = 8'hDF; #100;
A = 8'h12; B = 8'hE0; #100;
A = 8'h12; B = 8'hE1; #100;
A = 8'h12; B = 8'hE2; #100;
A = 8'h12; B = 8'hE3; #100;
A = 8'h12; B = 8'hE4; #100;
A = 8'h12; B = 8'hE5; #100;
A = 8'h12; B = 8'hE6; #100;
A = 8'h12; B = 8'hE7; #100;
A = 8'h12; B = 8'hE8; #100;
A = 8'h12; B = 8'hE9; #100;
A = 8'h12; B = 8'hEA; #100;
A = 8'h12; B = 8'hEB; #100;
A = 8'h12; B = 8'hEC; #100;
A = 8'h12; B = 8'hED; #100;
A = 8'h12; B = 8'hEE; #100;
A = 8'h12; B = 8'hEF; #100;
A = 8'h12; B = 8'hF0; #100;
A = 8'h12; B = 8'hF1; #100;
A = 8'h12; B = 8'hF2; #100;
A = 8'h12; B = 8'hF3; #100;
A = 8'h12; B = 8'hF4; #100;
A = 8'h12; B = 8'hF5; #100;
A = 8'h12; B = 8'hF6; #100;
A = 8'h12; B = 8'hF7; #100;
A = 8'h12; B = 8'hF8; #100;
A = 8'h12; B = 8'hF9; #100;
A = 8'h12; B = 8'hFA; #100;
A = 8'h12; B = 8'hFB; #100;
A = 8'h12; B = 8'hFC; #100;
A = 8'h12; B = 8'hFD; #100;
A = 8'h12; B = 8'hFE; #100;
A = 8'h12; B = 8'hFF; #100;
A = 8'h13; B = 8'h0; #100;
A = 8'h13; B = 8'h1; #100;
A = 8'h13; B = 8'h2; #100;
A = 8'h13; B = 8'h3; #100;
A = 8'h13; B = 8'h4; #100;
A = 8'h13; B = 8'h5; #100;
A = 8'h13; B = 8'h6; #100;
A = 8'h13; B = 8'h7; #100;
A = 8'h13; B = 8'h8; #100;
A = 8'h13; B = 8'h9; #100;
A = 8'h13; B = 8'hA; #100;
A = 8'h13; B = 8'hB; #100;
A = 8'h13; B = 8'hC; #100;
A = 8'h13; B = 8'hD; #100;
A = 8'h13; B = 8'hE; #100;
A = 8'h13; B = 8'hF; #100;
A = 8'h13; B = 8'h10; #100;
A = 8'h13; B = 8'h11; #100;
A = 8'h13; B = 8'h12; #100;
A = 8'h13; B = 8'h13; #100;
A = 8'h13; B = 8'h14; #100;
A = 8'h13; B = 8'h15; #100;
A = 8'h13; B = 8'h16; #100;
A = 8'h13; B = 8'h17; #100;
A = 8'h13; B = 8'h18; #100;
A = 8'h13; B = 8'h19; #100;
A = 8'h13; B = 8'h1A; #100;
A = 8'h13; B = 8'h1B; #100;
A = 8'h13; B = 8'h1C; #100;
A = 8'h13; B = 8'h1D; #100;
A = 8'h13; B = 8'h1E; #100;
A = 8'h13; B = 8'h1F; #100;
A = 8'h13; B = 8'h20; #100;
A = 8'h13; B = 8'h21; #100;
A = 8'h13; B = 8'h22; #100;
A = 8'h13; B = 8'h23; #100;
A = 8'h13; B = 8'h24; #100;
A = 8'h13; B = 8'h25; #100;
A = 8'h13; B = 8'h26; #100;
A = 8'h13; B = 8'h27; #100;
A = 8'h13; B = 8'h28; #100;
A = 8'h13; B = 8'h29; #100;
A = 8'h13; B = 8'h2A; #100;
A = 8'h13; B = 8'h2B; #100;
A = 8'h13; B = 8'h2C; #100;
A = 8'h13; B = 8'h2D; #100;
A = 8'h13; B = 8'h2E; #100;
A = 8'h13; B = 8'h2F; #100;
A = 8'h13; B = 8'h30; #100;
A = 8'h13; B = 8'h31; #100;
A = 8'h13; B = 8'h32; #100;
A = 8'h13; B = 8'h33; #100;
A = 8'h13; B = 8'h34; #100;
A = 8'h13; B = 8'h35; #100;
A = 8'h13; B = 8'h36; #100;
A = 8'h13; B = 8'h37; #100;
A = 8'h13; B = 8'h38; #100;
A = 8'h13; B = 8'h39; #100;
A = 8'h13; B = 8'h3A; #100;
A = 8'h13; B = 8'h3B; #100;
A = 8'h13; B = 8'h3C; #100;
A = 8'h13; B = 8'h3D; #100;
A = 8'h13; B = 8'h3E; #100;
A = 8'h13; B = 8'h3F; #100;
A = 8'h13; B = 8'h40; #100;
A = 8'h13; B = 8'h41; #100;
A = 8'h13; B = 8'h42; #100;
A = 8'h13; B = 8'h43; #100;
A = 8'h13; B = 8'h44; #100;
A = 8'h13; B = 8'h45; #100;
A = 8'h13; B = 8'h46; #100;
A = 8'h13; B = 8'h47; #100;
A = 8'h13; B = 8'h48; #100;
A = 8'h13; B = 8'h49; #100;
A = 8'h13; B = 8'h4A; #100;
A = 8'h13; B = 8'h4B; #100;
A = 8'h13; B = 8'h4C; #100;
A = 8'h13; B = 8'h4D; #100;
A = 8'h13; B = 8'h4E; #100;
A = 8'h13; B = 8'h4F; #100;
A = 8'h13; B = 8'h50; #100;
A = 8'h13; B = 8'h51; #100;
A = 8'h13; B = 8'h52; #100;
A = 8'h13; B = 8'h53; #100;
A = 8'h13; B = 8'h54; #100;
A = 8'h13; B = 8'h55; #100;
A = 8'h13; B = 8'h56; #100;
A = 8'h13; B = 8'h57; #100;
A = 8'h13; B = 8'h58; #100;
A = 8'h13; B = 8'h59; #100;
A = 8'h13; B = 8'h5A; #100;
A = 8'h13; B = 8'h5B; #100;
A = 8'h13; B = 8'h5C; #100;
A = 8'h13; B = 8'h5D; #100;
A = 8'h13; B = 8'h5E; #100;
A = 8'h13; B = 8'h5F; #100;
A = 8'h13; B = 8'h60; #100;
A = 8'h13; B = 8'h61; #100;
A = 8'h13; B = 8'h62; #100;
A = 8'h13; B = 8'h63; #100;
A = 8'h13; B = 8'h64; #100;
A = 8'h13; B = 8'h65; #100;
A = 8'h13; B = 8'h66; #100;
A = 8'h13; B = 8'h67; #100;
A = 8'h13; B = 8'h68; #100;
A = 8'h13; B = 8'h69; #100;
A = 8'h13; B = 8'h6A; #100;
A = 8'h13; B = 8'h6B; #100;
A = 8'h13; B = 8'h6C; #100;
A = 8'h13; B = 8'h6D; #100;
A = 8'h13; B = 8'h6E; #100;
A = 8'h13; B = 8'h6F; #100;
A = 8'h13; B = 8'h70; #100;
A = 8'h13; B = 8'h71; #100;
A = 8'h13; B = 8'h72; #100;
A = 8'h13; B = 8'h73; #100;
A = 8'h13; B = 8'h74; #100;
A = 8'h13; B = 8'h75; #100;
A = 8'h13; B = 8'h76; #100;
A = 8'h13; B = 8'h77; #100;
A = 8'h13; B = 8'h78; #100;
A = 8'h13; B = 8'h79; #100;
A = 8'h13; B = 8'h7A; #100;
A = 8'h13; B = 8'h7B; #100;
A = 8'h13; B = 8'h7C; #100;
A = 8'h13; B = 8'h7D; #100;
A = 8'h13; B = 8'h7E; #100;
A = 8'h13; B = 8'h7F; #100;
A = 8'h13; B = 8'h80; #100;
A = 8'h13; B = 8'h81; #100;
A = 8'h13; B = 8'h82; #100;
A = 8'h13; B = 8'h83; #100;
A = 8'h13; B = 8'h84; #100;
A = 8'h13; B = 8'h85; #100;
A = 8'h13; B = 8'h86; #100;
A = 8'h13; B = 8'h87; #100;
A = 8'h13; B = 8'h88; #100;
A = 8'h13; B = 8'h89; #100;
A = 8'h13; B = 8'h8A; #100;
A = 8'h13; B = 8'h8B; #100;
A = 8'h13; B = 8'h8C; #100;
A = 8'h13; B = 8'h8D; #100;
A = 8'h13; B = 8'h8E; #100;
A = 8'h13; B = 8'h8F; #100;
A = 8'h13; B = 8'h90; #100;
A = 8'h13; B = 8'h91; #100;
A = 8'h13; B = 8'h92; #100;
A = 8'h13; B = 8'h93; #100;
A = 8'h13; B = 8'h94; #100;
A = 8'h13; B = 8'h95; #100;
A = 8'h13; B = 8'h96; #100;
A = 8'h13; B = 8'h97; #100;
A = 8'h13; B = 8'h98; #100;
A = 8'h13; B = 8'h99; #100;
A = 8'h13; B = 8'h9A; #100;
A = 8'h13; B = 8'h9B; #100;
A = 8'h13; B = 8'h9C; #100;
A = 8'h13; B = 8'h9D; #100;
A = 8'h13; B = 8'h9E; #100;
A = 8'h13; B = 8'h9F; #100;
A = 8'h13; B = 8'hA0; #100;
A = 8'h13; B = 8'hA1; #100;
A = 8'h13; B = 8'hA2; #100;
A = 8'h13; B = 8'hA3; #100;
A = 8'h13; B = 8'hA4; #100;
A = 8'h13; B = 8'hA5; #100;
A = 8'h13; B = 8'hA6; #100;
A = 8'h13; B = 8'hA7; #100;
A = 8'h13; B = 8'hA8; #100;
A = 8'h13; B = 8'hA9; #100;
A = 8'h13; B = 8'hAA; #100;
A = 8'h13; B = 8'hAB; #100;
A = 8'h13; B = 8'hAC; #100;
A = 8'h13; B = 8'hAD; #100;
A = 8'h13; B = 8'hAE; #100;
A = 8'h13; B = 8'hAF; #100;
A = 8'h13; B = 8'hB0; #100;
A = 8'h13; B = 8'hB1; #100;
A = 8'h13; B = 8'hB2; #100;
A = 8'h13; B = 8'hB3; #100;
A = 8'h13; B = 8'hB4; #100;
A = 8'h13; B = 8'hB5; #100;
A = 8'h13; B = 8'hB6; #100;
A = 8'h13; B = 8'hB7; #100;
A = 8'h13; B = 8'hB8; #100;
A = 8'h13; B = 8'hB9; #100;
A = 8'h13; B = 8'hBA; #100;
A = 8'h13; B = 8'hBB; #100;
A = 8'h13; B = 8'hBC; #100;
A = 8'h13; B = 8'hBD; #100;
A = 8'h13; B = 8'hBE; #100;
A = 8'h13; B = 8'hBF; #100;
A = 8'h13; B = 8'hC0; #100;
A = 8'h13; B = 8'hC1; #100;
A = 8'h13; B = 8'hC2; #100;
A = 8'h13; B = 8'hC3; #100;
A = 8'h13; B = 8'hC4; #100;
A = 8'h13; B = 8'hC5; #100;
A = 8'h13; B = 8'hC6; #100;
A = 8'h13; B = 8'hC7; #100;
A = 8'h13; B = 8'hC8; #100;
A = 8'h13; B = 8'hC9; #100;
A = 8'h13; B = 8'hCA; #100;
A = 8'h13; B = 8'hCB; #100;
A = 8'h13; B = 8'hCC; #100;
A = 8'h13; B = 8'hCD; #100;
A = 8'h13; B = 8'hCE; #100;
A = 8'h13; B = 8'hCF; #100;
A = 8'h13; B = 8'hD0; #100;
A = 8'h13; B = 8'hD1; #100;
A = 8'h13; B = 8'hD2; #100;
A = 8'h13; B = 8'hD3; #100;
A = 8'h13; B = 8'hD4; #100;
A = 8'h13; B = 8'hD5; #100;
A = 8'h13; B = 8'hD6; #100;
A = 8'h13; B = 8'hD7; #100;
A = 8'h13; B = 8'hD8; #100;
A = 8'h13; B = 8'hD9; #100;
A = 8'h13; B = 8'hDA; #100;
A = 8'h13; B = 8'hDB; #100;
A = 8'h13; B = 8'hDC; #100;
A = 8'h13; B = 8'hDD; #100;
A = 8'h13; B = 8'hDE; #100;
A = 8'h13; B = 8'hDF; #100;
A = 8'h13; B = 8'hE0; #100;
A = 8'h13; B = 8'hE1; #100;
A = 8'h13; B = 8'hE2; #100;
A = 8'h13; B = 8'hE3; #100;
A = 8'h13; B = 8'hE4; #100;
A = 8'h13; B = 8'hE5; #100;
A = 8'h13; B = 8'hE6; #100;
A = 8'h13; B = 8'hE7; #100;
A = 8'h13; B = 8'hE8; #100;
A = 8'h13; B = 8'hE9; #100;
A = 8'h13; B = 8'hEA; #100;
A = 8'h13; B = 8'hEB; #100;
A = 8'h13; B = 8'hEC; #100;
A = 8'h13; B = 8'hED; #100;
A = 8'h13; B = 8'hEE; #100;
A = 8'h13; B = 8'hEF; #100;
A = 8'h13; B = 8'hF0; #100;
A = 8'h13; B = 8'hF1; #100;
A = 8'h13; B = 8'hF2; #100;
A = 8'h13; B = 8'hF3; #100;
A = 8'h13; B = 8'hF4; #100;
A = 8'h13; B = 8'hF5; #100;
A = 8'h13; B = 8'hF6; #100;
A = 8'h13; B = 8'hF7; #100;
A = 8'h13; B = 8'hF8; #100;
A = 8'h13; B = 8'hF9; #100;
A = 8'h13; B = 8'hFA; #100;
A = 8'h13; B = 8'hFB; #100;
A = 8'h13; B = 8'hFC; #100;
A = 8'h13; B = 8'hFD; #100;
A = 8'h13; B = 8'hFE; #100;
A = 8'h13; B = 8'hFF; #100;
A = 8'h14; B = 8'h0; #100;
A = 8'h14; B = 8'h1; #100;
A = 8'h14; B = 8'h2; #100;
A = 8'h14; B = 8'h3; #100;
A = 8'h14; B = 8'h4; #100;
A = 8'h14; B = 8'h5; #100;
A = 8'h14; B = 8'h6; #100;
A = 8'h14; B = 8'h7; #100;
A = 8'h14; B = 8'h8; #100;
A = 8'h14; B = 8'h9; #100;
A = 8'h14; B = 8'hA; #100;
A = 8'h14; B = 8'hB; #100;
A = 8'h14; B = 8'hC; #100;
A = 8'h14; B = 8'hD; #100;
A = 8'h14; B = 8'hE; #100;
A = 8'h14; B = 8'hF; #100;
A = 8'h14; B = 8'h10; #100;
A = 8'h14; B = 8'h11; #100;
A = 8'h14; B = 8'h12; #100;
A = 8'h14; B = 8'h13; #100;
A = 8'h14; B = 8'h14; #100;
A = 8'h14; B = 8'h15; #100;
A = 8'h14; B = 8'h16; #100;
A = 8'h14; B = 8'h17; #100;
A = 8'h14; B = 8'h18; #100;
A = 8'h14; B = 8'h19; #100;
A = 8'h14; B = 8'h1A; #100;
A = 8'h14; B = 8'h1B; #100;
A = 8'h14; B = 8'h1C; #100;
A = 8'h14; B = 8'h1D; #100;
A = 8'h14; B = 8'h1E; #100;
A = 8'h14; B = 8'h1F; #100;
A = 8'h14; B = 8'h20; #100;
A = 8'h14; B = 8'h21; #100;
A = 8'h14; B = 8'h22; #100;
A = 8'h14; B = 8'h23; #100;
A = 8'h14; B = 8'h24; #100;
A = 8'h14; B = 8'h25; #100;
A = 8'h14; B = 8'h26; #100;
A = 8'h14; B = 8'h27; #100;
A = 8'h14; B = 8'h28; #100;
A = 8'h14; B = 8'h29; #100;
A = 8'h14; B = 8'h2A; #100;
A = 8'h14; B = 8'h2B; #100;
A = 8'h14; B = 8'h2C; #100;
A = 8'h14; B = 8'h2D; #100;
A = 8'h14; B = 8'h2E; #100;
A = 8'h14; B = 8'h2F; #100;
A = 8'h14; B = 8'h30; #100;
A = 8'h14; B = 8'h31; #100;
A = 8'h14; B = 8'h32; #100;
A = 8'h14; B = 8'h33; #100;
A = 8'h14; B = 8'h34; #100;
A = 8'h14; B = 8'h35; #100;
A = 8'h14; B = 8'h36; #100;
A = 8'h14; B = 8'h37; #100;
A = 8'h14; B = 8'h38; #100;
A = 8'h14; B = 8'h39; #100;
A = 8'h14; B = 8'h3A; #100;
A = 8'h14; B = 8'h3B; #100;
A = 8'h14; B = 8'h3C; #100;
A = 8'h14; B = 8'h3D; #100;
A = 8'h14; B = 8'h3E; #100;
A = 8'h14; B = 8'h3F; #100;
A = 8'h14; B = 8'h40; #100;
A = 8'h14; B = 8'h41; #100;
A = 8'h14; B = 8'h42; #100;
A = 8'h14; B = 8'h43; #100;
A = 8'h14; B = 8'h44; #100;
A = 8'h14; B = 8'h45; #100;
A = 8'h14; B = 8'h46; #100;
A = 8'h14; B = 8'h47; #100;
A = 8'h14; B = 8'h48; #100;
A = 8'h14; B = 8'h49; #100;
A = 8'h14; B = 8'h4A; #100;
A = 8'h14; B = 8'h4B; #100;
A = 8'h14; B = 8'h4C; #100;
A = 8'h14; B = 8'h4D; #100;
A = 8'h14; B = 8'h4E; #100;
A = 8'h14; B = 8'h4F; #100;
A = 8'h14; B = 8'h50; #100;
A = 8'h14; B = 8'h51; #100;
A = 8'h14; B = 8'h52; #100;
A = 8'h14; B = 8'h53; #100;
A = 8'h14; B = 8'h54; #100;
A = 8'h14; B = 8'h55; #100;
A = 8'h14; B = 8'h56; #100;
A = 8'h14; B = 8'h57; #100;
A = 8'h14; B = 8'h58; #100;
A = 8'h14; B = 8'h59; #100;
A = 8'h14; B = 8'h5A; #100;
A = 8'h14; B = 8'h5B; #100;
A = 8'h14; B = 8'h5C; #100;
A = 8'h14; B = 8'h5D; #100;
A = 8'h14; B = 8'h5E; #100;
A = 8'h14; B = 8'h5F; #100;
A = 8'h14; B = 8'h60; #100;
A = 8'h14; B = 8'h61; #100;
A = 8'h14; B = 8'h62; #100;
A = 8'h14; B = 8'h63; #100;
A = 8'h14; B = 8'h64; #100;
A = 8'h14; B = 8'h65; #100;
A = 8'h14; B = 8'h66; #100;
A = 8'h14; B = 8'h67; #100;
A = 8'h14; B = 8'h68; #100;
A = 8'h14; B = 8'h69; #100;
A = 8'h14; B = 8'h6A; #100;
A = 8'h14; B = 8'h6B; #100;
A = 8'h14; B = 8'h6C; #100;
A = 8'h14; B = 8'h6D; #100;
A = 8'h14; B = 8'h6E; #100;
A = 8'h14; B = 8'h6F; #100;
A = 8'h14; B = 8'h70; #100;
A = 8'h14; B = 8'h71; #100;
A = 8'h14; B = 8'h72; #100;
A = 8'h14; B = 8'h73; #100;
A = 8'h14; B = 8'h74; #100;
A = 8'h14; B = 8'h75; #100;
A = 8'h14; B = 8'h76; #100;
A = 8'h14; B = 8'h77; #100;
A = 8'h14; B = 8'h78; #100;
A = 8'h14; B = 8'h79; #100;
A = 8'h14; B = 8'h7A; #100;
A = 8'h14; B = 8'h7B; #100;
A = 8'h14; B = 8'h7C; #100;
A = 8'h14; B = 8'h7D; #100;
A = 8'h14; B = 8'h7E; #100;
A = 8'h14; B = 8'h7F; #100;
A = 8'h14; B = 8'h80; #100;
A = 8'h14; B = 8'h81; #100;
A = 8'h14; B = 8'h82; #100;
A = 8'h14; B = 8'h83; #100;
A = 8'h14; B = 8'h84; #100;
A = 8'h14; B = 8'h85; #100;
A = 8'h14; B = 8'h86; #100;
A = 8'h14; B = 8'h87; #100;
A = 8'h14; B = 8'h88; #100;
A = 8'h14; B = 8'h89; #100;
A = 8'h14; B = 8'h8A; #100;
A = 8'h14; B = 8'h8B; #100;
A = 8'h14; B = 8'h8C; #100;
A = 8'h14; B = 8'h8D; #100;
A = 8'h14; B = 8'h8E; #100;
A = 8'h14; B = 8'h8F; #100;
A = 8'h14; B = 8'h90; #100;
A = 8'h14; B = 8'h91; #100;
A = 8'h14; B = 8'h92; #100;
A = 8'h14; B = 8'h93; #100;
A = 8'h14; B = 8'h94; #100;
A = 8'h14; B = 8'h95; #100;
A = 8'h14; B = 8'h96; #100;
A = 8'h14; B = 8'h97; #100;
A = 8'h14; B = 8'h98; #100;
A = 8'h14; B = 8'h99; #100;
A = 8'h14; B = 8'h9A; #100;
A = 8'h14; B = 8'h9B; #100;
A = 8'h14; B = 8'h9C; #100;
A = 8'h14; B = 8'h9D; #100;
A = 8'h14; B = 8'h9E; #100;
A = 8'h14; B = 8'h9F; #100;
A = 8'h14; B = 8'hA0; #100;
A = 8'h14; B = 8'hA1; #100;
A = 8'h14; B = 8'hA2; #100;
A = 8'h14; B = 8'hA3; #100;
A = 8'h14; B = 8'hA4; #100;
A = 8'h14; B = 8'hA5; #100;
A = 8'h14; B = 8'hA6; #100;
A = 8'h14; B = 8'hA7; #100;
A = 8'h14; B = 8'hA8; #100;
A = 8'h14; B = 8'hA9; #100;
A = 8'h14; B = 8'hAA; #100;
A = 8'h14; B = 8'hAB; #100;
A = 8'h14; B = 8'hAC; #100;
A = 8'h14; B = 8'hAD; #100;
A = 8'h14; B = 8'hAE; #100;
A = 8'h14; B = 8'hAF; #100;
A = 8'h14; B = 8'hB0; #100;
A = 8'h14; B = 8'hB1; #100;
A = 8'h14; B = 8'hB2; #100;
A = 8'h14; B = 8'hB3; #100;
A = 8'h14; B = 8'hB4; #100;
A = 8'h14; B = 8'hB5; #100;
A = 8'h14; B = 8'hB6; #100;
A = 8'h14; B = 8'hB7; #100;
A = 8'h14; B = 8'hB8; #100;
A = 8'h14; B = 8'hB9; #100;
A = 8'h14; B = 8'hBA; #100;
A = 8'h14; B = 8'hBB; #100;
A = 8'h14; B = 8'hBC; #100;
A = 8'h14; B = 8'hBD; #100;
A = 8'h14; B = 8'hBE; #100;
A = 8'h14; B = 8'hBF; #100;
A = 8'h14; B = 8'hC0; #100;
A = 8'h14; B = 8'hC1; #100;
A = 8'h14; B = 8'hC2; #100;
A = 8'h14; B = 8'hC3; #100;
A = 8'h14; B = 8'hC4; #100;
A = 8'h14; B = 8'hC5; #100;
A = 8'h14; B = 8'hC6; #100;
A = 8'h14; B = 8'hC7; #100;
A = 8'h14; B = 8'hC8; #100;
A = 8'h14; B = 8'hC9; #100;
A = 8'h14; B = 8'hCA; #100;
A = 8'h14; B = 8'hCB; #100;
A = 8'h14; B = 8'hCC; #100;
A = 8'h14; B = 8'hCD; #100;
A = 8'h14; B = 8'hCE; #100;
A = 8'h14; B = 8'hCF; #100;
A = 8'h14; B = 8'hD0; #100;
A = 8'h14; B = 8'hD1; #100;
A = 8'h14; B = 8'hD2; #100;
A = 8'h14; B = 8'hD3; #100;
A = 8'h14; B = 8'hD4; #100;
A = 8'h14; B = 8'hD5; #100;
A = 8'h14; B = 8'hD6; #100;
A = 8'h14; B = 8'hD7; #100;
A = 8'h14; B = 8'hD8; #100;
A = 8'h14; B = 8'hD9; #100;
A = 8'h14; B = 8'hDA; #100;
A = 8'h14; B = 8'hDB; #100;
A = 8'h14; B = 8'hDC; #100;
A = 8'h14; B = 8'hDD; #100;
A = 8'h14; B = 8'hDE; #100;
A = 8'h14; B = 8'hDF; #100;
A = 8'h14; B = 8'hE0; #100;
A = 8'h14; B = 8'hE1; #100;
A = 8'h14; B = 8'hE2; #100;
A = 8'h14; B = 8'hE3; #100;
A = 8'h14; B = 8'hE4; #100;
A = 8'h14; B = 8'hE5; #100;
A = 8'h14; B = 8'hE6; #100;
A = 8'h14; B = 8'hE7; #100;
A = 8'h14; B = 8'hE8; #100;
A = 8'h14; B = 8'hE9; #100;
A = 8'h14; B = 8'hEA; #100;
A = 8'h14; B = 8'hEB; #100;
A = 8'h14; B = 8'hEC; #100;
A = 8'h14; B = 8'hED; #100;
A = 8'h14; B = 8'hEE; #100;
A = 8'h14; B = 8'hEF; #100;
A = 8'h14; B = 8'hF0; #100;
A = 8'h14; B = 8'hF1; #100;
A = 8'h14; B = 8'hF2; #100;
A = 8'h14; B = 8'hF3; #100;
A = 8'h14; B = 8'hF4; #100;
A = 8'h14; B = 8'hF5; #100;
A = 8'h14; B = 8'hF6; #100;
A = 8'h14; B = 8'hF7; #100;
A = 8'h14; B = 8'hF8; #100;
A = 8'h14; B = 8'hF9; #100;
A = 8'h14; B = 8'hFA; #100;
A = 8'h14; B = 8'hFB; #100;
A = 8'h14; B = 8'hFC; #100;
A = 8'h14; B = 8'hFD; #100;
A = 8'h14; B = 8'hFE; #100;
A = 8'h14; B = 8'hFF; #100;
A = 8'h15; B = 8'h0; #100;
A = 8'h15; B = 8'h1; #100;
A = 8'h15; B = 8'h2; #100;
A = 8'h15; B = 8'h3; #100;
A = 8'h15; B = 8'h4; #100;
A = 8'h15; B = 8'h5; #100;
A = 8'h15; B = 8'h6; #100;
A = 8'h15; B = 8'h7; #100;
A = 8'h15; B = 8'h8; #100;
A = 8'h15; B = 8'h9; #100;
A = 8'h15; B = 8'hA; #100;
A = 8'h15; B = 8'hB; #100;
A = 8'h15; B = 8'hC; #100;
A = 8'h15; B = 8'hD; #100;
A = 8'h15; B = 8'hE; #100;
A = 8'h15; B = 8'hF; #100;
A = 8'h15; B = 8'h10; #100;
A = 8'h15; B = 8'h11; #100;
A = 8'h15; B = 8'h12; #100;
A = 8'h15; B = 8'h13; #100;
A = 8'h15; B = 8'h14; #100;
A = 8'h15; B = 8'h15; #100;
A = 8'h15; B = 8'h16; #100;
A = 8'h15; B = 8'h17; #100;
A = 8'h15; B = 8'h18; #100;
A = 8'h15; B = 8'h19; #100;
A = 8'h15; B = 8'h1A; #100;
A = 8'h15; B = 8'h1B; #100;
A = 8'h15; B = 8'h1C; #100;
A = 8'h15; B = 8'h1D; #100;
A = 8'h15; B = 8'h1E; #100;
A = 8'h15; B = 8'h1F; #100;
A = 8'h15; B = 8'h20; #100;
A = 8'h15; B = 8'h21; #100;
A = 8'h15; B = 8'h22; #100;
A = 8'h15; B = 8'h23; #100;
A = 8'h15; B = 8'h24; #100;
A = 8'h15; B = 8'h25; #100;
A = 8'h15; B = 8'h26; #100;
A = 8'h15; B = 8'h27; #100;
A = 8'h15; B = 8'h28; #100;
A = 8'h15; B = 8'h29; #100;
A = 8'h15; B = 8'h2A; #100;
A = 8'h15; B = 8'h2B; #100;
A = 8'h15; B = 8'h2C; #100;
A = 8'h15; B = 8'h2D; #100;
A = 8'h15; B = 8'h2E; #100;
A = 8'h15; B = 8'h2F; #100;
A = 8'h15; B = 8'h30; #100;
A = 8'h15; B = 8'h31; #100;
A = 8'h15; B = 8'h32; #100;
A = 8'h15; B = 8'h33; #100;
A = 8'h15; B = 8'h34; #100;
A = 8'h15; B = 8'h35; #100;
A = 8'h15; B = 8'h36; #100;
A = 8'h15; B = 8'h37; #100;
A = 8'h15; B = 8'h38; #100;
A = 8'h15; B = 8'h39; #100;
A = 8'h15; B = 8'h3A; #100;
A = 8'h15; B = 8'h3B; #100;
A = 8'h15; B = 8'h3C; #100;
A = 8'h15; B = 8'h3D; #100;
A = 8'h15; B = 8'h3E; #100;
A = 8'h15; B = 8'h3F; #100;
A = 8'h15; B = 8'h40; #100;
A = 8'h15; B = 8'h41; #100;
A = 8'h15; B = 8'h42; #100;
A = 8'h15; B = 8'h43; #100;
A = 8'h15; B = 8'h44; #100;
A = 8'h15; B = 8'h45; #100;
A = 8'h15; B = 8'h46; #100;
A = 8'h15; B = 8'h47; #100;
A = 8'h15; B = 8'h48; #100;
A = 8'h15; B = 8'h49; #100;
A = 8'h15; B = 8'h4A; #100;
A = 8'h15; B = 8'h4B; #100;
A = 8'h15; B = 8'h4C; #100;
A = 8'h15; B = 8'h4D; #100;
A = 8'h15; B = 8'h4E; #100;
A = 8'h15; B = 8'h4F; #100;
A = 8'h15; B = 8'h50; #100;
A = 8'h15; B = 8'h51; #100;
A = 8'h15; B = 8'h52; #100;
A = 8'h15; B = 8'h53; #100;
A = 8'h15; B = 8'h54; #100;
A = 8'h15; B = 8'h55; #100;
A = 8'h15; B = 8'h56; #100;
A = 8'h15; B = 8'h57; #100;
A = 8'h15; B = 8'h58; #100;
A = 8'h15; B = 8'h59; #100;
A = 8'h15; B = 8'h5A; #100;
A = 8'h15; B = 8'h5B; #100;
A = 8'h15; B = 8'h5C; #100;
A = 8'h15; B = 8'h5D; #100;
A = 8'h15; B = 8'h5E; #100;
A = 8'h15; B = 8'h5F; #100;
A = 8'h15; B = 8'h60; #100;
A = 8'h15; B = 8'h61; #100;
A = 8'h15; B = 8'h62; #100;
A = 8'h15; B = 8'h63; #100;
A = 8'h15; B = 8'h64; #100;
A = 8'h15; B = 8'h65; #100;
A = 8'h15; B = 8'h66; #100;
A = 8'h15; B = 8'h67; #100;
A = 8'h15; B = 8'h68; #100;
A = 8'h15; B = 8'h69; #100;
A = 8'h15; B = 8'h6A; #100;
A = 8'h15; B = 8'h6B; #100;
A = 8'h15; B = 8'h6C; #100;
A = 8'h15; B = 8'h6D; #100;
A = 8'h15; B = 8'h6E; #100;
A = 8'h15; B = 8'h6F; #100;
A = 8'h15; B = 8'h70; #100;
A = 8'h15; B = 8'h71; #100;
A = 8'h15; B = 8'h72; #100;
A = 8'h15; B = 8'h73; #100;
A = 8'h15; B = 8'h74; #100;
A = 8'h15; B = 8'h75; #100;
A = 8'h15; B = 8'h76; #100;
A = 8'h15; B = 8'h77; #100;
A = 8'h15; B = 8'h78; #100;
A = 8'h15; B = 8'h79; #100;
A = 8'h15; B = 8'h7A; #100;
A = 8'h15; B = 8'h7B; #100;
A = 8'h15; B = 8'h7C; #100;
A = 8'h15; B = 8'h7D; #100;
A = 8'h15; B = 8'h7E; #100;
A = 8'h15; B = 8'h7F; #100;
A = 8'h15; B = 8'h80; #100;
A = 8'h15; B = 8'h81; #100;
A = 8'h15; B = 8'h82; #100;
A = 8'h15; B = 8'h83; #100;
A = 8'h15; B = 8'h84; #100;
A = 8'h15; B = 8'h85; #100;
A = 8'h15; B = 8'h86; #100;
A = 8'h15; B = 8'h87; #100;
A = 8'h15; B = 8'h88; #100;
A = 8'h15; B = 8'h89; #100;
A = 8'h15; B = 8'h8A; #100;
A = 8'h15; B = 8'h8B; #100;
A = 8'h15; B = 8'h8C; #100;
A = 8'h15; B = 8'h8D; #100;
A = 8'h15; B = 8'h8E; #100;
A = 8'h15; B = 8'h8F; #100;
A = 8'h15; B = 8'h90; #100;
A = 8'h15; B = 8'h91; #100;
A = 8'h15; B = 8'h92; #100;
A = 8'h15; B = 8'h93; #100;
A = 8'h15; B = 8'h94; #100;
A = 8'h15; B = 8'h95; #100;
A = 8'h15; B = 8'h96; #100;
A = 8'h15; B = 8'h97; #100;
A = 8'h15; B = 8'h98; #100;
A = 8'h15; B = 8'h99; #100;
A = 8'h15; B = 8'h9A; #100;
A = 8'h15; B = 8'h9B; #100;
A = 8'h15; B = 8'h9C; #100;
A = 8'h15; B = 8'h9D; #100;
A = 8'h15; B = 8'h9E; #100;
A = 8'h15; B = 8'h9F; #100;
A = 8'h15; B = 8'hA0; #100;
A = 8'h15; B = 8'hA1; #100;
A = 8'h15; B = 8'hA2; #100;
A = 8'h15; B = 8'hA3; #100;
A = 8'h15; B = 8'hA4; #100;
A = 8'h15; B = 8'hA5; #100;
A = 8'h15; B = 8'hA6; #100;
A = 8'h15; B = 8'hA7; #100;
A = 8'h15; B = 8'hA8; #100;
A = 8'h15; B = 8'hA9; #100;
A = 8'h15; B = 8'hAA; #100;
A = 8'h15; B = 8'hAB; #100;
A = 8'h15; B = 8'hAC; #100;
A = 8'h15; B = 8'hAD; #100;
A = 8'h15; B = 8'hAE; #100;
A = 8'h15; B = 8'hAF; #100;
A = 8'h15; B = 8'hB0; #100;
A = 8'h15; B = 8'hB1; #100;
A = 8'h15; B = 8'hB2; #100;
A = 8'h15; B = 8'hB3; #100;
A = 8'h15; B = 8'hB4; #100;
A = 8'h15; B = 8'hB5; #100;
A = 8'h15; B = 8'hB6; #100;
A = 8'h15; B = 8'hB7; #100;
A = 8'h15; B = 8'hB8; #100;
A = 8'h15; B = 8'hB9; #100;
A = 8'h15; B = 8'hBA; #100;
A = 8'h15; B = 8'hBB; #100;
A = 8'h15; B = 8'hBC; #100;
A = 8'h15; B = 8'hBD; #100;
A = 8'h15; B = 8'hBE; #100;
A = 8'h15; B = 8'hBF; #100;
A = 8'h15; B = 8'hC0; #100;
A = 8'h15; B = 8'hC1; #100;
A = 8'h15; B = 8'hC2; #100;
A = 8'h15; B = 8'hC3; #100;
A = 8'h15; B = 8'hC4; #100;
A = 8'h15; B = 8'hC5; #100;
A = 8'h15; B = 8'hC6; #100;
A = 8'h15; B = 8'hC7; #100;
A = 8'h15; B = 8'hC8; #100;
A = 8'h15; B = 8'hC9; #100;
A = 8'h15; B = 8'hCA; #100;
A = 8'h15; B = 8'hCB; #100;
A = 8'h15; B = 8'hCC; #100;
A = 8'h15; B = 8'hCD; #100;
A = 8'h15; B = 8'hCE; #100;
A = 8'h15; B = 8'hCF; #100;
A = 8'h15; B = 8'hD0; #100;
A = 8'h15; B = 8'hD1; #100;
A = 8'h15; B = 8'hD2; #100;
A = 8'h15; B = 8'hD3; #100;
A = 8'h15; B = 8'hD4; #100;
A = 8'h15; B = 8'hD5; #100;
A = 8'h15; B = 8'hD6; #100;
A = 8'h15; B = 8'hD7; #100;
A = 8'h15; B = 8'hD8; #100;
A = 8'h15; B = 8'hD9; #100;
A = 8'h15; B = 8'hDA; #100;
A = 8'h15; B = 8'hDB; #100;
A = 8'h15; B = 8'hDC; #100;
A = 8'h15; B = 8'hDD; #100;
A = 8'h15; B = 8'hDE; #100;
A = 8'h15; B = 8'hDF; #100;
A = 8'h15; B = 8'hE0; #100;
A = 8'h15; B = 8'hE1; #100;
A = 8'h15; B = 8'hE2; #100;
A = 8'h15; B = 8'hE3; #100;
A = 8'h15; B = 8'hE4; #100;
A = 8'h15; B = 8'hE5; #100;
A = 8'h15; B = 8'hE6; #100;
A = 8'h15; B = 8'hE7; #100;
A = 8'h15; B = 8'hE8; #100;
A = 8'h15; B = 8'hE9; #100;
A = 8'h15; B = 8'hEA; #100;
A = 8'h15; B = 8'hEB; #100;
A = 8'h15; B = 8'hEC; #100;
A = 8'h15; B = 8'hED; #100;
A = 8'h15; B = 8'hEE; #100;
A = 8'h15; B = 8'hEF; #100;
A = 8'h15; B = 8'hF0; #100;
A = 8'h15; B = 8'hF1; #100;
A = 8'h15; B = 8'hF2; #100;
A = 8'h15; B = 8'hF3; #100;
A = 8'h15; B = 8'hF4; #100;
A = 8'h15; B = 8'hF5; #100;
A = 8'h15; B = 8'hF6; #100;
A = 8'h15; B = 8'hF7; #100;
A = 8'h15; B = 8'hF8; #100;
A = 8'h15; B = 8'hF9; #100;
A = 8'h15; B = 8'hFA; #100;
A = 8'h15; B = 8'hFB; #100;
A = 8'h15; B = 8'hFC; #100;
A = 8'h15; B = 8'hFD; #100;
A = 8'h15; B = 8'hFE; #100;
A = 8'h15; B = 8'hFF; #100;
A = 8'h16; B = 8'h0; #100;
A = 8'h16; B = 8'h1; #100;
A = 8'h16; B = 8'h2; #100;
A = 8'h16; B = 8'h3; #100;
A = 8'h16; B = 8'h4; #100;
A = 8'h16; B = 8'h5; #100;
A = 8'h16; B = 8'h6; #100;
A = 8'h16; B = 8'h7; #100;
A = 8'h16; B = 8'h8; #100;
A = 8'h16; B = 8'h9; #100;
A = 8'h16; B = 8'hA; #100;
A = 8'h16; B = 8'hB; #100;
A = 8'h16; B = 8'hC; #100;
A = 8'h16; B = 8'hD; #100;
A = 8'h16; B = 8'hE; #100;
A = 8'h16; B = 8'hF; #100;
A = 8'h16; B = 8'h10; #100;
A = 8'h16; B = 8'h11; #100;
A = 8'h16; B = 8'h12; #100;
A = 8'h16; B = 8'h13; #100;
A = 8'h16; B = 8'h14; #100;
A = 8'h16; B = 8'h15; #100;
A = 8'h16; B = 8'h16; #100;
A = 8'h16; B = 8'h17; #100;
A = 8'h16; B = 8'h18; #100;
A = 8'h16; B = 8'h19; #100;
A = 8'h16; B = 8'h1A; #100;
A = 8'h16; B = 8'h1B; #100;
A = 8'h16; B = 8'h1C; #100;
A = 8'h16; B = 8'h1D; #100;
A = 8'h16; B = 8'h1E; #100;
A = 8'h16; B = 8'h1F; #100;
A = 8'h16; B = 8'h20; #100;
A = 8'h16; B = 8'h21; #100;
A = 8'h16; B = 8'h22; #100;
A = 8'h16; B = 8'h23; #100;
A = 8'h16; B = 8'h24; #100;
A = 8'h16; B = 8'h25; #100;
A = 8'h16; B = 8'h26; #100;
A = 8'h16; B = 8'h27; #100;
A = 8'h16; B = 8'h28; #100;
A = 8'h16; B = 8'h29; #100;
A = 8'h16; B = 8'h2A; #100;
A = 8'h16; B = 8'h2B; #100;
A = 8'h16; B = 8'h2C; #100;
A = 8'h16; B = 8'h2D; #100;
A = 8'h16; B = 8'h2E; #100;
A = 8'h16; B = 8'h2F; #100;
A = 8'h16; B = 8'h30; #100;
A = 8'h16; B = 8'h31; #100;
A = 8'h16; B = 8'h32; #100;
A = 8'h16; B = 8'h33; #100;
A = 8'h16; B = 8'h34; #100;
A = 8'h16; B = 8'h35; #100;
A = 8'h16; B = 8'h36; #100;
A = 8'h16; B = 8'h37; #100;
A = 8'h16; B = 8'h38; #100;
A = 8'h16; B = 8'h39; #100;
A = 8'h16; B = 8'h3A; #100;
A = 8'h16; B = 8'h3B; #100;
A = 8'h16; B = 8'h3C; #100;
A = 8'h16; B = 8'h3D; #100;
A = 8'h16; B = 8'h3E; #100;
A = 8'h16; B = 8'h3F; #100;
A = 8'h16; B = 8'h40; #100;
A = 8'h16; B = 8'h41; #100;
A = 8'h16; B = 8'h42; #100;
A = 8'h16; B = 8'h43; #100;
A = 8'h16; B = 8'h44; #100;
A = 8'h16; B = 8'h45; #100;
A = 8'h16; B = 8'h46; #100;
A = 8'h16; B = 8'h47; #100;
A = 8'h16; B = 8'h48; #100;
A = 8'h16; B = 8'h49; #100;
A = 8'h16; B = 8'h4A; #100;
A = 8'h16; B = 8'h4B; #100;
A = 8'h16; B = 8'h4C; #100;
A = 8'h16; B = 8'h4D; #100;
A = 8'h16; B = 8'h4E; #100;
A = 8'h16; B = 8'h4F; #100;
A = 8'h16; B = 8'h50; #100;
A = 8'h16; B = 8'h51; #100;
A = 8'h16; B = 8'h52; #100;
A = 8'h16; B = 8'h53; #100;
A = 8'h16; B = 8'h54; #100;
A = 8'h16; B = 8'h55; #100;
A = 8'h16; B = 8'h56; #100;
A = 8'h16; B = 8'h57; #100;
A = 8'h16; B = 8'h58; #100;
A = 8'h16; B = 8'h59; #100;
A = 8'h16; B = 8'h5A; #100;
A = 8'h16; B = 8'h5B; #100;
A = 8'h16; B = 8'h5C; #100;
A = 8'h16; B = 8'h5D; #100;
A = 8'h16; B = 8'h5E; #100;
A = 8'h16; B = 8'h5F; #100;
A = 8'h16; B = 8'h60; #100;
A = 8'h16; B = 8'h61; #100;
A = 8'h16; B = 8'h62; #100;
A = 8'h16; B = 8'h63; #100;
A = 8'h16; B = 8'h64; #100;
A = 8'h16; B = 8'h65; #100;
A = 8'h16; B = 8'h66; #100;
A = 8'h16; B = 8'h67; #100;
A = 8'h16; B = 8'h68; #100;
A = 8'h16; B = 8'h69; #100;
A = 8'h16; B = 8'h6A; #100;
A = 8'h16; B = 8'h6B; #100;
A = 8'h16; B = 8'h6C; #100;
A = 8'h16; B = 8'h6D; #100;
A = 8'h16; B = 8'h6E; #100;
A = 8'h16; B = 8'h6F; #100;
A = 8'h16; B = 8'h70; #100;
A = 8'h16; B = 8'h71; #100;
A = 8'h16; B = 8'h72; #100;
A = 8'h16; B = 8'h73; #100;
A = 8'h16; B = 8'h74; #100;
A = 8'h16; B = 8'h75; #100;
A = 8'h16; B = 8'h76; #100;
A = 8'h16; B = 8'h77; #100;
A = 8'h16; B = 8'h78; #100;
A = 8'h16; B = 8'h79; #100;
A = 8'h16; B = 8'h7A; #100;
A = 8'h16; B = 8'h7B; #100;
A = 8'h16; B = 8'h7C; #100;
A = 8'h16; B = 8'h7D; #100;
A = 8'h16; B = 8'h7E; #100;
A = 8'h16; B = 8'h7F; #100;
A = 8'h16; B = 8'h80; #100;
A = 8'h16; B = 8'h81; #100;
A = 8'h16; B = 8'h82; #100;
A = 8'h16; B = 8'h83; #100;
A = 8'h16; B = 8'h84; #100;
A = 8'h16; B = 8'h85; #100;
A = 8'h16; B = 8'h86; #100;
A = 8'h16; B = 8'h87; #100;
A = 8'h16; B = 8'h88; #100;
A = 8'h16; B = 8'h89; #100;
A = 8'h16; B = 8'h8A; #100;
A = 8'h16; B = 8'h8B; #100;
A = 8'h16; B = 8'h8C; #100;
A = 8'h16; B = 8'h8D; #100;
A = 8'h16; B = 8'h8E; #100;
A = 8'h16; B = 8'h8F; #100;
A = 8'h16; B = 8'h90; #100;
A = 8'h16; B = 8'h91; #100;
A = 8'h16; B = 8'h92; #100;
A = 8'h16; B = 8'h93; #100;
A = 8'h16; B = 8'h94; #100;
A = 8'h16; B = 8'h95; #100;
A = 8'h16; B = 8'h96; #100;
A = 8'h16; B = 8'h97; #100;
A = 8'h16; B = 8'h98; #100;
A = 8'h16; B = 8'h99; #100;
A = 8'h16; B = 8'h9A; #100;
A = 8'h16; B = 8'h9B; #100;
A = 8'h16; B = 8'h9C; #100;
A = 8'h16; B = 8'h9D; #100;
A = 8'h16; B = 8'h9E; #100;
A = 8'h16; B = 8'h9F; #100;
A = 8'h16; B = 8'hA0; #100;
A = 8'h16; B = 8'hA1; #100;
A = 8'h16; B = 8'hA2; #100;
A = 8'h16; B = 8'hA3; #100;
A = 8'h16; B = 8'hA4; #100;
A = 8'h16; B = 8'hA5; #100;
A = 8'h16; B = 8'hA6; #100;
A = 8'h16; B = 8'hA7; #100;
A = 8'h16; B = 8'hA8; #100;
A = 8'h16; B = 8'hA9; #100;
A = 8'h16; B = 8'hAA; #100;
A = 8'h16; B = 8'hAB; #100;
A = 8'h16; B = 8'hAC; #100;
A = 8'h16; B = 8'hAD; #100;
A = 8'h16; B = 8'hAE; #100;
A = 8'h16; B = 8'hAF; #100;
A = 8'h16; B = 8'hB0; #100;
A = 8'h16; B = 8'hB1; #100;
A = 8'h16; B = 8'hB2; #100;
A = 8'h16; B = 8'hB3; #100;
A = 8'h16; B = 8'hB4; #100;
A = 8'h16; B = 8'hB5; #100;
A = 8'h16; B = 8'hB6; #100;
A = 8'h16; B = 8'hB7; #100;
A = 8'h16; B = 8'hB8; #100;
A = 8'h16; B = 8'hB9; #100;
A = 8'h16; B = 8'hBA; #100;
A = 8'h16; B = 8'hBB; #100;
A = 8'h16; B = 8'hBC; #100;
A = 8'h16; B = 8'hBD; #100;
A = 8'h16; B = 8'hBE; #100;
A = 8'h16; B = 8'hBF; #100;
A = 8'h16; B = 8'hC0; #100;
A = 8'h16; B = 8'hC1; #100;
A = 8'h16; B = 8'hC2; #100;
A = 8'h16; B = 8'hC3; #100;
A = 8'h16; B = 8'hC4; #100;
A = 8'h16; B = 8'hC5; #100;
A = 8'h16; B = 8'hC6; #100;
A = 8'h16; B = 8'hC7; #100;
A = 8'h16; B = 8'hC8; #100;
A = 8'h16; B = 8'hC9; #100;
A = 8'h16; B = 8'hCA; #100;
A = 8'h16; B = 8'hCB; #100;
A = 8'h16; B = 8'hCC; #100;
A = 8'h16; B = 8'hCD; #100;
A = 8'h16; B = 8'hCE; #100;
A = 8'h16; B = 8'hCF; #100;
A = 8'h16; B = 8'hD0; #100;
A = 8'h16; B = 8'hD1; #100;
A = 8'h16; B = 8'hD2; #100;
A = 8'h16; B = 8'hD3; #100;
A = 8'h16; B = 8'hD4; #100;
A = 8'h16; B = 8'hD5; #100;
A = 8'h16; B = 8'hD6; #100;
A = 8'h16; B = 8'hD7; #100;
A = 8'h16; B = 8'hD8; #100;
A = 8'h16; B = 8'hD9; #100;
A = 8'h16; B = 8'hDA; #100;
A = 8'h16; B = 8'hDB; #100;
A = 8'h16; B = 8'hDC; #100;
A = 8'h16; B = 8'hDD; #100;
A = 8'h16; B = 8'hDE; #100;
A = 8'h16; B = 8'hDF; #100;
A = 8'h16; B = 8'hE0; #100;
A = 8'h16; B = 8'hE1; #100;
A = 8'h16; B = 8'hE2; #100;
A = 8'h16; B = 8'hE3; #100;
A = 8'h16; B = 8'hE4; #100;
A = 8'h16; B = 8'hE5; #100;
A = 8'h16; B = 8'hE6; #100;
A = 8'h16; B = 8'hE7; #100;
A = 8'h16; B = 8'hE8; #100;
A = 8'h16; B = 8'hE9; #100;
A = 8'h16; B = 8'hEA; #100;
A = 8'h16; B = 8'hEB; #100;
A = 8'h16; B = 8'hEC; #100;
A = 8'h16; B = 8'hED; #100;
A = 8'h16; B = 8'hEE; #100;
A = 8'h16; B = 8'hEF; #100;
A = 8'h16; B = 8'hF0; #100;
A = 8'h16; B = 8'hF1; #100;
A = 8'h16; B = 8'hF2; #100;
A = 8'h16; B = 8'hF3; #100;
A = 8'h16; B = 8'hF4; #100;
A = 8'h16; B = 8'hF5; #100;
A = 8'h16; B = 8'hF6; #100;
A = 8'h16; B = 8'hF7; #100;
A = 8'h16; B = 8'hF8; #100;
A = 8'h16; B = 8'hF9; #100;
A = 8'h16; B = 8'hFA; #100;
A = 8'h16; B = 8'hFB; #100;
A = 8'h16; B = 8'hFC; #100;
A = 8'h16; B = 8'hFD; #100;
A = 8'h16; B = 8'hFE; #100;
A = 8'h16; B = 8'hFF; #100;
A = 8'h17; B = 8'h0; #100;
A = 8'h17; B = 8'h1; #100;
A = 8'h17; B = 8'h2; #100;
A = 8'h17; B = 8'h3; #100;
A = 8'h17; B = 8'h4; #100;
A = 8'h17; B = 8'h5; #100;
A = 8'h17; B = 8'h6; #100;
A = 8'h17; B = 8'h7; #100;
A = 8'h17; B = 8'h8; #100;
A = 8'h17; B = 8'h9; #100;
A = 8'h17; B = 8'hA; #100;
A = 8'h17; B = 8'hB; #100;
A = 8'h17; B = 8'hC; #100;
A = 8'h17; B = 8'hD; #100;
A = 8'h17; B = 8'hE; #100;
A = 8'h17; B = 8'hF; #100;
A = 8'h17; B = 8'h10; #100;
A = 8'h17; B = 8'h11; #100;
A = 8'h17; B = 8'h12; #100;
A = 8'h17; B = 8'h13; #100;
A = 8'h17; B = 8'h14; #100;
A = 8'h17; B = 8'h15; #100;
A = 8'h17; B = 8'h16; #100;
A = 8'h17; B = 8'h17; #100;
A = 8'h17; B = 8'h18; #100;
A = 8'h17; B = 8'h19; #100;
A = 8'h17; B = 8'h1A; #100;
A = 8'h17; B = 8'h1B; #100;
A = 8'h17; B = 8'h1C; #100;
A = 8'h17; B = 8'h1D; #100;
A = 8'h17; B = 8'h1E; #100;
A = 8'h17; B = 8'h1F; #100;
A = 8'h17; B = 8'h20; #100;
A = 8'h17; B = 8'h21; #100;
A = 8'h17; B = 8'h22; #100;
A = 8'h17; B = 8'h23; #100;
A = 8'h17; B = 8'h24; #100;
A = 8'h17; B = 8'h25; #100;
A = 8'h17; B = 8'h26; #100;
A = 8'h17; B = 8'h27; #100;
A = 8'h17; B = 8'h28; #100;
A = 8'h17; B = 8'h29; #100;
A = 8'h17; B = 8'h2A; #100;
A = 8'h17; B = 8'h2B; #100;
A = 8'h17; B = 8'h2C; #100;
A = 8'h17; B = 8'h2D; #100;
A = 8'h17; B = 8'h2E; #100;
A = 8'h17; B = 8'h2F; #100;
A = 8'h17; B = 8'h30; #100;
A = 8'h17; B = 8'h31; #100;
A = 8'h17; B = 8'h32; #100;
A = 8'h17; B = 8'h33; #100;
A = 8'h17; B = 8'h34; #100;
A = 8'h17; B = 8'h35; #100;
A = 8'h17; B = 8'h36; #100;
A = 8'h17; B = 8'h37; #100;
A = 8'h17; B = 8'h38; #100;
A = 8'h17; B = 8'h39; #100;
A = 8'h17; B = 8'h3A; #100;
A = 8'h17; B = 8'h3B; #100;
A = 8'h17; B = 8'h3C; #100;
A = 8'h17; B = 8'h3D; #100;
A = 8'h17; B = 8'h3E; #100;
A = 8'h17; B = 8'h3F; #100;
A = 8'h17; B = 8'h40; #100;
A = 8'h17; B = 8'h41; #100;
A = 8'h17; B = 8'h42; #100;
A = 8'h17; B = 8'h43; #100;
A = 8'h17; B = 8'h44; #100;
A = 8'h17; B = 8'h45; #100;
A = 8'h17; B = 8'h46; #100;
A = 8'h17; B = 8'h47; #100;
A = 8'h17; B = 8'h48; #100;
A = 8'h17; B = 8'h49; #100;
A = 8'h17; B = 8'h4A; #100;
A = 8'h17; B = 8'h4B; #100;
A = 8'h17; B = 8'h4C; #100;
A = 8'h17; B = 8'h4D; #100;
A = 8'h17; B = 8'h4E; #100;
A = 8'h17; B = 8'h4F; #100;
A = 8'h17; B = 8'h50; #100;
A = 8'h17; B = 8'h51; #100;
A = 8'h17; B = 8'h52; #100;
A = 8'h17; B = 8'h53; #100;
A = 8'h17; B = 8'h54; #100;
A = 8'h17; B = 8'h55; #100;
A = 8'h17; B = 8'h56; #100;
A = 8'h17; B = 8'h57; #100;
A = 8'h17; B = 8'h58; #100;
A = 8'h17; B = 8'h59; #100;
A = 8'h17; B = 8'h5A; #100;
A = 8'h17; B = 8'h5B; #100;
A = 8'h17; B = 8'h5C; #100;
A = 8'h17; B = 8'h5D; #100;
A = 8'h17; B = 8'h5E; #100;
A = 8'h17; B = 8'h5F; #100;
A = 8'h17; B = 8'h60; #100;
A = 8'h17; B = 8'h61; #100;
A = 8'h17; B = 8'h62; #100;
A = 8'h17; B = 8'h63; #100;
A = 8'h17; B = 8'h64; #100;
A = 8'h17; B = 8'h65; #100;
A = 8'h17; B = 8'h66; #100;
A = 8'h17; B = 8'h67; #100;
A = 8'h17; B = 8'h68; #100;
A = 8'h17; B = 8'h69; #100;
A = 8'h17; B = 8'h6A; #100;
A = 8'h17; B = 8'h6B; #100;
A = 8'h17; B = 8'h6C; #100;
A = 8'h17; B = 8'h6D; #100;
A = 8'h17; B = 8'h6E; #100;
A = 8'h17; B = 8'h6F; #100;
A = 8'h17; B = 8'h70; #100;
A = 8'h17; B = 8'h71; #100;
A = 8'h17; B = 8'h72; #100;
A = 8'h17; B = 8'h73; #100;
A = 8'h17; B = 8'h74; #100;
A = 8'h17; B = 8'h75; #100;
A = 8'h17; B = 8'h76; #100;
A = 8'h17; B = 8'h77; #100;
A = 8'h17; B = 8'h78; #100;
A = 8'h17; B = 8'h79; #100;
A = 8'h17; B = 8'h7A; #100;
A = 8'h17; B = 8'h7B; #100;
A = 8'h17; B = 8'h7C; #100;
A = 8'h17; B = 8'h7D; #100;
A = 8'h17; B = 8'h7E; #100;
A = 8'h17; B = 8'h7F; #100;
A = 8'h17; B = 8'h80; #100;
A = 8'h17; B = 8'h81; #100;
A = 8'h17; B = 8'h82; #100;
A = 8'h17; B = 8'h83; #100;
A = 8'h17; B = 8'h84; #100;
A = 8'h17; B = 8'h85; #100;
A = 8'h17; B = 8'h86; #100;
A = 8'h17; B = 8'h87; #100;
A = 8'h17; B = 8'h88; #100;
A = 8'h17; B = 8'h89; #100;
A = 8'h17; B = 8'h8A; #100;
A = 8'h17; B = 8'h8B; #100;
A = 8'h17; B = 8'h8C; #100;
A = 8'h17; B = 8'h8D; #100;
A = 8'h17; B = 8'h8E; #100;
A = 8'h17; B = 8'h8F; #100;
A = 8'h17; B = 8'h90; #100;
A = 8'h17; B = 8'h91; #100;
A = 8'h17; B = 8'h92; #100;
A = 8'h17; B = 8'h93; #100;
A = 8'h17; B = 8'h94; #100;
A = 8'h17; B = 8'h95; #100;
A = 8'h17; B = 8'h96; #100;
A = 8'h17; B = 8'h97; #100;
A = 8'h17; B = 8'h98; #100;
A = 8'h17; B = 8'h99; #100;
A = 8'h17; B = 8'h9A; #100;
A = 8'h17; B = 8'h9B; #100;
A = 8'h17; B = 8'h9C; #100;
A = 8'h17; B = 8'h9D; #100;
A = 8'h17; B = 8'h9E; #100;
A = 8'h17; B = 8'h9F; #100;
A = 8'h17; B = 8'hA0; #100;
A = 8'h17; B = 8'hA1; #100;
A = 8'h17; B = 8'hA2; #100;
A = 8'h17; B = 8'hA3; #100;
A = 8'h17; B = 8'hA4; #100;
A = 8'h17; B = 8'hA5; #100;
A = 8'h17; B = 8'hA6; #100;
A = 8'h17; B = 8'hA7; #100;
A = 8'h17; B = 8'hA8; #100;
A = 8'h17; B = 8'hA9; #100;
A = 8'h17; B = 8'hAA; #100;
A = 8'h17; B = 8'hAB; #100;
A = 8'h17; B = 8'hAC; #100;
A = 8'h17; B = 8'hAD; #100;
A = 8'h17; B = 8'hAE; #100;
A = 8'h17; B = 8'hAF; #100;
A = 8'h17; B = 8'hB0; #100;
A = 8'h17; B = 8'hB1; #100;
A = 8'h17; B = 8'hB2; #100;
A = 8'h17; B = 8'hB3; #100;
A = 8'h17; B = 8'hB4; #100;
A = 8'h17; B = 8'hB5; #100;
A = 8'h17; B = 8'hB6; #100;
A = 8'h17; B = 8'hB7; #100;
A = 8'h17; B = 8'hB8; #100;
A = 8'h17; B = 8'hB9; #100;
A = 8'h17; B = 8'hBA; #100;
A = 8'h17; B = 8'hBB; #100;
A = 8'h17; B = 8'hBC; #100;
A = 8'h17; B = 8'hBD; #100;
A = 8'h17; B = 8'hBE; #100;
A = 8'h17; B = 8'hBF; #100;
A = 8'h17; B = 8'hC0; #100;
A = 8'h17; B = 8'hC1; #100;
A = 8'h17; B = 8'hC2; #100;
A = 8'h17; B = 8'hC3; #100;
A = 8'h17; B = 8'hC4; #100;
A = 8'h17; B = 8'hC5; #100;
A = 8'h17; B = 8'hC6; #100;
A = 8'h17; B = 8'hC7; #100;
A = 8'h17; B = 8'hC8; #100;
A = 8'h17; B = 8'hC9; #100;
A = 8'h17; B = 8'hCA; #100;
A = 8'h17; B = 8'hCB; #100;
A = 8'h17; B = 8'hCC; #100;
A = 8'h17; B = 8'hCD; #100;
A = 8'h17; B = 8'hCE; #100;
A = 8'h17; B = 8'hCF; #100;
A = 8'h17; B = 8'hD0; #100;
A = 8'h17; B = 8'hD1; #100;
A = 8'h17; B = 8'hD2; #100;
A = 8'h17; B = 8'hD3; #100;
A = 8'h17; B = 8'hD4; #100;
A = 8'h17; B = 8'hD5; #100;
A = 8'h17; B = 8'hD6; #100;
A = 8'h17; B = 8'hD7; #100;
A = 8'h17; B = 8'hD8; #100;
A = 8'h17; B = 8'hD9; #100;
A = 8'h17; B = 8'hDA; #100;
A = 8'h17; B = 8'hDB; #100;
A = 8'h17; B = 8'hDC; #100;
A = 8'h17; B = 8'hDD; #100;
A = 8'h17; B = 8'hDE; #100;
A = 8'h17; B = 8'hDF; #100;
A = 8'h17; B = 8'hE0; #100;
A = 8'h17; B = 8'hE1; #100;
A = 8'h17; B = 8'hE2; #100;
A = 8'h17; B = 8'hE3; #100;
A = 8'h17; B = 8'hE4; #100;
A = 8'h17; B = 8'hE5; #100;
A = 8'h17; B = 8'hE6; #100;
A = 8'h17; B = 8'hE7; #100;
A = 8'h17; B = 8'hE8; #100;
A = 8'h17; B = 8'hE9; #100;
A = 8'h17; B = 8'hEA; #100;
A = 8'h17; B = 8'hEB; #100;
A = 8'h17; B = 8'hEC; #100;
A = 8'h17; B = 8'hED; #100;
A = 8'h17; B = 8'hEE; #100;
A = 8'h17; B = 8'hEF; #100;
A = 8'h17; B = 8'hF0; #100;
A = 8'h17; B = 8'hF1; #100;
A = 8'h17; B = 8'hF2; #100;
A = 8'h17; B = 8'hF3; #100;
A = 8'h17; B = 8'hF4; #100;
A = 8'h17; B = 8'hF5; #100;
A = 8'h17; B = 8'hF6; #100;
A = 8'h17; B = 8'hF7; #100;
A = 8'h17; B = 8'hF8; #100;
A = 8'h17; B = 8'hF9; #100;
A = 8'h17; B = 8'hFA; #100;
A = 8'h17; B = 8'hFB; #100;
A = 8'h17; B = 8'hFC; #100;
A = 8'h17; B = 8'hFD; #100;
A = 8'h17; B = 8'hFE; #100;
A = 8'h17; B = 8'hFF; #100;
A = 8'h18; B = 8'h0; #100;
A = 8'h18; B = 8'h1; #100;
A = 8'h18; B = 8'h2; #100;
A = 8'h18; B = 8'h3; #100;
A = 8'h18; B = 8'h4; #100;
A = 8'h18; B = 8'h5; #100;
A = 8'h18; B = 8'h6; #100;
A = 8'h18; B = 8'h7; #100;
A = 8'h18; B = 8'h8; #100;
A = 8'h18; B = 8'h9; #100;
A = 8'h18; B = 8'hA; #100;
A = 8'h18; B = 8'hB; #100;
A = 8'h18; B = 8'hC; #100;
A = 8'h18; B = 8'hD; #100;
A = 8'h18; B = 8'hE; #100;
A = 8'h18; B = 8'hF; #100;
A = 8'h18; B = 8'h10; #100;
A = 8'h18; B = 8'h11; #100;
A = 8'h18; B = 8'h12; #100;
A = 8'h18; B = 8'h13; #100;
A = 8'h18; B = 8'h14; #100;
A = 8'h18; B = 8'h15; #100;
A = 8'h18; B = 8'h16; #100;
A = 8'h18; B = 8'h17; #100;
A = 8'h18; B = 8'h18; #100;
A = 8'h18; B = 8'h19; #100;
A = 8'h18; B = 8'h1A; #100;
A = 8'h18; B = 8'h1B; #100;
A = 8'h18; B = 8'h1C; #100;
A = 8'h18; B = 8'h1D; #100;
A = 8'h18; B = 8'h1E; #100;
A = 8'h18; B = 8'h1F; #100;
A = 8'h18; B = 8'h20; #100;
A = 8'h18; B = 8'h21; #100;
A = 8'h18; B = 8'h22; #100;
A = 8'h18; B = 8'h23; #100;
A = 8'h18; B = 8'h24; #100;
A = 8'h18; B = 8'h25; #100;
A = 8'h18; B = 8'h26; #100;
A = 8'h18; B = 8'h27; #100;
A = 8'h18; B = 8'h28; #100;
A = 8'h18; B = 8'h29; #100;
A = 8'h18; B = 8'h2A; #100;
A = 8'h18; B = 8'h2B; #100;
A = 8'h18; B = 8'h2C; #100;
A = 8'h18; B = 8'h2D; #100;
A = 8'h18; B = 8'h2E; #100;
A = 8'h18; B = 8'h2F; #100;
A = 8'h18; B = 8'h30; #100;
A = 8'h18; B = 8'h31; #100;
A = 8'h18; B = 8'h32; #100;
A = 8'h18; B = 8'h33; #100;
A = 8'h18; B = 8'h34; #100;
A = 8'h18; B = 8'h35; #100;
A = 8'h18; B = 8'h36; #100;
A = 8'h18; B = 8'h37; #100;
A = 8'h18; B = 8'h38; #100;
A = 8'h18; B = 8'h39; #100;
A = 8'h18; B = 8'h3A; #100;
A = 8'h18; B = 8'h3B; #100;
A = 8'h18; B = 8'h3C; #100;
A = 8'h18; B = 8'h3D; #100;
A = 8'h18; B = 8'h3E; #100;
A = 8'h18; B = 8'h3F; #100;
A = 8'h18; B = 8'h40; #100;
A = 8'h18; B = 8'h41; #100;
A = 8'h18; B = 8'h42; #100;
A = 8'h18; B = 8'h43; #100;
A = 8'h18; B = 8'h44; #100;
A = 8'h18; B = 8'h45; #100;
A = 8'h18; B = 8'h46; #100;
A = 8'h18; B = 8'h47; #100;
A = 8'h18; B = 8'h48; #100;
A = 8'h18; B = 8'h49; #100;
A = 8'h18; B = 8'h4A; #100;
A = 8'h18; B = 8'h4B; #100;
A = 8'h18; B = 8'h4C; #100;
A = 8'h18; B = 8'h4D; #100;
A = 8'h18; B = 8'h4E; #100;
A = 8'h18; B = 8'h4F; #100;
A = 8'h18; B = 8'h50; #100;
A = 8'h18; B = 8'h51; #100;
A = 8'h18; B = 8'h52; #100;
A = 8'h18; B = 8'h53; #100;
A = 8'h18; B = 8'h54; #100;
A = 8'h18; B = 8'h55; #100;
A = 8'h18; B = 8'h56; #100;
A = 8'h18; B = 8'h57; #100;
A = 8'h18; B = 8'h58; #100;
A = 8'h18; B = 8'h59; #100;
A = 8'h18; B = 8'h5A; #100;
A = 8'h18; B = 8'h5B; #100;
A = 8'h18; B = 8'h5C; #100;
A = 8'h18; B = 8'h5D; #100;
A = 8'h18; B = 8'h5E; #100;
A = 8'h18; B = 8'h5F; #100;
A = 8'h18; B = 8'h60; #100;
A = 8'h18; B = 8'h61; #100;
A = 8'h18; B = 8'h62; #100;
A = 8'h18; B = 8'h63; #100;
A = 8'h18; B = 8'h64; #100;
A = 8'h18; B = 8'h65; #100;
A = 8'h18; B = 8'h66; #100;
A = 8'h18; B = 8'h67; #100;
A = 8'h18; B = 8'h68; #100;
A = 8'h18; B = 8'h69; #100;
A = 8'h18; B = 8'h6A; #100;
A = 8'h18; B = 8'h6B; #100;
A = 8'h18; B = 8'h6C; #100;
A = 8'h18; B = 8'h6D; #100;
A = 8'h18; B = 8'h6E; #100;
A = 8'h18; B = 8'h6F; #100;
A = 8'h18; B = 8'h70; #100;
A = 8'h18; B = 8'h71; #100;
A = 8'h18; B = 8'h72; #100;
A = 8'h18; B = 8'h73; #100;
A = 8'h18; B = 8'h74; #100;
A = 8'h18; B = 8'h75; #100;
A = 8'h18; B = 8'h76; #100;
A = 8'h18; B = 8'h77; #100;
A = 8'h18; B = 8'h78; #100;
A = 8'h18; B = 8'h79; #100;
A = 8'h18; B = 8'h7A; #100;
A = 8'h18; B = 8'h7B; #100;
A = 8'h18; B = 8'h7C; #100;
A = 8'h18; B = 8'h7D; #100;
A = 8'h18; B = 8'h7E; #100;
A = 8'h18; B = 8'h7F; #100;
A = 8'h18; B = 8'h80; #100;
A = 8'h18; B = 8'h81; #100;
A = 8'h18; B = 8'h82; #100;
A = 8'h18; B = 8'h83; #100;
A = 8'h18; B = 8'h84; #100;
A = 8'h18; B = 8'h85; #100;
A = 8'h18; B = 8'h86; #100;
A = 8'h18; B = 8'h87; #100;
A = 8'h18; B = 8'h88; #100;
A = 8'h18; B = 8'h89; #100;
A = 8'h18; B = 8'h8A; #100;
A = 8'h18; B = 8'h8B; #100;
A = 8'h18; B = 8'h8C; #100;
A = 8'h18; B = 8'h8D; #100;
A = 8'h18; B = 8'h8E; #100;
A = 8'h18; B = 8'h8F; #100;
A = 8'h18; B = 8'h90; #100;
A = 8'h18; B = 8'h91; #100;
A = 8'h18; B = 8'h92; #100;
A = 8'h18; B = 8'h93; #100;
A = 8'h18; B = 8'h94; #100;
A = 8'h18; B = 8'h95; #100;
A = 8'h18; B = 8'h96; #100;
A = 8'h18; B = 8'h97; #100;
A = 8'h18; B = 8'h98; #100;
A = 8'h18; B = 8'h99; #100;
A = 8'h18; B = 8'h9A; #100;
A = 8'h18; B = 8'h9B; #100;
A = 8'h18; B = 8'h9C; #100;
A = 8'h18; B = 8'h9D; #100;
A = 8'h18; B = 8'h9E; #100;
A = 8'h18; B = 8'h9F; #100;
A = 8'h18; B = 8'hA0; #100;
A = 8'h18; B = 8'hA1; #100;
A = 8'h18; B = 8'hA2; #100;
A = 8'h18; B = 8'hA3; #100;
A = 8'h18; B = 8'hA4; #100;
A = 8'h18; B = 8'hA5; #100;
A = 8'h18; B = 8'hA6; #100;
A = 8'h18; B = 8'hA7; #100;
A = 8'h18; B = 8'hA8; #100;
A = 8'h18; B = 8'hA9; #100;
A = 8'h18; B = 8'hAA; #100;
A = 8'h18; B = 8'hAB; #100;
A = 8'h18; B = 8'hAC; #100;
A = 8'h18; B = 8'hAD; #100;
A = 8'h18; B = 8'hAE; #100;
A = 8'h18; B = 8'hAF; #100;
A = 8'h18; B = 8'hB0; #100;
A = 8'h18; B = 8'hB1; #100;
A = 8'h18; B = 8'hB2; #100;
A = 8'h18; B = 8'hB3; #100;
A = 8'h18; B = 8'hB4; #100;
A = 8'h18; B = 8'hB5; #100;
A = 8'h18; B = 8'hB6; #100;
A = 8'h18; B = 8'hB7; #100;
A = 8'h18; B = 8'hB8; #100;
A = 8'h18; B = 8'hB9; #100;
A = 8'h18; B = 8'hBA; #100;
A = 8'h18; B = 8'hBB; #100;
A = 8'h18; B = 8'hBC; #100;
A = 8'h18; B = 8'hBD; #100;
A = 8'h18; B = 8'hBE; #100;
A = 8'h18; B = 8'hBF; #100;
A = 8'h18; B = 8'hC0; #100;
A = 8'h18; B = 8'hC1; #100;
A = 8'h18; B = 8'hC2; #100;
A = 8'h18; B = 8'hC3; #100;
A = 8'h18; B = 8'hC4; #100;
A = 8'h18; B = 8'hC5; #100;
A = 8'h18; B = 8'hC6; #100;
A = 8'h18; B = 8'hC7; #100;
A = 8'h18; B = 8'hC8; #100;
A = 8'h18; B = 8'hC9; #100;
A = 8'h18; B = 8'hCA; #100;
A = 8'h18; B = 8'hCB; #100;
A = 8'h18; B = 8'hCC; #100;
A = 8'h18; B = 8'hCD; #100;
A = 8'h18; B = 8'hCE; #100;
A = 8'h18; B = 8'hCF; #100;
A = 8'h18; B = 8'hD0; #100;
A = 8'h18; B = 8'hD1; #100;
A = 8'h18; B = 8'hD2; #100;
A = 8'h18; B = 8'hD3; #100;
A = 8'h18; B = 8'hD4; #100;
A = 8'h18; B = 8'hD5; #100;
A = 8'h18; B = 8'hD6; #100;
A = 8'h18; B = 8'hD7; #100;
A = 8'h18; B = 8'hD8; #100;
A = 8'h18; B = 8'hD9; #100;
A = 8'h18; B = 8'hDA; #100;
A = 8'h18; B = 8'hDB; #100;
A = 8'h18; B = 8'hDC; #100;
A = 8'h18; B = 8'hDD; #100;
A = 8'h18; B = 8'hDE; #100;
A = 8'h18; B = 8'hDF; #100;
A = 8'h18; B = 8'hE0; #100;
A = 8'h18; B = 8'hE1; #100;
A = 8'h18; B = 8'hE2; #100;
A = 8'h18; B = 8'hE3; #100;
A = 8'h18; B = 8'hE4; #100;
A = 8'h18; B = 8'hE5; #100;
A = 8'h18; B = 8'hE6; #100;
A = 8'h18; B = 8'hE7; #100;
A = 8'h18; B = 8'hE8; #100;
A = 8'h18; B = 8'hE9; #100;
A = 8'h18; B = 8'hEA; #100;
A = 8'h18; B = 8'hEB; #100;
A = 8'h18; B = 8'hEC; #100;
A = 8'h18; B = 8'hED; #100;
A = 8'h18; B = 8'hEE; #100;
A = 8'h18; B = 8'hEF; #100;
A = 8'h18; B = 8'hF0; #100;
A = 8'h18; B = 8'hF1; #100;
A = 8'h18; B = 8'hF2; #100;
A = 8'h18; B = 8'hF3; #100;
A = 8'h18; B = 8'hF4; #100;
A = 8'h18; B = 8'hF5; #100;
A = 8'h18; B = 8'hF6; #100;
A = 8'h18; B = 8'hF7; #100;
A = 8'h18; B = 8'hF8; #100;
A = 8'h18; B = 8'hF9; #100;
A = 8'h18; B = 8'hFA; #100;
A = 8'h18; B = 8'hFB; #100;
A = 8'h18; B = 8'hFC; #100;
A = 8'h18; B = 8'hFD; #100;
A = 8'h18; B = 8'hFE; #100;
A = 8'h18; B = 8'hFF; #100;
A = 8'h19; B = 8'h0; #100;
A = 8'h19; B = 8'h1; #100;
A = 8'h19; B = 8'h2; #100;
A = 8'h19; B = 8'h3; #100;
A = 8'h19; B = 8'h4; #100;
A = 8'h19; B = 8'h5; #100;
A = 8'h19; B = 8'h6; #100;
A = 8'h19; B = 8'h7; #100;
A = 8'h19; B = 8'h8; #100;
A = 8'h19; B = 8'h9; #100;
A = 8'h19; B = 8'hA; #100;
A = 8'h19; B = 8'hB; #100;
A = 8'h19; B = 8'hC; #100;
A = 8'h19; B = 8'hD; #100;
A = 8'h19; B = 8'hE; #100;
A = 8'h19; B = 8'hF; #100;
A = 8'h19; B = 8'h10; #100;
A = 8'h19; B = 8'h11; #100;
A = 8'h19; B = 8'h12; #100;
A = 8'h19; B = 8'h13; #100;
A = 8'h19; B = 8'h14; #100;
A = 8'h19; B = 8'h15; #100;
A = 8'h19; B = 8'h16; #100;
A = 8'h19; B = 8'h17; #100;
A = 8'h19; B = 8'h18; #100;
A = 8'h19; B = 8'h19; #100;
A = 8'h19; B = 8'h1A; #100;
A = 8'h19; B = 8'h1B; #100;
A = 8'h19; B = 8'h1C; #100;
A = 8'h19; B = 8'h1D; #100;
A = 8'h19; B = 8'h1E; #100;
A = 8'h19; B = 8'h1F; #100;
A = 8'h19; B = 8'h20; #100;
A = 8'h19; B = 8'h21; #100;
A = 8'h19; B = 8'h22; #100;
A = 8'h19; B = 8'h23; #100;
A = 8'h19; B = 8'h24; #100;
A = 8'h19; B = 8'h25; #100;
A = 8'h19; B = 8'h26; #100;
A = 8'h19; B = 8'h27; #100;
A = 8'h19; B = 8'h28; #100;
A = 8'h19; B = 8'h29; #100;
A = 8'h19; B = 8'h2A; #100;
A = 8'h19; B = 8'h2B; #100;
A = 8'h19; B = 8'h2C; #100;
A = 8'h19; B = 8'h2D; #100;
A = 8'h19; B = 8'h2E; #100;
A = 8'h19; B = 8'h2F; #100;
A = 8'h19; B = 8'h30; #100;
A = 8'h19; B = 8'h31; #100;
A = 8'h19; B = 8'h32; #100;
A = 8'h19; B = 8'h33; #100;
A = 8'h19; B = 8'h34; #100;
A = 8'h19; B = 8'h35; #100;
A = 8'h19; B = 8'h36; #100;
A = 8'h19; B = 8'h37; #100;
A = 8'h19; B = 8'h38; #100;
A = 8'h19; B = 8'h39; #100;
A = 8'h19; B = 8'h3A; #100;
A = 8'h19; B = 8'h3B; #100;
A = 8'h19; B = 8'h3C; #100;
A = 8'h19; B = 8'h3D; #100;
A = 8'h19; B = 8'h3E; #100;
A = 8'h19; B = 8'h3F; #100;
A = 8'h19; B = 8'h40; #100;
A = 8'h19; B = 8'h41; #100;
A = 8'h19; B = 8'h42; #100;
A = 8'h19; B = 8'h43; #100;
A = 8'h19; B = 8'h44; #100;
A = 8'h19; B = 8'h45; #100;
A = 8'h19; B = 8'h46; #100;
A = 8'h19; B = 8'h47; #100;
A = 8'h19; B = 8'h48; #100;
A = 8'h19; B = 8'h49; #100;
A = 8'h19; B = 8'h4A; #100;
A = 8'h19; B = 8'h4B; #100;
A = 8'h19; B = 8'h4C; #100;
A = 8'h19; B = 8'h4D; #100;
A = 8'h19; B = 8'h4E; #100;
A = 8'h19; B = 8'h4F; #100;
A = 8'h19; B = 8'h50; #100;
A = 8'h19; B = 8'h51; #100;
A = 8'h19; B = 8'h52; #100;
A = 8'h19; B = 8'h53; #100;
A = 8'h19; B = 8'h54; #100;
A = 8'h19; B = 8'h55; #100;
A = 8'h19; B = 8'h56; #100;
A = 8'h19; B = 8'h57; #100;
A = 8'h19; B = 8'h58; #100;
A = 8'h19; B = 8'h59; #100;
A = 8'h19; B = 8'h5A; #100;
A = 8'h19; B = 8'h5B; #100;
A = 8'h19; B = 8'h5C; #100;
A = 8'h19; B = 8'h5D; #100;
A = 8'h19; B = 8'h5E; #100;
A = 8'h19; B = 8'h5F; #100;
A = 8'h19; B = 8'h60; #100;
A = 8'h19; B = 8'h61; #100;
A = 8'h19; B = 8'h62; #100;
A = 8'h19; B = 8'h63; #100;
A = 8'h19; B = 8'h64; #100;
A = 8'h19; B = 8'h65; #100;
A = 8'h19; B = 8'h66; #100;
A = 8'h19; B = 8'h67; #100;
A = 8'h19; B = 8'h68; #100;
A = 8'h19; B = 8'h69; #100;
A = 8'h19; B = 8'h6A; #100;
A = 8'h19; B = 8'h6B; #100;
A = 8'h19; B = 8'h6C; #100;
A = 8'h19; B = 8'h6D; #100;
A = 8'h19; B = 8'h6E; #100;
A = 8'h19; B = 8'h6F; #100;
A = 8'h19; B = 8'h70; #100;
A = 8'h19; B = 8'h71; #100;
A = 8'h19; B = 8'h72; #100;
A = 8'h19; B = 8'h73; #100;
A = 8'h19; B = 8'h74; #100;
A = 8'h19; B = 8'h75; #100;
A = 8'h19; B = 8'h76; #100;
A = 8'h19; B = 8'h77; #100;
A = 8'h19; B = 8'h78; #100;
A = 8'h19; B = 8'h79; #100;
A = 8'h19; B = 8'h7A; #100;
A = 8'h19; B = 8'h7B; #100;
A = 8'h19; B = 8'h7C; #100;
A = 8'h19; B = 8'h7D; #100;
A = 8'h19; B = 8'h7E; #100;
A = 8'h19; B = 8'h7F; #100;
A = 8'h19; B = 8'h80; #100;
A = 8'h19; B = 8'h81; #100;
A = 8'h19; B = 8'h82; #100;
A = 8'h19; B = 8'h83; #100;
A = 8'h19; B = 8'h84; #100;
A = 8'h19; B = 8'h85; #100;
A = 8'h19; B = 8'h86; #100;
A = 8'h19; B = 8'h87; #100;
A = 8'h19; B = 8'h88; #100;
A = 8'h19; B = 8'h89; #100;
A = 8'h19; B = 8'h8A; #100;
A = 8'h19; B = 8'h8B; #100;
A = 8'h19; B = 8'h8C; #100;
A = 8'h19; B = 8'h8D; #100;
A = 8'h19; B = 8'h8E; #100;
A = 8'h19; B = 8'h8F; #100;
A = 8'h19; B = 8'h90; #100;
A = 8'h19; B = 8'h91; #100;
A = 8'h19; B = 8'h92; #100;
A = 8'h19; B = 8'h93; #100;
A = 8'h19; B = 8'h94; #100;
A = 8'h19; B = 8'h95; #100;
A = 8'h19; B = 8'h96; #100;
A = 8'h19; B = 8'h97; #100;
A = 8'h19; B = 8'h98; #100;
A = 8'h19; B = 8'h99; #100;
A = 8'h19; B = 8'h9A; #100;
A = 8'h19; B = 8'h9B; #100;
A = 8'h19; B = 8'h9C; #100;
A = 8'h19; B = 8'h9D; #100;
A = 8'h19; B = 8'h9E; #100;
A = 8'h19; B = 8'h9F; #100;
A = 8'h19; B = 8'hA0; #100;
A = 8'h19; B = 8'hA1; #100;
A = 8'h19; B = 8'hA2; #100;
A = 8'h19; B = 8'hA3; #100;
A = 8'h19; B = 8'hA4; #100;
A = 8'h19; B = 8'hA5; #100;
A = 8'h19; B = 8'hA6; #100;
A = 8'h19; B = 8'hA7; #100;
A = 8'h19; B = 8'hA8; #100;
A = 8'h19; B = 8'hA9; #100;
A = 8'h19; B = 8'hAA; #100;
A = 8'h19; B = 8'hAB; #100;
A = 8'h19; B = 8'hAC; #100;
A = 8'h19; B = 8'hAD; #100;
A = 8'h19; B = 8'hAE; #100;
A = 8'h19; B = 8'hAF; #100;
A = 8'h19; B = 8'hB0; #100;
A = 8'h19; B = 8'hB1; #100;
A = 8'h19; B = 8'hB2; #100;
A = 8'h19; B = 8'hB3; #100;
A = 8'h19; B = 8'hB4; #100;
A = 8'h19; B = 8'hB5; #100;
A = 8'h19; B = 8'hB6; #100;
A = 8'h19; B = 8'hB7; #100;
A = 8'h19; B = 8'hB8; #100;
A = 8'h19; B = 8'hB9; #100;
A = 8'h19; B = 8'hBA; #100;
A = 8'h19; B = 8'hBB; #100;
A = 8'h19; B = 8'hBC; #100;
A = 8'h19; B = 8'hBD; #100;
A = 8'h19; B = 8'hBE; #100;
A = 8'h19; B = 8'hBF; #100;
A = 8'h19; B = 8'hC0; #100;
A = 8'h19; B = 8'hC1; #100;
A = 8'h19; B = 8'hC2; #100;
A = 8'h19; B = 8'hC3; #100;
A = 8'h19; B = 8'hC4; #100;
A = 8'h19; B = 8'hC5; #100;
A = 8'h19; B = 8'hC6; #100;
A = 8'h19; B = 8'hC7; #100;
A = 8'h19; B = 8'hC8; #100;
A = 8'h19; B = 8'hC9; #100;
A = 8'h19; B = 8'hCA; #100;
A = 8'h19; B = 8'hCB; #100;
A = 8'h19; B = 8'hCC; #100;
A = 8'h19; B = 8'hCD; #100;
A = 8'h19; B = 8'hCE; #100;
A = 8'h19; B = 8'hCF; #100;
A = 8'h19; B = 8'hD0; #100;
A = 8'h19; B = 8'hD1; #100;
A = 8'h19; B = 8'hD2; #100;
A = 8'h19; B = 8'hD3; #100;
A = 8'h19; B = 8'hD4; #100;
A = 8'h19; B = 8'hD5; #100;
A = 8'h19; B = 8'hD6; #100;
A = 8'h19; B = 8'hD7; #100;
A = 8'h19; B = 8'hD8; #100;
A = 8'h19; B = 8'hD9; #100;
A = 8'h19; B = 8'hDA; #100;
A = 8'h19; B = 8'hDB; #100;
A = 8'h19; B = 8'hDC; #100;
A = 8'h19; B = 8'hDD; #100;
A = 8'h19; B = 8'hDE; #100;
A = 8'h19; B = 8'hDF; #100;
A = 8'h19; B = 8'hE0; #100;
A = 8'h19; B = 8'hE1; #100;
A = 8'h19; B = 8'hE2; #100;
A = 8'h19; B = 8'hE3; #100;
A = 8'h19; B = 8'hE4; #100;
A = 8'h19; B = 8'hE5; #100;
A = 8'h19; B = 8'hE6; #100;
A = 8'h19; B = 8'hE7; #100;
A = 8'h19; B = 8'hE8; #100;
A = 8'h19; B = 8'hE9; #100;
A = 8'h19; B = 8'hEA; #100;
A = 8'h19; B = 8'hEB; #100;
A = 8'h19; B = 8'hEC; #100;
A = 8'h19; B = 8'hED; #100;
A = 8'h19; B = 8'hEE; #100;
A = 8'h19; B = 8'hEF; #100;
A = 8'h19; B = 8'hF0; #100;
A = 8'h19; B = 8'hF1; #100;
A = 8'h19; B = 8'hF2; #100;
A = 8'h19; B = 8'hF3; #100;
A = 8'h19; B = 8'hF4; #100;
A = 8'h19; B = 8'hF5; #100;
A = 8'h19; B = 8'hF6; #100;
A = 8'h19; B = 8'hF7; #100;
A = 8'h19; B = 8'hF8; #100;
A = 8'h19; B = 8'hF9; #100;
A = 8'h19; B = 8'hFA; #100;
A = 8'h19; B = 8'hFB; #100;
A = 8'h19; B = 8'hFC; #100;
A = 8'h19; B = 8'hFD; #100;
A = 8'h19; B = 8'hFE; #100;
A = 8'h19; B = 8'hFF; #100;
A = 8'h1A; B = 8'h0; #100;
A = 8'h1A; B = 8'h1; #100;
A = 8'h1A; B = 8'h2; #100;
A = 8'h1A; B = 8'h3; #100;
A = 8'h1A; B = 8'h4; #100;
A = 8'h1A; B = 8'h5; #100;
A = 8'h1A; B = 8'h6; #100;
A = 8'h1A; B = 8'h7; #100;
A = 8'h1A; B = 8'h8; #100;
A = 8'h1A; B = 8'h9; #100;
A = 8'h1A; B = 8'hA; #100;
A = 8'h1A; B = 8'hB; #100;
A = 8'h1A; B = 8'hC; #100;
A = 8'h1A; B = 8'hD; #100;
A = 8'h1A; B = 8'hE; #100;
A = 8'h1A; B = 8'hF; #100;
A = 8'h1A; B = 8'h10; #100;
A = 8'h1A; B = 8'h11; #100;
A = 8'h1A; B = 8'h12; #100;
A = 8'h1A; B = 8'h13; #100;
A = 8'h1A; B = 8'h14; #100;
A = 8'h1A; B = 8'h15; #100;
A = 8'h1A; B = 8'h16; #100;
A = 8'h1A; B = 8'h17; #100;
A = 8'h1A; B = 8'h18; #100;
A = 8'h1A; B = 8'h19; #100;
A = 8'h1A; B = 8'h1A; #100;
A = 8'h1A; B = 8'h1B; #100;
A = 8'h1A; B = 8'h1C; #100;
A = 8'h1A; B = 8'h1D; #100;
A = 8'h1A; B = 8'h1E; #100;
A = 8'h1A; B = 8'h1F; #100;
A = 8'h1A; B = 8'h20; #100;
A = 8'h1A; B = 8'h21; #100;
A = 8'h1A; B = 8'h22; #100;
A = 8'h1A; B = 8'h23; #100;
A = 8'h1A; B = 8'h24; #100;
A = 8'h1A; B = 8'h25; #100;
A = 8'h1A; B = 8'h26; #100;
A = 8'h1A; B = 8'h27; #100;
A = 8'h1A; B = 8'h28; #100;
A = 8'h1A; B = 8'h29; #100;
A = 8'h1A; B = 8'h2A; #100;
A = 8'h1A; B = 8'h2B; #100;
A = 8'h1A; B = 8'h2C; #100;
A = 8'h1A; B = 8'h2D; #100;
A = 8'h1A; B = 8'h2E; #100;
A = 8'h1A; B = 8'h2F; #100;
A = 8'h1A; B = 8'h30; #100;
A = 8'h1A; B = 8'h31; #100;
A = 8'h1A; B = 8'h32; #100;
A = 8'h1A; B = 8'h33; #100;
A = 8'h1A; B = 8'h34; #100;
A = 8'h1A; B = 8'h35; #100;
A = 8'h1A; B = 8'h36; #100;
A = 8'h1A; B = 8'h37; #100;
A = 8'h1A; B = 8'h38; #100;
A = 8'h1A; B = 8'h39; #100;
A = 8'h1A; B = 8'h3A; #100;
A = 8'h1A; B = 8'h3B; #100;
A = 8'h1A; B = 8'h3C; #100;
A = 8'h1A; B = 8'h3D; #100;
A = 8'h1A; B = 8'h3E; #100;
A = 8'h1A; B = 8'h3F; #100;
A = 8'h1A; B = 8'h40; #100;
A = 8'h1A; B = 8'h41; #100;
A = 8'h1A; B = 8'h42; #100;
A = 8'h1A; B = 8'h43; #100;
A = 8'h1A; B = 8'h44; #100;
A = 8'h1A; B = 8'h45; #100;
A = 8'h1A; B = 8'h46; #100;
A = 8'h1A; B = 8'h47; #100;
A = 8'h1A; B = 8'h48; #100;
A = 8'h1A; B = 8'h49; #100;
A = 8'h1A; B = 8'h4A; #100;
A = 8'h1A; B = 8'h4B; #100;
A = 8'h1A; B = 8'h4C; #100;
A = 8'h1A; B = 8'h4D; #100;
A = 8'h1A; B = 8'h4E; #100;
A = 8'h1A; B = 8'h4F; #100;
A = 8'h1A; B = 8'h50; #100;
A = 8'h1A; B = 8'h51; #100;
A = 8'h1A; B = 8'h52; #100;
A = 8'h1A; B = 8'h53; #100;
A = 8'h1A; B = 8'h54; #100;
A = 8'h1A; B = 8'h55; #100;
A = 8'h1A; B = 8'h56; #100;
A = 8'h1A; B = 8'h57; #100;
A = 8'h1A; B = 8'h58; #100;
A = 8'h1A; B = 8'h59; #100;
A = 8'h1A; B = 8'h5A; #100;
A = 8'h1A; B = 8'h5B; #100;
A = 8'h1A; B = 8'h5C; #100;
A = 8'h1A; B = 8'h5D; #100;
A = 8'h1A; B = 8'h5E; #100;
A = 8'h1A; B = 8'h5F; #100;
A = 8'h1A; B = 8'h60; #100;
A = 8'h1A; B = 8'h61; #100;
A = 8'h1A; B = 8'h62; #100;
A = 8'h1A; B = 8'h63; #100;
A = 8'h1A; B = 8'h64; #100;
A = 8'h1A; B = 8'h65; #100;
A = 8'h1A; B = 8'h66; #100;
A = 8'h1A; B = 8'h67; #100;
A = 8'h1A; B = 8'h68; #100;
A = 8'h1A; B = 8'h69; #100;
A = 8'h1A; B = 8'h6A; #100;
A = 8'h1A; B = 8'h6B; #100;
A = 8'h1A; B = 8'h6C; #100;
A = 8'h1A; B = 8'h6D; #100;
A = 8'h1A; B = 8'h6E; #100;
A = 8'h1A; B = 8'h6F; #100;
A = 8'h1A; B = 8'h70; #100;
A = 8'h1A; B = 8'h71; #100;
A = 8'h1A; B = 8'h72; #100;
A = 8'h1A; B = 8'h73; #100;
A = 8'h1A; B = 8'h74; #100;
A = 8'h1A; B = 8'h75; #100;
A = 8'h1A; B = 8'h76; #100;
A = 8'h1A; B = 8'h77; #100;
A = 8'h1A; B = 8'h78; #100;
A = 8'h1A; B = 8'h79; #100;
A = 8'h1A; B = 8'h7A; #100;
A = 8'h1A; B = 8'h7B; #100;
A = 8'h1A; B = 8'h7C; #100;
A = 8'h1A; B = 8'h7D; #100;
A = 8'h1A; B = 8'h7E; #100;
A = 8'h1A; B = 8'h7F; #100;
A = 8'h1A; B = 8'h80; #100;
A = 8'h1A; B = 8'h81; #100;
A = 8'h1A; B = 8'h82; #100;
A = 8'h1A; B = 8'h83; #100;
A = 8'h1A; B = 8'h84; #100;
A = 8'h1A; B = 8'h85; #100;
A = 8'h1A; B = 8'h86; #100;
A = 8'h1A; B = 8'h87; #100;
A = 8'h1A; B = 8'h88; #100;
A = 8'h1A; B = 8'h89; #100;
A = 8'h1A; B = 8'h8A; #100;
A = 8'h1A; B = 8'h8B; #100;
A = 8'h1A; B = 8'h8C; #100;
A = 8'h1A; B = 8'h8D; #100;
A = 8'h1A; B = 8'h8E; #100;
A = 8'h1A; B = 8'h8F; #100;
A = 8'h1A; B = 8'h90; #100;
A = 8'h1A; B = 8'h91; #100;
A = 8'h1A; B = 8'h92; #100;
A = 8'h1A; B = 8'h93; #100;
A = 8'h1A; B = 8'h94; #100;
A = 8'h1A; B = 8'h95; #100;
A = 8'h1A; B = 8'h96; #100;
A = 8'h1A; B = 8'h97; #100;
A = 8'h1A; B = 8'h98; #100;
A = 8'h1A; B = 8'h99; #100;
A = 8'h1A; B = 8'h9A; #100;
A = 8'h1A; B = 8'h9B; #100;
A = 8'h1A; B = 8'h9C; #100;
A = 8'h1A; B = 8'h9D; #100;
A = 8'h1A; B = 8'h9E; #100;
A = 8'h1A; B = 8'h9F; #100;
A = 8'h1A; B = 8'hA0; #100;
A = 8'h1A; B = 8'hA1; #100;
A = 8'h1A; B = 8'hA2; #100;
A = 8'h1A; B = 8'hA3; #100;
A = 8'h1A; B = 8'hA4; #100;
A = 8'h1A; B = 8'hA5; #100;
A = 8'h1A; B = 8'hA6; #100;
A = 8'h1A; B = 8'hA7; #100;
A = 8'h1A; B = 8'hA8; #100;
A = 8'h1A; B = 8'hA9; #100;
A = 8'h1A; B = 8'hAA; #100;
A = 8'h1A; B = 8'hAB; #100;
A = 8'h1A; B = 8'hAC; #100;
A = 8'h1A; B = 8'hAD; #100;
A = 8'h1A; B = 8'hAE; #100;
A = 8'h1A; B = 8'hAF; #100;
A = 8'h1A; B = 8'hB0; #100;
A = 8'h1A; B = 8'hB1; #100;
A = 8'h1A; B = 8'hB2; #100;
A = 8'h1A; B = 8'hB3; #100;
A = 8'h1A; B = 8'hB4; #100;
A = 8'h1A; B = 8'hB5; #100;
A = 8'h1A; B = 8'hB6; #100;
A = 8'h1A; B = 8'hB7; #100;
A = 8'h1A; B = 8'hB8; #100;
A = 8'h1A; B = 8'hB9; #100;
A = 8'h1A; B = 8'hBA; #100;
A = 8'h1A; B = 8'hBB; #100;
A = 8'h1A; B = 8'hBC; #100;
A = 8'h1A; B = 8'hBD; #100;
A = 8'h1A; B = 8'hBE; #100;
A = 8'h1A; B = 8'hBF; #100;
A = 8'h1A; B = 8'hC0; #100;
A = 8'h1A; B = 8'hC1; #100;
A = 8'h1A; B = 8'hC2; #100;
A = 8'h1A; B = 8'hC3; #100;
A = 8'h1A; B = 8'hC4; #100;
A = 8'h1A; B = 8'hC5; #100;
A = 8'h1A; B = 8'hC6; #100;
A = 8'h1A; B = 8'hC7; #100;
A = 8'h1A; B = 8'hC8; #100;
A = 8'h1A; B = 8'hC9; #100;
A = 8'h1A; B = 8'hCA; #100;
A = 8'h1A; B = 8'hCB; #100;
A = 8'h1A; B = 8'hCC; #100;
A = 8'h1A; B = 8'hCD; #100;
A = 8'h1A; B = 8'hCE; #100;
A = 8'h1A; B = 8'hCF; #100;
A = 8'h1A; B = 8'hD0; #100;
A = 8'h1A; B = 8'hD1; #100;
A = 8'h1A; B = 8'hD2; #100;
A = 8'h1A; B = 8'hD3; #100;
A = 8'h1A; B = 8'hD4; #100;
A = 8'h1A; B = 8'hD5; #100;
A = 8'h1A; B = 8'hD6; #100;
A = 8'h1A; B = 8'hD7; #100;
A = 8'h1A; B = 8'hD8; #100;
A = 8'h1A; B = 8'hD9; #100;
A = 8'h1A; B = 8'hDA; #100;
A = 8'h1A; B = 8'hDB; #100;
A = 8'h1A; B = 8'hDC; #100;
A = 8'h1A; B = 8'hDD; #100;
A = 8'h1A; B = 8'hDE; #100;
A = 8'h1A; B = 8'hDF; #100;
A = 8'h1A; B = 8'hE0; #100;
A = 8'h1A; B = 8'hE1; #100;
A = 8'h1A; B = 8'hE2; #100;
A = 8'h1A; B = 8'hE3; #100;
A = 8'h1A; B = 8'hE4; #100;
A = 8'h1A; B = 8'hE5; #100;
A = 8'h1A; B = 8'hE6; #100;
A = 8'h1A; B = 8'hE7; #100;
A = 8'h1A; B = 8'hE8; #100;
A = 8'h1A; B = 8'hE9; #100;
A = 8'h1A; B = 8'hEA; #100;
A = 8'h1A; B = 8'hEB; #100;
A = 8'h1A; B = 8'hEC; #100;
A = 8'h1A; B = 8'hED; #100;
A = 8'h1A; B = 8'hEE; #100;
A = 8'h1A; B = 8'hEF; #100;
A = 8'h1A; B = 8'hF0; #100;
A = 8'h1A; B = 8'hF1; #100;
A = 8'h1A; B = 8'hF2; #100;
A = 8'h1A; B = 8'hF3; #100;
A = 8'h1A; B = 8'hF4; #100;
A = 8'h1A; B = 8'hF5; #100;
A = 8'h1A; B = 8'hF6; #100;
A = 8'h1A; B = 8'hF7; #100;
A = 8'h1A; B = 8'hF8; #100;
A = 8'h1A; B = 8'hF9; #100;
A = 8'h1A; B = 8'hFA; #100;
A = 8'h1A; B = 8'hFB; #100;
A = 8'h1A; B = 8'hFC; #100;
A = 8'h1A; B = 8'hFD; #100;
A = 8'h1A; B = 8'hFE; #100;
A = 8'h1A; B = 8'hFF; #100;
A = 8'h1B; B = 8'h0; #100;
A = 8'h1B; B = 8'h1; #100;
A = 8'h1B; B = 8'h2; #100;
A = 8'h1B; B = 8'h3; #100;
A = 8'h1B; B = 8'h4; #100;
A = 8'h1B; B = 8'h5; #100;
A = 8'h1B; B = 8'h6; #100;
A = 8'h1B; B = 8'h7; #100;
A = 8'h1B; B = 8'h8; #100;
A = 8'h1B; B = 8'h9; #100;
A = 8'h1B; B = 8'hA; #100;
A = 8'h1B; B = 8'hB; #100;
A = 8'h1B; B = 8'hC; #100;
A = 8'h1B; B = 8'hD; #100;
A = 8'h1B; B = 8'hE; #100;
A = 8'h1B; B = 8'hF; #100;
A = 8'h1B; B = 8'h10; #100;
A = 8'h1B; B = 8'h11; #100;
A = 8'h1B; B = 8'h12; #100;
A = 8'h1B; B = 8'h13; #100;
A = 8'h1B; B = 8'h14; #100;
A = 8'h1B; B = 8'h15; #100;
A = 8'h1B; B = 8'h16; #100;
A = 8'h1B; B = 8'h17; #100;
A = 8'h1B; B = 8'h18; #100;
A = 8'h1B; B = 8'h19; #100;
A = 8'h1B; B = 8'h1A; #100;
A = 8'h1B; B = 8'h1B; #100;
A = 8'h1B; B = 8'h1C; #100;
A = 8'h1B; B = 8'h1D; #100;
A = 8'h1B; B = 8'h1E; #100;
A = 8'h1B; B = 8'h1F; #100;
A = 8'h1B; B = 8'h20; #100;
A = 8'h1B; B = 8'h21; #100;
A = 8'h1B; B = 8'h22; #100;
A = 8'h1B; B = 8'h23; #100;
A = 8'h1B; B = 8'h24; #100;
A = 8'h1B; B = 8'h25; #100;
A = 8'h1B; B = 8'h26; #100;
A = 8'h1B; B = 8'h27; #100;
A = 8'h1B; B = 8'h28; #100;
A = 8'h1B; B = 8'h29; #100;
A = 8'h1B; B = 8'h2A; #100;
A = 8'h1B; B = 8'h2B; #100;
A = 8'h1B; B = 8'h2C; #100;
A = 8'h1B; B = 8'h2D; #100;
A = 8'h1B; B = 8'h2E; #100;
A = 8'h1B; B = 8'h2F; #100;
A = 8'h1B; B = 8'h30; #100;
A = 8'h1B; B = 8'h31; #100;
A = 8'h1B; B = 8'h32; #100;
A = 8'h1B; B = 8'h33; #100;
A = 8'h1B; B = 8'h34; #100;
A = 8'h1B; B = 8'h35; #100;
A = 8'h1B; B = 8'h36; #100;
A = 8'h1B; B = 8'h37; #100;
A = 8'h1B; B = 8'h38; #100;
A = 8'h1B; B = 8'h39; #100;
A = 8'h1B; B = 8'h3A; #100;
A = 8'h1B; B = 8'h3B; #100;
A = 8'h1B; B = 8'h3C; #100;
A = 8'h1B; B = 8'h3D; #100;
A = 8'h1B; B = 8'h3E; #100;
A = 8'h1B; B = 8'h3F; #100;
A = 8'h1B; B = 8'h40; #100;
A = 8'h1B; B = 8'h41; #100;
A = 8'h1B; B = 8'h42; #100;
A = 8'h1B; B = 8'h43; #100;
A = 8'h1B; B = 8'h44; #100;
A = 8'h1B; B = 8'h45; #100;
A = 8'h1B; B = 8'h46; #100;
A = 8'h1B; B = 8'h47; #100;
A = 8'h1B; B = 8'h48; #100;
A = 8'h1B; B = 8'h49; #100;
A = 8'h1B; B = 8'h4A; #100;
A = 8'h1B; B = 8'h4B; #100;
A = 8'h1B; B = 8'h4C; #100;
A = 8'h1B; B = 8'h4D; #100;
A = 8'h1B; B = 8'h4E; #100;
A = 8'h1B; B = 8'h4F; #100;
A = 8'h1B; B = 8'h50; #100;
A = 8'h1B; B = 8'h51; #100;
A = 8'h1B; B = 8'h52; #100;
A = 8'h1B; B = 8'h53; #100;
A = 8'h1B; B = 8'h54; #100;
A = 8'h1B; B = 8'h55; #100;
A = 8'h1B; B = 8'h56; #100;
A = 8'h1B; B = 8'h57; #100;
A = 8'h1B; B = 8'h58; #100;
A = 8'h1B; B = 8'h59; #100;
A = 8'h1B; B = 8'h5A; #100;
A = 8'h1B; B = 8'h5B; #100;
A = 8'h1B; B = 8'h5C; #100;
A = 8'h1B; B = 8'h5D; #100;
A = 8'h1B; B = 8'h5E; #100;
A = 8'h1B; B = 8'h5F; #100;
A = 8'h1B; B = 8'h60; #100;
A = 8'h1B; B = 8'h61; #100;
A = 8'h1B; B = 8'h62; #100;
A = 8'h1B; B = 8'h63; #100;
A = 8'h1B; B = 8'h64; #100;
A = 8'h1B; B = 8'h65; #100;
A = 8'h1B; B = 8'h66; #100;
A = 8'h1B; B = 8'h67; #100;
A = 8'h1B; B = 8'h68; #100;
A = 8'h1B; B = 8'h69; #100;
A = 8'h1B; B = 8'h6A; #100;
A = 8'h1B; B = 8'h6B; #100;
A = 8'h1B; B = 8'h6C; #100;
A = 8'h1B; B = 8'h6D; #100;
A = 8'h1B; B = 8'h6E; #100;
A = 8'h1B; B = 8'h6F; #100;
A = 8'h1B; B = 8'h70; #100;
A = 8'h1B; B = 8'h71; #100;
A = 8'h1B; B = 8'h72; #100;
A = 8'h1B; B = 8'h73; #100;
A = 8'h1B; B = 8'h74; #100;
A = 8'h1B; B = 8'h75; #100;
A = 8'h1B; B = 8'h76; #100;
A = 8'h1B; B = 8'h77; #100;
A = 8'h1B; B = 8'h78; #100;
A = 8'h1B; B = 8'h79; #100;
A = 8'h1B; B = 8'h7A; #100;
A = 8'h1B; B = 8'h7B; #100;
A = 8'h1B; B = 8'h7C; #100;
A = 8'h1B; B = 8'h7D; #100;
A = 8'h1B; B = 8'h7E; #100;
A = 8'h1B; B = 8'h7F; #100;
A = 8'h1B; B = 8'h80; #100;
A = 8'h1B; B = 8'h81; #100;
A = 8'h1B; B = 8'h82; #100;
A = 8'h1B; B = 8'h83; #100;
A = 8'h1B; B = 8'h84; #100;
A = 8'h1B; B = 8'h85; #100;
A = 8'h1B; B = 8'h86; #100;
A = 8'h1B; B = 8'h87; #100;
A = 8'h1B; B = 8'h88; #100;
A = 8'h1B; B = 8'h89; #100;
A = 8'h1B; B = 8'h8A; #100;
A = 8'h1B; B = 8'h8B; #100;
A = 8'h1B; B = 8'h8C; #100;
A = 8'h1B; B = 8'h8D; #100;
A = 8'h1B; B = 8'h8E; #100;
A = 8'h1B; B = 8'h8F; #100;
A = 8'h1B; B = 8'h90; #100;
A = 8'h1B; B = 8'h91; #100;
A = 8'h1B; B = 8'h92; #100;
A = 8'h1B; B = 8'h93; #100;
A = 8'h1B; B = 8'h94; #100;
A = 8'h1B; B = 8'h95; #100;
A = 8'h1B; B = 8'h96; #100;
A = 8'h1B; B = 8'h97; #100;
A = 8'h1B; B = 8'h98; #100;
A = 8'h1B; B = 8'h99; #100;
A = 8'h1B; B = 8'h9A; #100;
A = 8'h1B; B = 8'h9B; #100;
A = 8'h1B; B = 8'h9C; #100;
A = 8'h1B; B = 8'h9D; #100;
A = 8'h1B; B = 8'h9E; #100;
A = 8'h1B; B = 8'h9F; #100;
A = 8'h1B; B = 8'hA0; #100;
A = 8'h1B; B = 8'hA1; #100;
A = 8'h1B; B = 8'hA2; #100;
A = 8'h1B; B = 8'hA3; #100;
A = 8'h1B; B = 8'hA4; #100;
A = 8'h1B; B = 8'hA5; #100;
A = 8'h1B; B = 8'hA6; #100;
A = 8'h1B; B = 8'hA7; #100;
A = 8'h1B; B = 8'hA8; #100;
A = 8'h1B; B = 8'hA9; #100;
A = 8'h1B; B = 8'hAA; #100;
A = 8'h1B; B = 8'hAB; #100;
A = 8'h1B; B = 8'hAC; #100;
A = 8'h1B; B = 8'hAD; #100;
A = 8'h1B; B = 8'hAE; #100;
A = 8'h1B; B = 8'hAF; #100;
A = 8'h1B; B = 8'hB0; #100;
A = 8'h1B; B = 8'hB1; #100;
A = 8'h1B; B = 8'hB2; #100;
A = 8'h1B; B = 8'hB3; #100;
A = 8'h1B; B = 8'hB4; #100;
A = 8'h1B; B = 8'hB5; #100;
A = 8'h1B; B = 8'hB6; #100;
A = 8'h1B; B = 8'hB7; #100;
A = 8'h1B; B = 8'hB8; #100;
A = 8'h1B; B = 8'hB9; #100;
A = 8'h1B; B = 8'hBA; #100;
A = 8'h1B; B = 8'hBB; #100;
A = 8'h1B; B = 8'hBC; #100;
A = 8'h1B; B = 8'hBD; #100;
A = 8'h1B; B = 8'hBE; #100;
A = 8'h1B; B = 8'hBF; #100;
A = 8'h1B; B = 8'hC0; #100;
A = 8'h1B; B = 8'hC1; #100;
A = 8'h1B; B = 8'hC2; #100;
A = 8'h1B; B = 8'hC3; #100;
A = 8'h1B; B = 8'hC4; #100;
A = 8'h1B; B = 8'hC5; #100;
A = 8'h1B; B = 8'hC6; #100;
A = 8'h1B; B = 8'hC7; #100;
A = 8'h1B; B = 8'hC8; #100;
A = 8'h1B; B = 8'hC9; #100;
A = 8'h1B; B = 8'hCA; #100;
A = 8'h1B; B = 8'hCB; #100;
A = 8'h1B; B = 8'hCC; #100;
A = 8'h1B; B = 8'hCD; #100;
A = 8'h1B; B = 8'hCE; #100;
A = 8'h1B; B = 8'hCF; #100;
A = 8'h1B; B = 8'hD0; #100;
A = 8'h1B; B = 8'hD1; #100;
A = 8'h1B; B = 8'hD2; #100;
A = 8'h1B; B = 8'hD3; #100;
A = 8'h1B; B = 8'hD4; #100;
A = 8'h1B; B = 8'hD5; #100;
A = 8'h1B; B = 8'hD6; #100;
A = 8'h1B; B = 8'hD7; #100;
A = 8'h1B; B = 8'hD8; #100;
A = 8'h1B; B = 8'hD9; #100;
A = 8'h1B; B = 8'hDA; #100;
A = 8'h1B; B = 8'hDB; #100;
A = 8'h1B; B = 8'hDC; #100;
A = 8'h1B; B = 8'hDD; #100;
A = 8'h1B; B = 8'hDE; #100;
A = 8'h1B; B = 8'hDF; #100;
A = 8'h1B; B = 8'hE0; #100;
A = 8'h1B; B = 8'hE1; #100;
A = 8'h1B; B = 8'hE2; #100;
A = 8'h1B; B = 8'hE3; #100;
A = 8'h1B; B = 8'hE4; #100;
A = 8'h1B; B = 8'hE5; #100;
A = 8'h1B; B = 8'hE6; #100;
A = 8'h1B; B = 8'hE7; #100;
A = 8'h1B; B = 8'hE8; #100;
A = 8'h1B; B = 8'hE9; #100;
A = 8'h1B; B = 8'hEA; #100;
A = 8'h1B; B = 8'hEB; #100;
A = 8'h1B; B = 8'hEC; #100;
A = 8'h1B; B = 8'hED; #100;
A = 8'h1B; B = 8'hEE; #100;
A = 8'h1B; B = 8'hEF; #100;
A = 8'h1B; B = 8'hF0; #100;
A = 8'h1B; B = 8'hF1; #100;
A = 8'h1B; B = 8'hF2; #100;
A = 8'h1B; B = 8'hF3; #100;
A = 8'h1B; B = 8'hF4; #100;
A = 8'h1B; B = 8'hF5; #100;
A = 8'h1B; B = 8'hF6; #100;
A = 8'h1B; B = 8'hF7; #100;
A = 8'h1B; B = 8'hF8; #100;
A = 8'h1B; B = 8'hF9; #100;
A = 8'h1B; B = 8'hFA; #100;
A = 8'h1B; B = 8'hFB; #100;
A = 8'h1B; B = 8'hFC; #100;
A = 8'h1B; B = 8'hFD; #100;
A = 8'h1B; B = 8'hFE; #100;
A = 8'h1B; B = 8'hFF; #100;
A = 8'h1C; B = 8'h0; #100;
A = 8'h1C; B = 8'h1; #100;
A = 8'h1C; B = 8'h2; #100;
A = 8'h1C; B = 8'h3; #100;
A = 8'h1C; B = 8'h4; #100;
A = 8'h1C; B = 8'h5; #100;
A = 8'h1C; B = 8'h6; #100;
A = 8'h1C; B = 8'h7; #100;
A = 8'h1C; B = 8'h8; #100;
A = 8'h1C; B = 8'h9; #100;
A = 8'h1C; B = 8'hA; #100;
A = 8'h1C; B = 8'hB; #100;
A = 8'h1C; B = 8'hC; #100;
A = 8'h1C; B = 8'hD; #100;
A = 8'h1C; B = 8'hE; #100;
A = 8'h1C; B = 8'hF; #100;
A = 8'h1C; B = 8'h10; #100;
A = 8'h1C; B = 8'h11; #100;
A = 8'h1C; B = 8'h12; #100;
A = 8'h1C; B = 8'h13; #100;
A = 8'h1C; B = 8'h14; #100;
A = 8'h1C; B = 8'h15; #100;
A = 8'h1C; B = 8'h16; #100;
A = 8'h1C; B = 8'h17; #100;
A = 8'h1C; B = 8'h18; #100;
A = 8'h1C; B = 8'h19; #100;
A = 8'h1C; B = 8'h1A; #100;
A = 8'h1C; B = 8'h1B; #100;
A = 8'h1C; B = 8'h1C; #100;
A = 8'h1C; B = 8'h1D; #100;
A = 8'h1C; B = 8'h1E; #100;
A = 8'h1C; B = 8'h1F; #100;
A = 8'h1C; B = 8'h20; #100;
A = 8'h1C; B = 8'h21; #100;
A = 8'h1C; B = 8'h22; #100;
A = 8'h1C; B = 8'h23; #100;
A = 8'h1C; B = 8'h24; #100;
A = 8'h1C; B = 8'h25; #100;
A = 8'h1C; B = 8'h26; #100;
A = 8'h1C; B = 8'h27; #100;
A = 8'h1C; B = 8'h28; #100;
A = 8'h1C; B = 8'h29; #100;
A = 8'h1C; B = 8'h2A; #100;
A = 8'h1C; B = 8'h2B; #100;
A = 8'h1C; B = 8'h2C; #100;
A = 8'h1C; B = 8'h2D; #100;
A = 8'h1C; B = 8'h2E; #100;
A = 8'h1C; B = 8'h2F; #100;
A = 8'h1C; B = 8'h30; #100;
A = 8'h1C; B = 8'h31; #100;
A = 8'h1C; B = 8'h32; #100;
A = 8'h1C; B = 8'h33; #100;
A = 8'h1C; B = 8'h34; #100;
A = 8'h1C; B = 8'h35; #100;
A = 8'h1C; B = 8'h36; #100;
A = 8'h1C; B = 8'h37; #100;
A = 8'h1C; B = 8'h38; #100;
A = 8'h1C; B = 8'h39; #100;
A = 8'h1C; B = 8'h3A; #100;
A = 8'h1C; B = 8'h3B; #100;
A = 8'h1C; B = 8'h3C; #100;
A = 8'h1C; B = 8'h3D; #100;
A = 8'h1C; B = 8'h3E; #100;
A = 8'h1C; B = 8'h3F; #100;
A = 8'h1C; B = 8'h40; #100;
A = 8'h1C; B = 8'h41; #100;
A = 8'h1C; B = 8'h42; #100;
A = 8'h1C; B = 8'h43; #100;
A = 8'h1C; B = 8'h44; #100;
A = 8'h1C; B = 8'h45; #100;
A = 8'h1C; B = 8'h46; #100;
A = 8'h1C; B = 8'h47; #100;
A = 8'h1C; B = 8'h48; #100;
A = 8'h1C; B = 8'h49; #100;
A = 8'h1C; B = 8'h4A; #100;
A = 8'h1C; B = 8'h4B; #100;
A = 8'h1C; B = 8'h4C; #100;
A = 8'h1C; B = 8'h4D; #100;
A = 8'h1C; B = 8'h4E; #100;
A = 8'h1C; B = 8'h4F; #100;
A = 8'h1C; B = 8'h50; #100;
A = 8'h1C; B = 8'h51; #100;
A = 8'h1C; B = 8'h52; #100;
A = 8'h1C; B = 8'h53; #100;
A = 8'h1C; B = 8'h54; #100;
A = 8'h1C; B = 8'h55; #100;
A = 8'h1C; B = 8'h56; #100;
A = 8'h1C; B = 8'h57; #100;
A = 8'h1C; B = 8'h58; #100;
A = 8'h1C; B = 8'h59; #100;
A = 8'h1C; B = 8'h5A; #100;
A = 8'h1C; B = 8'h5B; #100;
A = 8'h1C; B = 8'h5C; #100;
A = 8'h1C; B = 8'h5D; #100;
A = 8'h1C; B = 8'h5E; #100;
A = 8'h1C; B = 8'h5F; #100;
A = 8'h1C; B = 8'h60; #100;
A = 8'h1C; B = 8'h61; #100;
A = 8'h1C; B = 8'h62; #100;
A = 8'h1C; B = 8'h63; #100;
A = 8'h1C; B = 8'h64; #100;
A = 8'h1C; B = 8'h65; #100;
A = 8'h1C; B = 8'h66; #100;
A = 8'h1C; B = 8'h67; #100;
A = 8'h1C; B = 8'h68; #100;
A = 8'h1C; B = 8'h69; #100;
A = 8'h1C; B = 8'h6A; #100;
A = 8'h1C; B = 8'h6B; #100;
A = 8'h1C; B = 8'h6C; #100;
A = 8'h1C; B = 8'h6D; #100;
A = 8'h1C; B = 8'h6E; #100;
A = 8'h1C; B = 8'h6F; #100;
A = 8'h1C; B = 8'h70; #100;
A = 8'h1C; B = 8'h71; #100;
A = 8'h1C; B = 8'h72; #100;
A = 8'h1C; B = 8'h73; #100;
A = 8'h1C; B = 8'h74; #100;
A = 8'h1C; B = 8'h75; #100;
A = 8'h1C; B = 8'h76; #100;
A = 8'h1C; B = 8'h77; #100;
A = 8'h1C; B = 8'h78; #100;
A = 8'h1C; B = 8'h79; #100;
A = 8'h1C; B = 8'h7A; #100;
A = 8'h1C; B = 8'h7B; #100;
A = 8'h1C; B = 8'h7C; #100;
A = 8'h1C; B = 8'h7D; #100;
A = 8'h1C; B = 8'h7E; #100;
A = 8'h1C; B = 8'h7F; #100;
A = 8'h1C; B = 8'h80; #100;
A = 8'h1C; B = 8'h81; #100;
A = 8'h1C; B = 8'h82; #100;
A = 8'h1C; B = 8'h83; #100;
A = 8'h1C; B = 8'h84; #100;
A = 8'h1C; B = 8'h85; #100;
A = 8'h1C; B = 8'h86; #100;
A = 8'h1C; B = 8'h87; #100;
A = 8'h1C; B = 8'h88; #100;
A = 8'h1C; B = 8'h89; #100;
A = 8'h1C; B = 8'h8A; #100;
A = 8'h1C; B = 8'h8B; #100;
A = 8'h1C; B = 8'h8C; #100;
A = 8'h1C; B = 8'h8D; #100;
A = 8'h1C; B = 8'h8E; #100;
A = 8'h1C; B = 8'h8F; #100;
A = 8'h1C; B = 8'h90; #100;
A = 8'h1C; B = 8'h91; #100;
A = 8'h1C; B = 8'h92; #100;
A = 8'h1C; B = 8'h93; #100;
A = 8'h1C; B = 8'h94; #100;
A = 8'h1C; B = 8'h95; #100;
A = 8'h1C; B = 8'h96; #100;
A = 8'h1C; B = 8'h97; #100;
A = 8'h1C; B = 8'h98; #100;
A = 8'h1C; B = 8'h99; #100;
A = 8'h1C; B = 8'h9A; #100;
A = 8'h1C; B = 8'h9B; #100;
A = 8'h1C; B = 8'h9C; #100;
A = 8'h1C; B = 8'h9D; #100;
A = 8'h1C; B = 8'h9E; #100;
A = 8'h1C; B = 8'h9F; #100;
A = 8'h1C; B = 8'hA0; #100;
A = 8'h1C; B = 8'hA1; #100;
A = 8'h1C; B = 8'hA2; #100;
A = 8'h1C; B = 8'hA3; #100;
A = 8'h1C; B = 8'hA4; #100;
A = 8'h1C; B = 8'hA5; #100;
A = 8'h1C; B = 8'hA6; #100;
A = 8'h1C; B = 8'hA7; #100;
A = 8'h1C; B = 8'hA8; #100;
A = 8'h1C; B = 8'hA9; #100;
A = 8'h1C; B = 8'hAA; #100;
A = 8'h1C; B = 8'hAB; #100;
A = 8'h1C; B = 8'hAC; #100;
A = 8'h1C; B = 8'hAD; #100;
A = 8'h1C; B = 8'hAE; #100;
A = 8'h1C; B = 8'hAF; #100;
A = 8'h1C; B = 8'hB0; #100;
A = 8'h1C; B = 8'hB1; #100;
A = 8'h1C; B = 8'hB2; #100;
A = 8'h1C; B = 8'hB3; #100;
A = 8'h1C; B = 8'hB4; #100;
A = 8'h1C; B = 8'hB5; #100;
A = 8'h1C; B = 8'hB6; #100;
A = 8'h1C; B = 8'hB7; #100;
A = 8'h1C; B = 8'hB8; #100;
A = 8'h1C; B = 8'hB9; #100;
A = 8'h1C; B = 8'hBA; #100;
A = 8'h1C; B = 8'hBB; #100;
A = 8'h1C; B = 8'hBC; #100;
A = 8'h1C; B = 8'hBD; #100;
A = 8'h1C; B = 8'hBE; #100;
A = 8'h1C; B = 8'hBF; #100;
A = 8'h1C; B = 8'hC0; #100;
A = 8'h1C; B = 8'hC1; #100;
A = 8'h1C; B = 8'hC2; #100;
A = 8'h1C; B = 8'hC3; #100;
A = 8'h1C; B = 8'hC4; #100;
A = 8'h1C; B = 8'hC5; #100;
A = 8'h1C; B = 8'hC6; #100;
A = 8'h1C; B = 8'hC7; #100;
A = 8'h1C; B = 8'hC8; #100;
A = 8'h1C; B = 8'hC9; #100;
A = 8'h1C; B = 8'hCA; #100;
A = 8'h1C; B = 8'hCB; #100;
A = 8'h1C; B = 8'hCC; #100;
A = 8'h1C; B = 8'hCD; #100;
A = 8'h1C; B = 8'hCE; #100;
A = 8'h1C; B = 8'hCF; #100;
A = 8'h1C; B = 8'hD0; #100;
A = 8'h1C; B = 8'hD1; #100;
A = 8'h1C; B = 8'hD2; #100;
A = 8'h1C; B = 8'hD3; #100;
A = 8'h1C; B = 8'hD4; #100;
A = 8'h1C; B = 8'hD5; #100;
A = 8'h1C; B = 8'hD6; #100;
A = 8'h1C; B = 8'hD7; #100;
A = 8'h1C; B = 8'hD8; #100;
A = 8'h1C; B = 8'hD9; #100;
A = 8'h1C; B = 8'hDA; #100;
A = 8'h1C; B = 8'hDB; #100;
A = 8'h1C; B = 8'hDC; #100;
A = 8'h1C; B = 8'hDD; #100;
A = 8'h1C; B = 8'hDE; #100;
A = 8'h1C; B = 8'hDF; #100;
A = 8'h1C; B = 8'hE0; #100;
A = 8'h1C; B = 8'hE1; #100;
A = 8'h1C; B = 8'hE2; #100;
A = 8'h1C; B = 8'hE3; #100;
A = 8'h1C; B = 8'hE4; #100;
A = 8'h1C; B = 8'hE5; #100;
A = 8'h1C; B = 8'hE6; #100;
A = 8'h1C; B = 8'hE7; #100;
A = 8'h1C; B = 8'hE8; #100;
A = 8'h1C; B = 8'hE9; #100;
A = 8'h1C; B = 8'hEA; #100;
A = 8'h1C; B = 8'hEB; #100;
A = 8'h1C; B = 8'hEC; #100;
A = 8'h1C; B = 8'hED; #100;
A = 8'h1C; B = 8'hEE; #100;
A = 8'h1C; B = 8'hEF; #100;
A = 8'h1C; B = 8'hF0; #100;
A = 8'h1C; B = 8'hF1; #100;
A = 8'h1C; B = 8'hF2; #100;
A = 8'h1C; B = 8'hF3; #100;
A = 8'h1C; B = 8'hF4; #100;
A = 8'h1C; B = 8'hF5; #100;
A = 8'h1C; B = 8'hF6; #100;
A = 8'h1C; B = 8'hF7; #100;
A = 8'h1C; B = 8'hF8; #100;
A = 8'h1C; B = 8'hF9; #100;
A = 8'h1C; B = 8'hFA; #100;
A = 8'h1C; B = 8'hFB; #100;
A = 8'h1C; B = 8'hFC; #100;
A = 8'h1C; B = 8'hFD; #100;
A = 8'h1C; B = 8'hFE; #100;
A = 8'h1C; B = 8'hFF; #100;
A = 8'h1D; B = 8'h0; #100;
A = 8'h1D; B = 8'h1; #100;
A = 8'h1D; B = 8'h2; #100;
A = 8'h1D; B = 8'h3; #100;
A = 8'h1D; B = 8'h4; #100;
A = 8'h1D; B = 8'h5; #100;
A = 8'h1D; B = 8'h6; #100;
A = 8'h1D; B = 8'h7; #100;
A = 8'h1D; B = 8'h8; #100;
A = 8'h1D; B = 8'h9; #100;
A = 8'h1D; B = 8'hA; #100;
A = 8'h1D; B = 8'hB; #100;
A = 8'h1D; B = 8'hC; #100;
A = 8'h1D; B = 8'hD; #100;
A = 8'h1D; B = 8'hE; #100;
A = 8'h1D; B = 8'hF; #100;
A = 8'h1D; B = 8'h10; #100;
A = 8'h1D; B = 8'h11; #100;
A = 8'h1D; B = 8'h12; #100;
A = 8'h1D; B = 8'h13; #100;
A = 8'h1D; B = 8'h14; #100;
A = 8'h1D; B = 8'h15; #100;
A = 8'h1D; B = 8'h16; #100;
A = 8'h1D; B = 8'h17; #100;
A = 8'h1D; B = 8'h18; #100;
A = 8'h1D; B = 8'h19; #100;
A = 8'h1D; B = 8'h1A; #100;
A = 8'h1D; B = 8'h1B; #100;
A = 8'h1D; B = 8'h1C; #100;
A = 8'h1D; B = 8'h1D; #100;
A = 8'h1D; B = 8'h1E; #100;
A = 8'h1D; B = 8'h1F; #100;
A = 8'h1D; B = 8'h20; #100;
A = 8'h1D; B = 8'h21; #100;
A = 8'h1D; B = 8'h22; #100;
A = 8'h1D; B = 8'h23; #100;
A = 8'h1D; B = 8'h24; #100;
A = 8'h1D; B = 8'h25; #100;
A = 8'h1D; B = 8'h26; #100;
A = 8'h1D; B = 8'h27; #100;
A = 8'h1D; B = 8'h28; #100;
A = 8'h1D; B = 8'h29; #100;
A = 8'h1D; B = 8'h2A; #100;
A = 8'h1D; B = 8'h2B; #100;
A = 8'h1D; B = 8'h2C; #100;
A = 8'h1D; B = 8'h2D; #100;
A = 8'h1D; B = 8'h2E; #100;
A = 8'h1D; B = 8'h2F; #100;
A = 8'h1D; B = 8'h30; #100;
A = 8'h1D; B = 8'h31; #100;
A = 8'h1D; B = 8'h32; #100;
A = 8'h1D; B = 8'h33; #100;
A = 8'h1D; B = 8'h34; #100;
A = 8'h1D; B = 8'h35; #100;
A = 8'h1D; B = 8'h36; #100;
A = 8'h1D; B = 8'h37; #100;
A = 8'h1D; B = 8'h38; #100;
A = 8'h1D; B = 8'h39; #100;
A = 8'h1D; B = 8'h3A; #100;
A = 8'h1D; B = 8'h3B; #100;
A = 8'h1D; B = 8'h3C; #100;
A = 8'h1D; B = 8'h3D; #100;
A = 8'h1D; B = 8'h3E; #100;
A = 8'h1D; B = 8'h3F; #100;
A = 8'h1D; B = 8'h40; #100;
A = 8'h1D; B = 8'h41; #100;
A = 8'h1D; B = 8'h42; #100;
A = 8'h1D; B = 8'h43; #100;
A = 8'h1D; B = 8'h44; #100;
A = 8'h1D; B = 8'h45; #100;
A = 8'h1D; B = 8'h46; #100;
A = 8'h1D; B = 8'h47; #100;
A = 8'h1D; B = 8'h48; #100;
A = 8'h1D; B = 8'h49; #100;
A = 8'h1D; B = 8'h4A; #100;
A = 8'h1D; B = 8'h4B; #100;
A = 8'h1D; B = 8'h4C; #100;
A = 8'h1D; B = 8'h4D; #100;
A = 8'h1D; B = 8'h4E; #100;
A = 8'h1D; B = 8'h4F; #100;
A = 8'h1D; B = 8'h50; #100;
A = 8'h1D; B = 8'h51; #100;
A = 8'h1D; B = 8'h52; #100;
A = 8'h1D; B = 8'h53; #100;
A = 8'h1D; B = 8'h54; #100;
A = 8'h1D; B = 8'h55; #100;
A = 8'h1D; B = 8'h56; #100;
A = 8'h1D; B = 8'h57; #100;
A = 8'h1D; B = 8'h58; #100;
A = 8'h1D; B = 8'h59; #100;
A = 8'h1D; B = 8'h5A; #100;
A = 8'h1D; B = 8'h5B; #100;
A = 8'h1D; B = 8'h5C; #100;
A = 8'h1D; B = 8'h5D; #100;
A = 8'h1D; B = 8'h5E; #100;
A = 8'h1D; B = 8'h5F; #100;
A = 8'h1D; B = 8'h60; #100;
A = 8'h1D; B = 8'h61; #100;
A = 8'h1D; B = 8'h62; #100;
A = 8'h1D; B = 8'h63; #100;
A = 8'h1D; B = 8'h64; #100;
A = 8'h1D; B = 8'h65; #100;
A = 8'h1D; B = 8'h66; #100;
A = 8'h1D; B = 8'h67; #100;
A = 8'h1D; B = 8'h68; #100;
A = 8'h1D; B = 8'h69; #100;
A = 8'h1D; B = 8'h6A; #100;
A = 8'h1D; B = 8'h6B; #100;
A = 8'h1D; B = 8'h6C; #100;
A = 8'h1D; B = 8'h6D; #100;
A = 8'h1D; B = 8'h6E; #100;
A = 8'h1D; B = 8'h6F; #100;
A = 8'h1D; B = 8'h70; #100;
A = 8'h1D; B = 8'h71; #100;
A = 8'h1D; B = 8'h72; #100;
A = 8'h1D; B = 8'h73; #100;
A = 8'h1D; B = 8'h74; #100;
A = 8'h1D; B = 8'h75; #100;
A = 8'h1D; B = 8'h76; #100;
A = 8'h1D; B = 8'h77; #100;
A = 8'h1D; B = 8'h78; #100;
A = 8'h1D; B = 8'h79; #100;
A = 8'h1D; B = 8'h7A; #100;
A = 8'h1D; B = 8'h7B; #100;
A = 8'h1D; B = 8'h7C; #100;
A = 8'h1D; B = 8'h7D; #100;
A = 8'h1D; B = 8'h7E; #100;
A = 8'h1D; B = 8'h7F; #100;
A = 8'h1D; B = 8'h80; #100;
A = 8'h1D; B = 8'h81; #100;
A = 8'h1D; B = 8'h82; #100;
A = 8'h1D; B = 8'h83; #100;
A = 8'h1D; B = 8'h84; #100;
A = 8'h1D; B = 8'h85; #100;
A = 8'h1D; B = 8'h86; #100;
A = 8'h1D; B = 8'h87; #100;
A = 8'h1D; B = 8'h88; #100;
A = 8'h1D; B = 8'h89; #100;
A = 8'h1D; B = 8'h8A; #100;
A = 8'h1D; B = 8'h8B; #100;
A = 8'h1D; B = 8'h8C; #100;
A = 8'h1D; B = 8'h8D; #100;
A = 8'h1D; B = 8'h8E; #100;
A = 8'h1D; B = 8'h8F; #100;
A = 8'h1D; B = 8'h90; #100;
A = 8'h1D; B = 8'h91; #100;
A = 8'h1D; B = 8'h92; #100;
A = 8'h1D; B = 8'h93; #100;
A = 8'h1D; B = 8'h94; #100;
A = 8'h1D; B = 8'h95; #100;
A = 8'h1D; B = 8'h96; #100;
A = 8'h1D; B = 8'h97; #100;
A = 8'h1D; B = 8'h98; #100;
A = 8'h1D; B = 8'h99; #100;
A = 8'h1D; B = 8'h9A; #100;
A = 8'h1D; B = 8'h9B; #100;
A = 8'h1D; B = 8'h9C; #100;
A = 8'h1D; B = 8'h9D; #100;
A = 8'h1D; B = 8'h9E; #100;
A = 8'h1D; B = 8'h9F; #100;
A = 8'h1D; B = 8'hA0; #100;
A = 8'h1D; B = 8'hA1; #100;
A = 8'h1D; B = 8'hA2; #100;
A = 8'h1D; B = 8'hA3; #100;
A = 8'h1D; B = 8'hA4; #100;
A = 8'h1D; B = 8'hA5; #100;
A = 8'h1D; B = 8'hA6; #100;
A = 8'h1D; B = 8'hA7; #100;
A = 8'h1D; B = 8'hA8; #100;
A = 8'h1D; B = 8'hA9; #100;
A = 8'h1D; B = 8'hAA; #100;
A = 8'h1D; B = 8'hAB; #100;
A = 8'h1D; B = 8'hAC; #100;
A = 8'h1D; B = 8'hAD; #100;
A = 8'h1D; B = 8'hAE; #100;
A = 8'h1D; B = 8'hAF; #100;
A = 8'h1D; B = 8'hB0; #100;
A = 8'h1D; B = 8'hB1; #100;
A = 8'h1D; B = 8'hB2; #100;
A = 8'h1D; B = 8'hB3; #100;
A = 8'h1D; B = 8'hB4; #100;
A = 8'h1D; B = 8'hB5; #100;
A = 8'h1D; B = 8'hB6; #100;
A = 8'h1D; B = 8'hB7; #100;
A = 8'h1D; B = 8'hB8; #100;
A = 8'h1D; B = 8'hB9; #100;
A = 8'h1D; B = 8'hBA; #100;
A = 8'h1D; B = 8'hBB; #100;
A = 8'h1D; B = 8'hBC; #100;
A = 8'h1D; B = 8'hBD; #100;
A = 8'h1D; B = 8'hBE; #100;
A = 8'h1D; B = 8'hBF; #100;
A = 8'h1D; B = 8'hC0; #100;
A = 8'h1D; B = 8'hC1; #100;
A = 8'h1D; B = 8'hC2; #100;
A = 8'h1D; B = 8'hC3; #100;
A = 8'h1D; B = 8'hC4; #100;
A = 8'h1D; B = 8'hC5; #100;
A = 8'h1D; B = 8'hC6; #100;
A = 8'h1D; B = 8'hC7; #100;
A = 8'h1D; B = 8'hC8; #100;
A = 8'h1D; B = 8'hC9; #100;
A = 8'h1D; B = 8'hCA; #100;
A = 8'h1D; B = 8'hCB; #100;
A = 8'h1D; B = 8'hCC; #100;
A = 8'h1D; B = 8'hCD; #100;
A = 8'h1D; B = 8'hCE; #100;
A = 8'h1D; B = 8'hCF; #100;
A = 8'h1D; B = 8'hD0; #100;
A = 8'h1D; B = 8'hD1; #100;
A = 8'h1D; B = 8'hD2; #100;
A = 8'h1D; B = 8'hD3; #100;
A = 8'h1D; B = 8'hD4; #100;
A = 8'h1D; B = 8'hD5; #100;
A = 8'h1D; B = 8'hD6; #100;
A = 8'h1D; B = 8'hD7; #100;
A = 8'h1D; B = 8'hD8; #100;
A = 8'h1D; B = 8'hD9; #100;
A = 8'h1D; B = 8'hDA; #100;
A = 8'h1D; B = 8'hDB; #100;
A = 8'h1D; B = 8'hDC; #100;
A = 8'h1D; B = 8'hDD; #100;
A = 8'h1D; B = 8'hDE; #100;
A = 8'h1D; B = 8'hDF; #100;
A = 8'h1D; B = 8'hE0; #100;
A = 8'h1D; B = 8'hE1; #100;
A = 8'h1D; B = 8'hE2; #100;
A = 8'h1D; B = 8'hE3; #100;
A = 8'h1D; B = 8'hE4; #100;
A = 8'h1D; B = 8'hE5; #100;
A = 8'h1D; B = 8'hE6; #100;
A = 8'h1D; B = 8'hE7; #100;
A = 8'h1D; B = 8'hE8; #100;
A = 8'h1D; B = 8'hE9; #100;
A = 8'h1D; B = 8'hEA; #100;
A = 8'h1D; B = 8'hEB; #100;
A = 8'h1D; B = 8'hEC; #100;
A = 8'h1D; B = 8'hED; #100;
A = 8'h1D; B = 8'hEE; #100;
A = 8'h1D; B = 8'hEF; #100;
A = 8'h1D; B = 8'hF0; #100;
A = 8'h1D; B = 8'hF1; #100;
A = 8'h1D; B = 8'hF2; #100;
A = 8'h1D; B = 8'hF3; #100;
A = 8'h1D; B = 8'hF4; #100;
A = 8'h1D; B = 8'hF5; #100;
A = 8'h1D; B = 8'hF6; #100;
A = 8'h1D; B = 8'hF7; #100;
A = 8'h1D; B = 8'hF8; #100;
A = 8'h1D; B = 8'hF9; #100;
A = 8'h1D; B = 8'hFA; #100;
A = 8'h1D; B = 8'hFB; #100;
A = 8'h1D; B = 8'hFC; #100;
A = 8'h1D; B = 8'hFD; #100;
A = 8'h1D; B = 8'hFE; #100;
A = 8'h1D; B = 8'hFF; #100;
A = 8'h1E; B = 8'h0; #100;
A = 8'h1E; B = 8'h1; #100;
A = 8'h1E; B = 8'h2; #100;
A = 8'h1E; B = 8'h3; #100;
A = 8'h1E; B = 8'h4; #100;
A = 8'h1E; B = 8'h5; #100;
A = 8'h1E; B = 8'h6; #100;
A = 8'h1E; B = 8'h7; #100;
A = 8'h1E; B = 8'h8; #100;
A = 8'h1E; B = 8'h9; #100;
A = 8'h1E; B = 8'hA; #100;
A = 8'h1E; B = 8'hB; #100;
A = 8'h1E; B = 8'hC; #100;
A = 8'h1E; B = 8'hD; #100;
A = 8'h1E; B = 8'hE; #100;
A = 8'h1E; B = 8'hF; #100;
A = 8'h1E; B = 8'h10; #100;
A = 8'h1E; B = 8'h11; #100;
A = 8'h1E; B = 8'h12; #100;
A = 8'h1E; B = 8'h13; #100;
A = 8'h1E; B = 8'h14; #100;
A = 8'h1E; B = 8'h15; #100;
A = 8'h1E; B = 8'h16; #100;
A = 8'h1E; B = 8'h17; #100;
A = 8'h1E; B = 8'h18; #100;
A = 8'h1E; B = 8'h19; #100;
A = 8'h1E; B = 8'h1A; #100;
A = 8'h1E; B = 8'h1B; #100;
A = 8'h1E; B = 8'h1C; #100;
A = 8'h1E; B = 8'h1D; #100;
A = 8'h1E; B = 8'h1E; #100;
A = 8'h1E; B = 8'h1F; #100;
A = 8'h1E; B = 8'h20; #100;
A = 8'h1E; B = 8'h21; #100;
A = 8'h1E; B = 8'h22; #100;
A = 8'h1E; B = 8'h23; #100;
A = 8'h1E; B = 8'h24; #100;
A = 8'h1E; B = 8'h25; #100;
A = 8'h1E; B = 8'h26; #100;
A = 8'h1E; B = 8'h27; #100;
A = 8'h1E; B = 8'h28; #100;
A = 8'h1E; B = 8'h29; #100;
A = 8'h1E; B = 8'h2A; #100;
A = 8'h1E; B = 8'h2B; #100;
A = 8'h1E; B = 8'h2C; #100;
A = 8'h1E; B = 8'h2D; #100;
A = 8'h1E; B = 8'h2E; #100;
A = 8'h1E; B = 8'h2F; #100;
A = 8'h1E; B = 8'h30; #100;
A = 8'h1E; B = 8'h31; #100;
A = 8'h1E; B = 8'h32; #100;
A = 8'h1E; B = 8'h33; #100;
A = 8'h1E; B = 8'h34; #100;
A = 8'h1E; B = 8'h35; #100;
A = 8'h1E; B = 8'h36; #100;
A = 8'h1E; B = 8'h37; #100;
A = 8'h1E; B = 8'h38; #100;
A = 8'h1E; B = 8'h39; #100;
A = 8'h1E; B = 8'h3A; #100;
A = 8'h1E; B = 8'h3B; #100;
A = 8'h1E; B = 8'h3C; #100;
A = 8'h1E; B = 8'h3D; #100;
A = 8'h1E; B = 8'h3E; #100;
A = 8'h1E; B = 8'h3F; #100;
A = 8'h1E; B = 8'h40; #100;
A = 8'h1E; B = 8'h41; #100;
A = 8'h1E; B = 8'h42; #100;
A = 8'h1E; B = 8'h43; #100;
A = 8'h1E; B = 8'h44; #100;
A = 8'h1E; B = 8'h45; #100;
A = 8'h1E; B = 8'h46; #100;
A = 8'h1E; B = 8'h47; #100;
A = 8'h1E; B = 8'h48; #100;
A = 8'h1E; B = 8'h49; #100;
A = 8'h1E; B = 8'h4A; #100;
A = 8'h1E; B = 8'h4B; #100;
A = 8'h1E; B = 8'h4C; #100;
A = 8'h1E; B = 8'h4D; #100;
A = 8'h1E; B = 8'h4E; #100;
A = 8'h1E; B = 8'h4F; #100;
A = 8'h1E; B = 8'h50; #100;
A = 8'h1E; B = 8'h51; #100;
A = 8'h1E; B = 8'h52; #100;
A = 8'h1E; B = 8'h53; #100;
A = 8'h1E; B = 8'h54; #100;
A = 8'h1E; B = 8'h55; #100;
A = 8'h1E; B = 8'h56; #100;
A = 8'h1E; B = 8'h57; #100;
A = 8'h1E; B = 8'h58; #100;
A = 8'h1E; B = 8'h59; #100;
A = 8'h1E; B = 8'h5A; #100;
A = 8'h1E; B = 8'h5B; #100;
A = 8'h1E; B = 8'h5C; #100;
A = 8'h1E; B = 8'h5D; #100;
A = 8'h1E; B = 8'h5E; #100;
A = 8'h1E; B = 8'h5F; #100;
A = 8'h1E; B = 8'h60; #100;
A = 8'h1E; B = 8'h61; #100;
A = 8'h1E; B = 8'h62; #100;
A = 8'h1E; B = 8'h63; #100;
A = 8'h1E; B = 8'h64; #100;
A = 8'h1E; B = 8'h65; #100;
A = 8'h1E; B = 8'h66; #100;
A = 8'h1E; B = 8'h67; #100;
A = 8'h1E; B = 8'h68; #100;
A = 8'h1E; B = 8'h69; #100;
A = 8'h1E; B = 8'h6A; #100;
A = 8'h1E; B = 8'h6B; #100;
A = 8'h1E; B = 8'h6C; #100;
A = 8'h1E; B = 8'h6D; #100;
A = 8'h1E; B = 8'h6E; #100;
A = 8'h1E; B = 8'h6F; #100;
A = 8'h1E; B = 8'h70; #100;
A = 8'h1E; B = 8'h71; #100;
A = 8'h1E; B = 8'h72; #100;
A = 8'h1E; B = 8'h73; #100;
A = 8'h1E; B = 8'h74; #100;
A = 8'h1E; B = 8'h75; #100;
A = 8'h1E; B = 8'h76; #100;
A = 8'h1E; B = 8'h77; #100;
A = 8'h1E; B = 8'h78; #100;
A = 8'h1E; B = 8'h79; #100;
A = 8'h1E; B = 8'h7A; #100;
A = 8'h1E; B = 8'h7B; #100;
A = 8'h1E; B = 8'h7C; #100;
A = 8'h1E; B = 8'h7D; #100;
A = 8'h1E; B = 8'h7E; #100;
A = 8'h1E; B = 8'h7F; #100;
A = 8'h1E; B = 8'h80; #100;
A = 8'h1E; B = 8'h81; #100;
A = 8'h1E; B = 8'h82; #100;
A = 8'h1E; B = 8'h83; #100;
A = 8'h1E; B = 8'h84; #100;
A = 8'h1E; B = 8'h85; #100;
A = 8'h1E; B = 8'h86; #100;
A = 8'h1E; B = 8'h87; #100;
A = 8'h1E; B = 8'h88; #100;
A = 8'h1E; B = 8'h89; #100;
A = 8'h1E; B = 8'h8A; #100;
A = 8'h1E; B = 8'h8B; #100;
A = 8'h1E; B = 8'h8C; #100;
A = 8'h1E; B = 8'h8D; #100;
A = 8'h1E; B = 8'h8E; #100;
A = 8'h1E; B = 8'h8F; #100;
A = 8'h1E; B = 8'h90; #100;
A = 8'h1E; B = 8'h91; #100;
A = 8'h1E; B = 8'h92; #100;
A = 8'h1E; B = 8'h93; #100;
A = 8'h1E; B = 8'h94; #100;
A = 8'h1E; B = 8'h95; #100;
A = 8'h1E; B = 8'h96; #100;
A = 8'h1E; B = 8'h97; #100;
A = 8'h1E; B = 8'h98; #100;
A = 8'h1E; B = 8'h99; #100;
A = 8'h1E; B = 8'h9A; #100;
A = 8'h1E; B = 8'h9B; #100;
A = 8'h1E; B = 8'h9C; #100;
A = 8'h1E; B = 8'h9D; #100;
A = 8'h1E; B = 8'h9E; #100;
A = 8'h1E; B = 8'h9F; #100;
A = 8'h1E; B = 8'hA0; #100;
A = 8'h1E; B = 8'hA1; #100;
A = 8'h1E; B = 8'hA2; #100;
A = 8'h1E; B = 8'hA3; #100;
A = 8'h1E; B = 8'hA4; #100;
A = 8'h1E; B = 8'hA5; #100;
A = 8'h1E; B = 8'hA6; #100;
A = 8'h1E; B = 8'hA7; #100;
A = 8'h1E; B = 8'hA8; #100;
A = 8'h1E; B = 8'hA9; #100;
A = 8'h1E; B = 8'hAA; #100;
A = 8'h1E; B = 8'hAB; #100;
A = 8'h1E; B = 8'hAC; #100;
A = 8'h1E; B = 8'hAD; #100;
A = 8'h1E; B = 8'hAE; #100;
A = 8'h1E; B = 8'hAF; #100;
A = 8'h1E; B = 8'hB0; #100;
A = 8'h1E; B = 8'hB1; #100;
A = 8'h1E; B = 8'hB2; #100;
A = 8'h1E; B = 8'hB3; #100;
A = 8'h1E; B = 8'hB4; #100;
A = 8'h1E; B = 8'hB5; #100;
A = 8'h1E; B = 8'hB6; #100;
A = 8'h1E; B = 8'hB7; #100;
A = 8'h1E; B = 8'hB8; #100;
A = 8'h1E; B = 8'hB9; #100;
A = 8'h1E; B = 8'hBA; #100;
A = 8'h1E; B = 8'hBB; #100;
A = 8'h1E; B = 8'hBC; #100;
A = 8'h1E; B = 8'hBD; #100;
A = 8'h1E; B = 8'hBE; #100;
A = 8'h1E; B = 8'hBF; #100;
A = 8'h1E; B = 8'hC0; #100;
A = 8'h1E; B = 8'hC1; #100;
A = 8'h1E; B = 8'hC2; #100;
A = 8'h1E; B = 8'hC3; #100;
A = 8'h1E; B = 8'hC4; #100;
A = 8'h1E; B = 8'hC5; #100;
A = 8'h1E; B = 8'hC6; #100;
A = 8'h1E; B = 8'hC7; #100;
A = 8'h1E; B = 8'hC8; #100;
A = 8'h1E; B = 8'hC9; #100;
A = 8'h1E; B = 8'hCA; #100;
A = 8'h1E; B = 8'hCB; #100;
A = 8'h1E; B = 8'hCC; #100;
A = 8'h1E; B = 8'hCD; #100;
A = 8'h1E; B = 8'hCE; #100;
A = 8'h1E; B = 8'hCF; #100;
A = 8'h1E; B = 8'hD0; #100;
A = 8'h1E; B = 8'hD1; #100;
A = 8'h1E; B = 8'hD2; #100;
A = 8'h1E; B = 8'hD3; #100;
A = 8'h1E; B = 8'hD4; #100;
A = 8'h1E; B = 8'hD5; #100;
A = 8'h1E; B = 8'hD6; #100;
A = 8'h1E; B = 8'hD7; #100;
A = 8'h1E; B = 8'hD8; #100;
A = 8'h1E; B = 8'hD9; #100;
A = 8'h1E; B = 8'hDA; #100;
A = 8'h1E; B = 8'hDB; #100;
A = 8'h1E; B = 8'hDC; #100;
A = 8'h1E; B = 8'hDD; #100;
A = 8'h1E; B = 8'hDE; #100;
A = 8'h1E; B = 8'hDF; #100;
A = 8'h1E; B = 8'hE0; #100;
A = 8'h1E; B = 8'hE1; #100;
A = 8'h1E; B = 8'hE2; #100;
A = 8'h1E; B = 8'hE3; #100;
A = 8'h1E; B = 8'hE4; #100;
A = 8'h1E; B = 8'hE5; #100;
A = 8'h1E; B = 8'hE6; #100;
A = 8'h1E; B = 8'hE7; #100;
A = 8'h1E; B = 8'hE8; #100;
A = 8'h1E; B = 8'hE9; #100;
A = 8'h1E; B = 8'hEA; #100;
A = 8'h1E; B = 8'hEB; #100;
A = 8'h1E; B = 8'hEC; #100;
A = 8'h1E; B = 8'hED; #100;
A = 8'h1E; B = 8'hEE; #100;
A = 8'h1E; B = 8'hEF; #100;
A = 8'h1E; B = 8'hF0; #100;
A = 8'h1E; B = 8'hF1; #100;
A = 8'h1E; B = 8'hF2; #100;
A = 8'h1E; B = 8'hF3; #100;
A = 8'h1E; B = 8'hF4; #100;
A = 8'h1E; B = 8'hF5; #100;
A = 8'h1E; B = 8'hF6; #100;
A = 8'h1E; B = 8'hF7; #100;
A = 8'h1E; B = 8'hF8; #100;
A = 8'h1E; B = 8'hF9; #100;
A = 8'h1E; B = 8'hFA; #100;
A = 8'h1E; B = 8'hFB; #100;
A = 8'h1E; B = 8'hFC; #100;
A = 8'h1E; B = 8'hFD; #100;
A = 8'h1E; B = 8'hFE; #100;
A = 8'h1E; B = 8'hFF; #100;
A = 8'h1F; B = 8'h0; #100;
A = 8'h1F; B = 8'h1; #100;
A = 8'h1F; B = 8'h2; #100;
A = 8'h1F; B = 8'h3; #100;
A = 8'h1F; B = 8'h4; #100;
A = 8'h1F; B = 8'h5; #100;
A = 8'h1F; B = 8'h6; #100;
A = 8'h1F; B = 8'h7; #100;
A = 8'h1F; B = 8'h8; #100;
A = 8'h1F; B = 8'h9; #100;
A = 8'h1F; B = 8'hA; #100;
A = 8'h1F; B = 8'hB; #100;
A = 8'h1F; B = 8'hC; #100;
A = 8'h1F; B = 8'hD; #100;
A = 8'h1F; B = 8'hE; #100;
A = 8'h1F; B = 8'hF; #100;
A = 8'h1F; B = 8'h10; #100;
A = 8'h1F; B = 8'h11; #100;
A = 8'h1F; B = 8'h12; #100;
A = 8'h1F; B = 8'h13; #100;
A = 8'h1F; B = 8'h14; #100;
A = 8'h1F; B = 8'h15; #100;
A = 8'h1F; B = 8'h16; #100;
A = 8'h1F; B = 8'h17; #100;
A = 8'h1F; B = 8'h18; #100;
A = 8'h1F; B = 8'h19; #100;
A = 8'h1F; B = 8'h1A; #100;
A = 8'h1F; B = 8'h1B; #100;
A = 8'h1F; B = 8'h1C; #100;
A = 8'h1F; B = 8'h1D; #100;
A = 8'h1F; B = 8'h1E; #100;
A = 8'h1F; B = 8'h1F; #100;
A = 8'h1F; B = 8'h20; #100;
A = 8'h1F; B = 8'h21; #100;
A = 8'h1F; B = 8'h22; #100;
A = 8'h1F; B = 8'h23; #100;
A = 8'h1F; B = 8'h24; #100;
A = 8'h1F; B = 8'h25; #100;
A = 8'h1F; B = 8'h26; #100;
A = 8'h1F; B = 8'h27; #100;
A = 8'h1F; B = 8'h28; #100;
A = 8'h1F; B = 8'h29; #100;
A = 8'h1F; B = 8'h2A; #100;
A = 8'h1F; B = 8'h2B; #100;
A = 8'h1F; B = 8'h2C; #100;
A = 8'h1F; B = 8'h2D; #100;
A = 8'h1F; B = 8'h2E; #100;
A = 8'h1F; B = 8'h2F; #100;
A = 8'h1F; B = 8'h30; #100;
A = 8'h1F; B = 8'h31; #100;
A = 8'h1F; B = 8'h32; #100;
A = 8'h1F; B = 8'h33; #100;
A = 8'h1F; B = 8'h34; #100;
A = 8'h1F; B = 8'h35; #100;
A = 8'h1F; B = 8'h36; #100;
A = 8'h1F; B = 8'h37; #100;
A = 8'h1F; B = 8'h38; #100;
A = 8'h1F; B = 8'h39; #100;
A = 8'h1F; B = 8'h3A; #100;
A = 8'h1F; B = 8'h3B; #100;
A = 8'h1F; B = 8'h3C; #100;
A = 8'h1F; B = 8'h3D; #100;
A = 8'h1F; B = 8'h3E; #100;
A = 8'h1F; B = 8'h3F; #100;
A = 8'h1F; B = 8'h40; #100;
A = 8'h1F; B = 8'h41; #100;
A = 8'h1F; B = 8'h42; #100;
A = 8'h1F; B = 8'h43; #100;
A = 8'h1F; B = 8'h44; #100;
A = 8'h1F; B = 8'h45; #100;
A = 8'h1F; B = 8'h46; #100;
A = 8'h1F; B = 8'h47; #100;
A = 8'h1F; B = 8'h48; #100;
A = 8'h1F; B = 8'h49; #100;
A = 8'h1F; B = 8'h4A; #100;
A = 8'h1F; B = 8'h4B; #100;
A = 8'h1F; B = 8'h4C; #100;
A = 8'h1F; B = 8'h4D; #100;
A = 8'h1F; B = 8'h4E; #100;
A = 8'h1F; B = 8'h4F; #100;
A = 8'h1F; B = 8'h50; #100;
A = 8'h1F; B = 8'h51; #100;
A = 8'h1F; B = 8'h52; #100;
A = 8'h1F; B = 8'h53; #100;
A = 8'h1F; B = 8'h54; #100;
A = 8'h1F; B = 8'h55; #100;
A = 8'h1F; B = 8'h56; #100;
A = 8'h1F; B = 8'h57; #100;
A = 8'h1F; B = 8'h58; #100;
A = 8'h1F; B = 8'h59; #100;
A = 8'h1F; B = 8'h5A; #100;
A = 8'h1F; B = 8'h5B; #100;
A = 8'h1F; B = 8'h5C; #100;
A = 8'h1F; B = 8'h5D; #100;
A = 8'h1F; B = 8'h5E; #100;
A = 8'h1F; B = 8'h5F; #100;
A = 8'h1F; B = 8'h60; #100;
A = 8'h1F; B = 8'h61; #100;
A = 8'h1F; B = 8'h62; #100;
A = 8'h1F; B = 8'h63; #100;
A = 8'h1F; B = 8'h64; #100;
A = 8'h1F; B = 8'h65; #100;
A = 8'h1F; B = 8'h66; #100;
A = 8'h1F; B = 8'h67; #100;
A = 8'h1F; B = 8'h68; #100;
A = 8'h1F; B = 8'h69; #100;
A = 8'h1F; B = 8'h6A; #100;
A = 8'h1F; B = 8'h6B; #100;
A = 8'h1F; B = 8'h6C; #100;
A = 8'h1F; B = 8'h6D; #100;
A = 8'h1F; B = 8'h6E; #100;
A = 8'h1F; B = 8'h6F; #100;
A = 8'h1F; B = 8'h70; #100;
A = 8'h1F; B = 8'h71; #100;
A = 8'h1F; B = 8'h72; #100;
A = 8'h1F; B = 8'h73; #100;
A = 8'h1F; B = 8'h74; #100;
A = 8'h1F; B = 8'h75; #100;
A = 8'h1F; B = 8'h76; #100;
A = 8'h1F; B = 8'h77; #100;
A = 8'h1F; B = 8'h78; #100;
A = 8'h1F; B = 8'h79; #100;
A = 8'h1F; B = 8'h7A; #100;
A = 8'h1F; B = 8'h7B; #100;
A = 8'h1F; B = 8'h7C; #100;
A = 8'h1F; B = 8'h7D; #100;
A = 8'h1F; B = 8'h7E; #100;
A = 8'h1F; B = 8'h7F; #100;
A = 8'h1F; B = 8'h80; #100;
A = 8'h1F; B = 8'h81; #100;
A = 8'h1F; B = 8'h82; #100;
A = 8'h1F; B = 8'h83; #100;
A = 8'h1F; B = 8'h84; #100;
A = 8'h1F; B = 8'h85; #100;
A = 8'h1F; B = 8'h86; #100;
A = 8'h1F; B = 8'h87; #100;
A = 8'h1F; B = 8'h88; #100;
A = 8'h1F; B = 8'h89; #100;
A = 8'h1F; B = 8'h8A; #100;
A = 8'h1F; B = 8'h8B; #100;
A = 8'h1F; B = 8'h8C; #100;
A = 8'h1F; B = 8'h8D; #100;
A = 8'h1F; B = 8'h8E; #100;
A = 8'h1F; B = 8'h8F; #100;
A = 8'h1F; B = 8'h90; #100;
A = 8'h1F; B = 8'h91; #100;
A = 8'h1F; B = 8'h92; #100;
A = 8'h1F; B = 8'h93; #100;
A = 8'h1F; B = 8'h94; #100;
A = 8'h1F; B = 8'h95; #100;
A = 8'h1F; B = 8'h96; #100;
A = 8'h1F; B = 8'h97; #100;
A = 8'h1F; B = 8'h98; #100;
A = 8'h1F; B = 8'h99; #100;
A = 8'h1F; B = 8'h9A; #100;
A = 8'h1F; B = 8'h9B; #100;
A = 8'h1F; B = 8'h9C; #100;
A = 8'h1F; B = 8'h9D; #100;
A = 8'h1F; B = 8'h9E; #100;
A = 8'h1F; B = 8'h9F; #100;
A = 8'h1F; B = 8'hA0; #100;
A = 8'h1F; B = 8'hA1; #100;
A = 8'h1F; B = 8'hA2; #100;
A = 8'h1F; B = 8'hA3; #100;
A = 8'h1F; B = 8'hA4; #100;
A = 8'h1F; B = 8'hA5; #100;
A = 8'h1F; B = 8'hA6; #100;
A = 8'h1F; B = 8'hA7; #100;
A = 8'h1F; B = 8'hA8; #100;
A = 8'h1F; B = 8'hA9; #100;
A = 8'h1F; B = 8'hAA; #100;
A = 8'h1F; B = 8'hAB; #100;
A = 8'h1F; B = 8'hAC; #100;
A = 8'h1F; B = 8'hAD; #100;
A = 8'h1F; B = 8'hAE; #100;
A = 8'h1F; B = 8'hAF; #100;
A = 8'h1F; B = 8'hB0; #100;
A = 8'h1F; B = 8'hB1; #100;
A = 8'h1F; B = 8'hB2; #100;
A = 8'h1F; B = 8'hB3; #100;
A = 8'h1F; B = 8'hB4; #100;
A = 8'h1F; B = 8'hB5; #100;
A = 8'h1F; B = 8'hB6; #100;
A = 8'h1F; B = 8'hB7; #100;
A = 8'h1F; B = 8'hB8; #100;
A = 8'h1F; B = 8'hB9; #100;
A = 8'h1F; B = 8'hBA; #100;
A = 8'h1F; B = 8'hBB; #100;
A = 8'h1F; B = 8'hBC; #100;
A = 8'h1F; B = 8'hBD; #100;
A = 8'h1F; B = 8'hBE; #100;
A = 8'h1F; B = 8'hBF; #100;
A = 8'h1F; B = 8'hC0; #100;
A = 8'h1F; B = 8'hC1; #100;
A = 8'h1F; B = 8'hC2; #100;
A = 8'h1F; B = 8'hC3; #100;
A = 8'h1F; B = 8'hC4; #100;
A = 8'h1F; B = 8'hC5; #100;
A = 8'h1F; B = 8'hC6; #100;
A = 8'h1F; B = 8'hC7; #100;
A = 8'h1F; B = 8'hC8; #100;
A = 8'h1F; B = 8'hC9; #100;
A = 8'h1F; B = 8'hCA; #100;
A = 8'h1F; B = 8'hCB; #100;
A = 8'h1F; B = 8'hCC; #100;
A = 8'h1F; B = 8'hCD; #100;
A = 8'h1F; B = 8'hCE; #100;
A = 8'h1F; B = 8'hCF; #100;
A = 8'h1F; B = 8'hD0; #100;
A = 8'h1F; B = 8'hD1; #100;
A = 8'h1F; B = 8'hD2; #100;
A = 8'h1F; B = 8'hD3; #100;
A = 8'h1F; B = 8'hD4; #100;
A = 8'h1F; B = 8'hD5; #100;
A = 8'h1F; B = 8'hD6; #100;
A = 8'h1F; B = 8'hD7; #100;
A = 8'h1F; B = 8'hD8; #100;
A = 8'h1F; B = 8'hD9; #100;
A = 8'h1F; B = 8'hDA; #100;
A = 8'h1F; B = 8'hDB; #100;
A = 8'h1F; B = 8'hDC; #100;
A = 8'h1F; B = 8'hDD; #100;
A = 8'h1F; B = 8'hDE; #100;
A = 8'h1F; B = 8'hDF; #100;
A = 8'h1F; B = 8'hE0; #100;
A = 8'h1F; B = 8'hE1; #100;
A = 8'h1F; B = 8'hE2; #100;
A = 8'h1F; B = 8'hE3; #100;
A = 8'h1F; B = 8'hE4; #100;
A = 8'h1F; B = 8'hE5; #100;
A = 8'h1F; B = 8'hE6; #100;
A = 8'h1F; B = 8'hE7; #100;
A = 8'h1F; B = 8'hE8; #100;
A = 8'h1F; B = 8'hE9; #100;
A = 8'h1F; B = 8'hEA; #100;
A = 8'h1F; B = 8'hEB; #100;
A = 8'h1F; B = 8'hEC; #100;
A = 8'h1F; B = 8'hED; #100;
A = 8'h1F; B = 8'hEE; #100;
A = 8'h1F; B = 8'hEF; #100;
A = 8'h1F; B = 8'hF0; #100;
A = 8'h1F; B = 8'hF1; #100;
A = 8'h1F; B = 8'hF2; #100;
A = 8'h1F; B = 8'hF3; #100;
A = 8'h1F; B = 8'hF4; #100;
A = 8'h1F; B = 8'hF5; #100;
A = 8'h1F; B = 8'hF6; #100;
A = 8'h1F; B = 8'hF7; #100;
A = 8'h1F; B = 8'hF8; #100;
A = 8'h1F; B = 8'hF9; #100;
A = 8'h1F; B = 8'hFA; #100;
A = 8'h1F; B = 8'hFB; #100;
A = 8'h1F; B = 8'hFC; #100;
A = 8'h1F; B = 8'hFD; #100;
A = 8'h1F; B = 8'hFE; #100;
A = 8'h1F; B = 8'hFF; #100;
A = 8'h20; B = 8'h0; #100;
A = 8'h20; B = 8'h1; #100;
A = 8'h20; B = 8'h2; #100;
A = 8'h20; B = 8'h3; #100;
A = 8'h20; B = 8'h4; #100;
A = 8'h20; B = 8'h5; #100;
A = 8'h20; B = 8'h6; #100;
A = 8'h20; B = 8'h7; #100;
A = 8'h20; B = 8'h8; #100;
A = 8'h20; B = 8'h9; #100;
A = 8'h20; B = 8'hA; #100;
A = 8'h20; B = 8'hB; #100;
A = 8'h20; B = 8'hC; #100;
A = 8'h20; B = 8'hD; #100;
A = 8'h20; B = 8'hE; #100;
A = 8'h20; B = 8'hF; #100;
A = 8'h20; B = 8'h10; #100;
A = 8'h20; B = 8'h11; #100;
A = 8'h20; B = 8'h12; #100;
A = 8'h20; B = 8'h13; #100;
A = 8'h20; B = 8'h14; #100;
A = 8'h20; B = 8'h15; #100;
A = 8'h20; B = 8'h16; #100;
A = 8'h20; B = 8'h17; #100;
A = 8'h20; B = 8'h18; #100;
A = 8'h20; B = 8'h19; #100;
A = 8'h20; B = 8'h1A; #100;
A = 8'h20; B = 8'h1B; #100;
A = 8'h20; B = 8'h1C; #100;
A = 8'h20; B = 8'h1D; #100;
A = 8'h20; B = 8'h1E; #100;
A = 8'h20; B = 8'h1F; #100;
A = 8'h20; B = 8'h20; #100;
A = 8'h20; B = 8'h21; #100;
A = 8'h20; B = 8'h22; #100;
A = 8'h20; B = 8'h23; #100;
A = 8'h20; B = 8'h24; #100;
A = 8'h20; B = 8'h25; #100;
A = 8'h20; B = 8'h26; #100;
A = 8'h20; B = 8'h27; #100;
A = 8'h20; B = 8'h28; #100;
A = 8'h20; B = 8'h29; #100;
A = 8'h20; B = 8'h2A; #100;
A = 8'h20; B = 8'h2B; #100;
A = 8'h20; B = 8'h2C; #100;
A = 8'h20; B = 8'h2D; #100;
A = 8'h20; B = 8'h2E; #100;
A = 8'h20; B = 8'h2F; #100;
A = 8'h20; B = 8'h30; #100;
A = 8'h20; B = 8'h31; #100;
A = 8'h20; B = 8'h32; #100;
A = 8'h20; B = 8'h33; #100;
A = 8'h20; B = 8'h34; #100;
A = 8'h20; B = 8'h35; #100;
A = 8'h20; B = 8'h36; #100;
A = 8'h20; B = 8'h37; #100;
A = 8'h20; B = 8'h38; #100;
A = 8'h20; B = 8'h39; #100;
A = 8'h20; B = 8'h3A; #100;
A = 8'h20; B = 8'h3B; #100;
A = 8'h20; B = 8'h3C; #100;
A = 8'h20; B = 8'h3D; #100;
A = 8'h20; B = 8'h3E; #100;
A = 8'h20; B = 8'h3F; #100;
A = 8'h20; B = 8'h40; #100;
A = 8'h20; B = 8'h41; #100;
A = 8'h20; B = 8'h42; #100;
A = 8'h20; B = 8'h43; #100;
A = 8'h20; B = 8'h44; #100;
A = 8'h20; B = 8'h45; #100;
A = 8'h20; B = 8'h46; #100;
A = 8'h20; B = 8'h47; #100;
A = 8'h20; B = 8'h48; #100;
A = 8'h20; B = 8'h49; #100;
A = 8'h20; B = 8'h4A; #100;
A = 8'h20; B = 8'h4B; #100;
A = 8'h20; B = 8'h4C; #100;
A = 8'h20; B = 8'h4D; #100;
A = 8'h20; B = 8'h4E; #100;
A = 8'h20; B = 8'h4F; #100;
A = 8'h20; B = 8'h50; #100;
A = 8'h20; B = 8'h51; #100;
A = 8'h20; B = 8'h52; #100;
A = 8'h20; B = 8'h53; #100;
A = 8'h20; B = 8'h54; #100;
A = 8'h20; B = 8'h55; #100;
A = 8'h20; B = 8'h56; #100;
A = 8'h20; B = 8'h57; #100;
A = 8'h20; B = 8'h58; #100;
A = 8'h20; B = 8'h59; #100;
A = 8'h20; B = 8'h5A; #100;
A = 8'h20; B = 8'h5B; #100;
A = 8'h20; B = 8'h5C; #100;
A = 8'h20; B = 8'h5D; #100;
A = 8'h20; B = 8'h5E; #100;
A = 8'h20; B = 8'h5F; #100;
A = 8'h20; B = 8'h60; #100;
A = 8'h20; B = 8'h61; #100;
A = 8'h20; B = 8'h62; #100;
A = 8'h20; B = 8'h63; #100;
A = 8'h20; B = 8'h64; #100;
A = 8'h20; B = 8'h65; #100;
A = 8'h20; B = 8'h66; #100;
A = 8'h20; B = 8'h67; #100;
A = 8'h20; B = 8'h68; #100;
A = 8'h20; B = 8'h69; #100;
A = 8'h20; B = 8'h6A; #100;
A = 8'h20; B = 8'h6B; #100;
A = 8'h20; B = 8'h6C; #100;
A = 8'h20; B = 8'h6D; #100;
A = 8'h20; B = 8'h6E; #100;
A = 8'h20; B = 8'h6F; #100;
A = 8'h20; B = 8'h70; #100;
A = 8'h20; B = 8'h71; #100;
A = 8'h20; B = 8'h72; #100;
A = 8'h20; B = 8'h73; #100;
A = 8'h20; B = 8'h74; #100;
A = 8'h20; B = 8'h75; #100;
A = 8'h20; B = 8'h76; #100;
A = 8'h20; B = 8'h77; #100;
A = 8'h20; B = 8'h78; #100;
A = 8'h20; B = 8'h79; #100;
A = 8'h20; B = 8'h7A; #100;
A = 8'h20; B = 8'h7B; #100;
A = 8'h20; B = 8'h7C; #100;
A = 8'h20; B = 8'h7D; #100;
A = 8'h20; B = 8'h7E; #100;
A = 8'h20; B = 8'h7F; #100;
A = 8'h20; B = 8'h80; #100;
A = 8'h20; B = 8'h81; #100;
A = 8'h20; B = 8'h82; #100;
A = 8'h20; B = 8'h83; #100;
A = 8'h20; B = 8'h84; #100;
A = 8'h20; B = 8'h85; #100;
A = 8'h20; B = 8'h86; #100;
A = 8'h20; B = 8'h87; #100;
A = 8'h20; B = 8'h88; #100;
A = 8'h20; B = 8'h89; #100;
A = 8'h20; B = 8'h8A; #100;
A = 8'h20; B = 8'h8B; #100;
A = 8'h20; B = 8'h8C; #100;
A = 8'h20; B = 8'h8D; #100;
A = 8'h20; B = 8'h8E; #100;
A = 8'h20; B = 8'h8F; #100;
A = 8'h20; B = 8'h90; #100;
A = 8'h20; B = 8'h91; #100;
A = 8'h20; B = 8'h92; #100;
A = 8'h20; B = 8'h93; #100;
A = 8'h20; B = 8'h94; #100;
A = 8'h20; B = 8'h95; #100;
A = 8'h20; B = 8'h96; #100;
A = 8'h20; B = 8'h97; #100;
A = 8'h20; B = 8'h98; #100;
A = 8'h20; B = 8'h99; #100;
A = 8'h20; B = 8'h9A; #100;
A = 8'h20; B = 8'h9B; #100;
A = 8'h20; B = 8'h9C; #100;
A = 8'h20; B = 8'h9D; #100;
A = 8'h20; B = 8'h9E; #100;
A = 8'h20; B = 8'h9F; #100;
A = 8'h20; B = 8'hA0; #100;
A = 8'h20; B = 8'hA1; #100;
A = 8'h20; B = 8'hA2; #100;
A = 8'h20; B = 8'hA3; #100;
A = 8'h20; B = 8'hA4; #100;
A = 8'h20; B = 8'hA5; #100;
A = 8'h20; B = 8'hA6; #100;
A = 8'h20; B = 8'hA7; #100;
A = 8'h20; B = 8'hA8; #100;
A = 8'h20; B = 8'hA9; #100;
A = 8'h20; B = 8'hAA; #100;
A = 8'h20; B = 8'hAB; #100;
A = 8'h20; B = 8'hAC; #100;
A = 8'h20; B = 8'hAD; #100;
A = 8'h20; B = 8'hAE; #100;
A = 8'h20; B = 8'hAF; #100;
A = 8'h20; B = 8'hB0; #100;
A = 8'h20; B = 8'hB1; #100;
A = 8'h20; B = 8'hB2; #100;
A = 8'h20; B = 8'hB3; #100;
A = 8'h20; B = 8'hB4; #100;
A = 8'h20; B = 8'hB5; #100;
A = 8'h20; B = 8'hB6; #100;
A = 8'h20; B = 8'hB7; #100;
A = 8'h20; B = 8'hB8; #100;
A = 8'h20; B = 8'hB9; #100;
A = 8'h20; B = 8'hBA; #100;
A = 8'h20; B = 8'hBB; #100;
A = 8'h20; B = 8'hBC; #100;
A = 8'h20; B = 8'hBD; #100;
A = 8'h20; B = 8'hBE; #100;
A = 8'h20; B = 8'hBF; #100;
A = 8'h20; B = 8'hC0; #100;
A = 8'h20; B = 8'hC1; #100;
A = 8'h20; B = 8'hC2; #100;
A = 8'h20; B = 8'hC3; #100;
A = 8'h20; B = 8'hC4; #100;
A = 8'h20; B = 8'hC5; #100;
A = 8'h20; B = 8'hC6; #100;
A = 8'h20; B = 8'hC7; #100;
A = 8'h20; B = 8'hC8; #100;
A = 8'h20; B = 8'hC9; #100;
A = 8'h20; B = 8'hCA; #100;
A = 8'h20; B = 8'hCB; #100;
A = 8'h20; B = 8'hCC; #100;
A = 8'h20; B = 8'hCD; #100;
A = 8'h20; B = 8'hCE; #100;
A = 8'h20; B = 8'hCF; #100;
A = 8'h20; B = 8'hD0; #100;
A = 8'h20; B = 8'hD1; #100;
A = 8'h20; B = 8'hD2; #100;
A = 8'h20; B = 8'hD3; #100;
A = 8'h20; B = 8'hD4; #100;
A = 8'h20; B = 8'hD5; #100;
A = 8'h20; B = 8'hD6; #100;
A = 8'h20; B = 8'hD7; #100;
A = 8'h20; B = 8'hD8; #100;
A = 8'h20; B = 8'hD9; #100;
A = 8'h20; B = 8'hDA; #100;
A = 8'h20; B = 8'hDB; #100;
A = 8'h20; B = 8'hDC; #100;
A = 8'h20; B = 8'hDD; #100;
A = 8'h20; B = 8'hDE; #100;
A = 8'h20; B = 8'hDF; #100;
A = 8'h20; B = 8'hE0; #100;
A = 8'h20; B = 8'hE1; #100;
A = 8'h20; B = 8'hE2; #100;
A = 8'h20; B = 8'hE3; #100;
A = 8'h20; B = 8'hE4; #100;
A = 8'h20; B = 8'hE5; #100;
A = 8'h20; B = 8'hE6; #100;
A = 8'h20; B = 8'hE7; #100;
A = 8'h20; B = 8'hE8; #100;
A = 8'h20; B = 8'hE9; #100;
A = 8'h20; B = 8'hEA; #100;
A = 8'h20; B = 8'hEB; #100;
A = 8'h20; B = 8'hEC; #100;
A = 8'h20; B = 8'hED; #100;
A = 8'h20; B = 8'hEE; #100;
A = 8'h20; B = 8'hEF; #100;
A = 8'h20; B = 8'hF0; #100;
A = 8'h20; B = 8'hF1; #100;
A = 8'h20; B = 8'hF2; #100;
A = 8'h20; B = 8'hF3; #100;
A = 8'h20; B = 8'hF4; #100;
A = 8'h20; B = 8'hF5; #100;
A = 8'h20; B = 8'hF6; #100;
A = 8'h20; B = 8'hF7; #100;
A = 8'h20; B = 8'hF8; #100;
A = 8'h20; B = 8'hF9; #100;
A = 8'h20; B = 8'hFA; #100;
A = 8'h20; B = 8'hFB; #100;
A = 8'h20; B = 8'hFC; #100;
A = 8'h20; B = 8'hFD; #100;
A = 8'h20; B = 8'hFE; #100;
A = 8'h20; B = 8'hFF; #100;
A = 8'h21; B = 8'h0; #100;
A = 8'h21; B = 8'h1; #100;
A = 8'h21; B = 8'h2; #100;
A = 8'h21; B = 8'h3; #100;
A = 8'h21; B = 8'h4; #100;
A = 8'h21; B = 8'h5; #100;
A = 8'h21; B = 8'h6; #100;
A = 8'h21; B = 8'h7; #100;
A = 8'h21; B = 8'h8; #100;
A = 8'h21; B = 8'h9; #100;
A = 8'h21; B = 8'hA; #100;
A = 8'h21; B = 8'hB; #100;
A = 8'h21; B = 8'hC; #100;
A = 8'h21; B = 8'hD; #100;
A = 8'h21; B = 8'hE; #100;
A = 8'h21; B = 8'hF; #100;
A = 8'h21; B = 8'h10; #100;
A = 8'h21; B = 8'h11; #100;
A = 8'h21; B = 8'h12; #100;
A = 8'h21; B = 8'h13; #100;
A = 8'h21; B = 8'h14; #100;
A = 8'h21; B = 8'h15; #100;
A = 8'h21; B = 8'h16; #100;
A = 8'h21; B = 8'h17; #100;
A = 8'h21; B = 8'h18; #100;
A = 8'h21; B = 8'h19; #100;
A = 8'h21; B = 8'h1A; #100;
A = 8'h21; B = 8'h1B; #100;
A = 8'h21; B = 8'h1C; #100;
A = 8'h21; B = 8'h1D; #100;
A = 8'h21; B = 8'h1E; #100;
A = 8'h21; B = 8'h1F; #100;
A = 8'h21; B = 8'h20; #100;
A = 8'h21; B = 8'h21; #100;
A = 8'h21; B = 8'h22; #100;
A = 8'h21; B = 8'h23; #100;
A = 8'h21; B = 8'h24; #100;
A = 8'h21; B = 8'h25; #100;
A = 8'h21; B = 8'h26; #100;
A = 8'h21; B = 8'h27; #100;
A = 8'h21; B = 8'h28; #100;
A = 8'h21; B = 8'h29; #100;
A = 8'h21; B = 8'h2A; #100;
A = 8'h21; B = 8'h2B; #100;
A = 8'h21; B = 8'h2C; #100;
A = 8'h21; B = 8'h2D; #100;
A = 8'h21; B = 8'h2E; #100;
A = 8'h21; B = 8'h2F; #100;
A = 8'h21; B = 8'h30; #100;
A = 8'h21; B = 8'h31; #100;
A = 8'h21; B = 8'h32; #100;
A = 8'h21; B = 8'h33; #100;
A = 8'h21; B = 8'h34; #100;
A = 8'h21; B = 8'h35; #100;
A = 8'h21; B = 8'h36; #100;
A = 8'h21; B = 8'h37; #100;
A = 8'h21; B = 8'h38; #100;
A = 8'h21; B = 8'h39; #100;
A = 8'h21; B = 8'h3A; #100;
A = 8'h21; B = 8'h3B; #100;
A = 8'h21; B = 8'h3C; #100;
A = 8'h21; B = 8'h3D; #100;
A = 8'h21; B = 8'h3E; #100;
A = 8'h21; B = 8'h3F; #100;
A = 8'h21; B = 8'h40; #100;
A = 8'h21; B = 8'h41; #100;
A = 8'h21; B = 8'h42; #100;
A = 8'h21; B = 8'h43; #100;
A = 8'h21; B = 8'h44; #100;
A = 8'h21; B = 8'h45; #100;
A = 8'h21; B = 8'h46; #100;
A = 8'h21; B = 8'h47; #100;
A = 8'h21; B = 8'h48; #100;
A = 8'h21; B = 8'h49; #100;
A = 8'h21; B = 8'h4A; #100;
A = 8'h21; B = 8'h4B; #100;
A = 8'h21; B = 8'h4C; #100;
A = 8'h21; B = 8'h4D; #100;
A = 8'h21; B = 8'h4E; #100;
A = 8'h21; B = 8'h4F; #100;
A = 8'h21; B = 8'h50; #100;
A = 8'h21; B = 8'h51; #100;
A = 8'h21; B = 8'h52; #100;
A = 8'h21; B = 8'h53; #100;
A = 8'h21; B = 8'h54; #100;
A = 8'h21; B = 8'h55; #100;
A = 8'h21; B = 8'h56; #100;
A = 8'h21; B = 8'h57; #100;
A = 8'h21; B = 8'h58; #100;
A = 8'h21; B = 8'h59; #100;
A = 8'h21; B = 8'h5A; #100;
A = 8'h21; B = 8'h5B; #100;
A = 8'h21; B = 8'h5C; #100;
A = 8'h21; B = 8'h5D; #100;
A = 8'h21; B = 8'h5E; #100;
A = 8'h21; B = 8'h5F; #100;
A = 8'h21; B = 8'h60; #100;
A = 8'h21; B = 8'h61; #100;
A = 8'h21; B = 8'h62; #100;
A = 8'h21; B = 8'h63; #100;
A = 8'h21; B = 8'h64; #100;
A = 8'h21; B = 8'h65; #100;
A = 8'h21; B = 8'h66; #100;
A = 8'h21; B = 8'h67; #100;
A = 8'h21; B = 8'h68; #100;
A = 8'h21; B = 8'h69; #100;
A = 8'h21; B = 8'h6A; #100;
A = 8'h21; B = 8'h6B; #100;
A = 8'h21; B = 8'h6C; #100;
A = 8'h21; B = 8'h6D; #100;
A = 8'h21; B = 8'h6E; #100;
A = 8'h21; B = 8'h6F; #100;
A = 8'h21; B = 8'h70; #100;
A = 8'h21; B = 8'h71; #100;
A = 8'h21; B = 8'h72; #100;
A = 8'h21; B = 8'h73; #100;
A = 8'h21; B = 8'h74; #100;
A = 8'h21; B = 8'h75; #100;
A = 8'h21; B = 8'h76; #100;
A = 8'h21; B = 8'h77; #100;
A = 8'h21; B = 8'h78; #100;
A = 8'h21; B = 8'h79; #100;
A = 8'h21; B = 8'h7A; #100;
A = 8'h21; B = 8'h7B; #100;
A = 8'h21; B = 8'h7C; #100;
A = 8'h21; B = 8'h7D; #100;
A = 8'h21; B = 8'h7E; #100;
A = 8'h21; B = 8'h7F; #100;
A = 8'h21; B = 8'h80; #100;
A = 8'h21; B = 8'h81; #100;
A = 8'h21; B = 8'h82; #100;
A = 8'h21; B = 8'h83; #100;
A = 8'h21; B = 8'h84; #100;
A = 8'h21; B = 8'h85; #100;
A = 8'h21; B = 8'h86; #100;
A = 8'h21; B = 8'h87; #100;
A = 8'h21; B = 8'h88; #100;
A = 8'h21; B = 8'h89; #100;
A = 8'h21; B = 8'h8A; #100;
A = 8'h21; B = 8'h8B; #100;
A = 8'h21; B = 8'h8C; #100;
A = 8'h21; B = 8'h8D; #100;
A = 8'h21; B = 8'h8E; #100;
A = 8'h21; B = 8'h8F; #100;
A = 8'h21; B = 8'h90; #100;
A = 8'h21; B = 8'h91; #100;
A = 8'h21; B = 8'h92; #100;
A = 8'h21; B = 8'h93; #100;
A = 8'h21; B = 8'h94; #100;
A = 8'h21; B = 8'h95; #100;
A = 8'h21; B = 8'h96; #100;
A = 8'h21; B = 8'h97; #100;
A = 8'h21; B = 8'h98; #100;
A = 8'h21; B = 8'h99; #100;
A = 8'h21; B = 8'h9A; #100;
A = 8'h21; B = 8'h9B; #100;
A = 8'h21; B = 8'h9C; #100;
A = 8'h21; B = 8'h9D; #100;
A = 8'h21; B = 8'h9E; #100;
A = 8'h21; B = 8'h9F; #100;
A = 8'h21; B = 8'hA0; #100;
A = 8'h21; B = 8'hA1; #100;
A = 8'h21; B = 8'hA2; #100;
A = 8'h21; B = 8'hA3; #100;
A = 8'h21; B = 8'hA4; #100;
A = 8'h21; B = 8'hA5; #100;
A = 8'h21; B = 8'hA6; #100;
A = 8'h21; B = 8'hA7; #100;
A = 8'h21; B = 8'hA8; #100;
A = 8'h21; B = 8'hA9; #100;
A = 8'h21; B = 8'hAA; #100;
A = 8'h21; B = 8'hAB; #100;
A = 8'h21; B = 8'hAC; #100;
A = 8'h21; B = 8'hAD; #100;
A = 8'h21; B = 8'hAE; #100;
A = 8'h21; B = 8'hAF; #100;
A = 8'h21; B = 8'hB0; #100;
A = 8'h21; B = 8'hB1; #100;
A = 8'h21; B = 8'hB2; #100;
A = 8'h21; B = 8'hB3; #100;
A = 8'h21; B = 8'hB4; #100;
A = 8'h21; B = 8'hB5; #100;
A = 8'h21; B = 8'hB6; #100;
A = 8'h21; B = 8'hB7; #100;
A = 8'h21; B = 8'hB8; #100;
A = 8'h21; B = 8'hB9; #100;
A = 8'h21; B = 8'hBA; #100;
A = 8'h21; B = 8'hBB; #100;
A = 8'h21; B = 8'hBC; #100;
A = 8'h21; B = 8'hBD; #100;
A = 8'h21; B = 8'hBE; #100;
A = 8'h21; B = 8'hBF; #100;
A = 8'h21; B = 8'hC0; #100;
A = 8'h21; B = 8'hC1; #100;
A = 8'h21; B = 8'hC2; #100;
A = 8'h21; B = 8'hC3; #100;
A = 8'h21; B = 8'hC4; #100;
A = 8'h21; B = 8'hC5; #100;
A = 8'h21; B = 8'hC6; #100;
A = 8'h21; B = 8'hC7; #100;
A = 8'h21; B = 8'hC8; #100;
A = 8'h21; B = 8'hC9; #100;
A = 8'h21; B = 8'hCA; #100;
A = 8'h21; B = 8'hCB; #100;
A = 8'h21; B = 8'hCC; #100;
A = 8'h21; B = 8'hCD; #100;
A = 8'h21; B = 8'hCE; #100;
A = 8'h21; B = 8'hCF; #100;
A = 8'h21; B = 8'hD0; #100;
A = 8'h21; B = 8'hD1; #100;
A = 8'h21; B = 8'hD2; #100;
A = 8'h21; B = 8'hD3; #100;
A = 8'h21; B = 8'hD4; #100;
A = 8'h21; B = 8'hD5; #100;
A = 8'h21; B = 8'hD6; #100;
A = 8'h21; B = 8'hD7; #100;
A = 8'h21; B = 8'hD8; #100;
A = 8'h21; B = 8'hD9; #100;
A = 8'h21; B = 8'hDA; #100;
A = 8'h21; B = 8'hDB; #100;
A = 8'h21; B = 8'hDC; #100;
A = 8'h21; B = 8'hDD; #100;
A = 8'h21; B = 8'hDE; #100;
A = 8'h21; B = 8'hDF; #100;
A = 8'h21; B = 8'hE0; #100;
A = 8'h21; B = 8'hE1; #100;
A = 8'h21; B = 8'hE2; #100;
A = 8'h21; B = 8'hE3; #100;
A = 8'h21; B = 8'hE4; #100;
A = 8'h21; B = 8'hE5; #100;
A = 8'h21; B = 8'hE6; #100;
A = 8'h21; B = 8'hE7; #100;
A = 8'h21; B = 8'hE8; #100;
A = 8'h21; B = 8'hE9; #100;
A = 8'h21; B = 8'hEA; #100;
A = 8'h21; B = 8'hEB; #100;
A = 8'h21; B = 8'hEC; #100;
A = 8'h21; B = 8'hED; #100;
A = 8'h21; B = 8'hEE; #100;
A = 8'h21; B = 8'hEF; #100;
A = 8'h21; B = 8'hF0; #100;
A = 8'h21; B = 8'hF1; #100;
A = 8'h21; B = 8'hF2; #100;
A = 8'h21; B = 8'hF3; #100;
A = 8'h21; B = 8'hF4; #100;
A = 8'h21; B = 8'hF5; #100;
A = 8'h21; B = 8'hF6; #100;
A = 8'h21; B = 8'hF7; #100;
A = 8'h21; B = 8'hF8; #100;
A = 8'h21; B = 8'hF9; #100;
A = 8'h21; B = 8'hFA; #100;
A = 8'h21; B = 8'hFB; #100;
A = 8'h21; B = 8'hFC; #100;
A = 8'h21; B = 8'hFD; #100;
A = 8'h21; B = 8'hFE; #100;
A = 8'h21; B = 8'hFF; #100;
A = 8'h22; B = 8'h0; #100;
A = 8'h22; B = 8'h1; #100;
A = 8'h22; B = 8'h2; #100;
A = 8'h22; B = 8'h3; #100;
A = 8'h22; B = 8'h4; #100;
A = 8'h22; B = 8'h5; #100;
A = 8'h22; B = 8'h6; #100;
A = 8'h22; B = 8'h7; #100;
A = 8'h22; B = 8'h8; #100;
A = 8'h22; B = 8'h9; #100;
A = 8'h22; B = 8'hA; #100;
A = 8'h22; B = 8'hB; #100;
A = 8'h22; B = 8'hC; #100;
A = 8'h22; B = 8'hD; #100;
A = 8'h22; B = 8'hE; #100;
A = 8'h22; B = 8'hF; #100;
A = 8'h22; B = 8'h10; #100;
A = 8'h22; B = 8'h11; #100;
A = 8'h22; B = 8'h12; #100;
A = 8'h22; B = 8'h13; #100;
A = 8'h22; B = 8'h14; #100;
A = 8'h22; B = 8'h15; #100;
A = 8'h22; B = 8'h16; #100;
A = 8'h22; B = 8'h17; #100;
A = 8'h22; B = 8'h18; #100;
A = 8'h22; B = 8'h19; #100;
A = 8'h22; B = 8'h1A; #100;
A = 8'h22; B = 8'h1B; #100;
A = 8'h22; B = 8'h1C; #100;
A = 8'h22; B = 8'h1D; #100;
A = 8'h22; B = 8'h1E; #100;
A = 8'h22; B = 8'h1F; #100;
A = 8'h22; B = 8'h20; #100;
A = 8'h22; B = 8'h21; #100;
A = 8'h22; B = 8'h22; #100;
A = 8'h22; B = 8'h23; #100;
A = 8'h22; B = 8'h24; #100;
A = 8'h22; B = 8'h25; #100;
A = 8'h22; B = 8'h26; #100;
A = 8'h22; B = 8'h27; #100;
A = 8'h22; B = 8'h28; #100;
A = 8'h22; B = 8'h29; #100;
A = 8'h22; B = 8'h2A; #100;
A = 8'h22; B = 8'h2B; #100;
A = 8'h22; B = 8'h2C; #100;
A = 8'h22; B = 8'h2D; #100;
A = 8'h22; B = 8'h2E; #100;
A = 8'h22; B = 8'h2F; #100;
A = 8'h22; B = 8'h30; #100;
A = 8'h22; B = 8'h31; #100;
A = 8'h22; B = 8'h32; #100;
A = 8'h22; B = 8'h33; #100;
A = 8'h22; B = 8'h34; #100;
A = 8'h22; B = 8'h35; #100;
A = 8'h22; B = 8'h36; #100;
A = 8'h22; B = 8'h37; #100;
A = 8'h22; B = 8'h38; #100;
A = 8'h22; B = 8'h39; #100;
A = 8'h22; B = 8'h3A; #100;
A = 8'h22; B = 8'h3B; #100;
A = 8'h22; B = 8'h3C; #100;
A = 8'h22; B = 8'h3D; #100;
A = 8'h22; B = 8'h3E; #100;
A = 8'h22; B = 8'h3F; #100;
A = 8'h22; B = 8'h40; #100;
A = 8'h22; B = 8'h41; #100;
A = 8'h22; B = 8'h42; #100;
A = 8'h22; B = 8'h43; #100;
A = 8'h22; B = 8'h44; #100;
A = 8'h22; B = 8'h45; #100;
A = 8'h22; B = 8'h46; #100;
A = 8'h22; B = 8'h47; #100;
A = 8'h22; B = 8'h48; #100;
A = 8'h22; B = 8'h49; #100;
A = 8'h22; B = 8'h4A; #100;
A = 8'h22; B = 8'h4B; #100;
A = 8'h22; B = 8'h4C; #100;
A = 8'h22; B = 8'h4D; #100;
A = 8'h22; B = 8'h4E; #100;
A = 8'h22; B = 8'h4F; #100;
A = 8'h22; B = 8'h50; #100;
A = 8'h22; B = 8'h51; #100;
A = 8'h22; B = 8'h52; #100;
A = 8'h22; B = 8'h53; #100;
A = 8'h22; B = 8'h54; #100;
A = 8'h22; B = 8'h55; #100;
A = 8'h22; B = 8'h56; #100;
A = 8'h22; B = 8'h57; #100;
A = 8'h22; B = 8'h58; #100;
A = 8'h22; B = 8'h59; #100;
A = 8'h22; B = 8'h5A; #100;
A = 8'h22; B = 8'h5B; #100;
A = 8'h22; B = 8'h5C; #100;
A = 8'h22; B = 8'h5D; #100;
A = 8'h22; B = 8'h5E; #100;
A = 8'h22; B = 8'h5F; #100;
A = 8'h22; B = 8'h60; #100;
A = 8'h22; B = 8'h61; #100;
A = 8'h22; B = 8'h62; #100;
A = 8'h22; B = 8'h63; #100;
A = 8'h22; B = 8'h64; #100;
A = 8'h22; B = 8'h65; #100;
A = 8'h22; B = 8'h66; #100;
A = 8'h22; B = 8'h67; #100;
A = 8'h22; B = 8'h68; #100;
A = 8'h22; B = 8'h69; #100;
A = 8'h22; B = 8'h6A; #100;
A = 8'h22; B = 8'h6B; #100;
A = 8'h22; B = 8'h6C; #100;
A = 8'h22; B = 8'h6D; #100;
A = 8'h22; B = 8'h6E; #100;
A = 8'h22; B = 8'h6F; #100;
A = 8'h22; B = 8'h70; #100;
A = 8'h22; B = 8'h71; #100;
A = 8'h22; B = 8'h72; #100;
A = 8'h22; B = 8'h73; #100;
A = 8'h22; B = 8'h74; #100;
A = 8'h22; B = 8'h75; #100;
A = 8'h22; B = 8'h76; #100;
A = 8'h22; B = 8'h77; #100;
A = 8'h22; B = 8'h78; #100;
A = 8'h22; B = 8'h79; #100;
A = 8'h22; B = 8'h7A; #100;
A = 8'h22; B = 8'h7B; #100;
A = 8'h22; B = 8'h7C; #100;
A = 8'h22; B = 8'h7D; #100;
A = 8'h22; B = 8'h7E; #100;
A = 8'h22; B = 8'h7F; #100;
A = 8'h22; B = 8'h80; #100;
A = 8'h22; B = 8'h81; #100;
A = 8'h22; B = 8'h82; #100;
A = 8'h22; B = 8'h83; #100;
A = 8'h22; B = 8'h84; #100;
A = 8'h22; B = 8'h85; #100;
A = 8'h22; B = 8'h86; #100;
A = 8'h22; B = 8'h87; #100;
A = 8'h22; B = 8'h88; #100;
A = 8'h22; B = 8'h89; #100;
A = 8'h22; B = 8'h8A; #100;
A = 8'h22; B = 8'h8B; #100;
A = 8'h22; B = 8'h8C; #100;
A = 8'h22; B = 8'h8D; #100;
A = 8'h22; B = 8'h8E; #100;
A = 8'h22; B = 8'h8F; #100;
A = 8'h22; B = 8'h90; #100;
A = 8'h22; B = 8'h91; #100;
A = 8'h22; B = 8'h92; #100;
A = 8'h22; B = 8'h93; #100;
A = 8'h22; B = 8'h94; #100;
A = 8'h22; B = 8'h95; #100;
A = 8'h22; B = 8'h96; #100;
A = 8'h22; B = 8'h97; #100;
A = 8'h22; B = 8'h98; #100;
A = 8'h22; B = 8'h99; #100;
A = 8'h22; B = 8'h9A; #100;
A = 8'h22; B = 8'h9B; #100;
A = 8'h22; B = 8'h9C; #100;
A = 8'h22; B = 8'h9D; #100;
A = 8'h22; B = 8'h9E; #100;
A = 8'h22; B = 8'h9F; #100;
A = 8'h22; B = 8'hA0; #100;
A = 8'h22; B = 8'hA1; #100;
A = 8'h22; B = 8'hA2; #100;
A = 8'h22; B = 8'hA3; #100;
A = 8'h22; B = 8'hA4; #100;
A = 8'h22; B = 8'hA5; #100;
A = 8'h22; B = 8'hA6; #100;
A = 8'h22; B = 8'hA7; #100;
A = 8'h22; B = 8'hA8; #100;
A = 8'h22; B = 8'hA9; #100;
A = 8'h22; B = 8'hAA; #100;
A = 8'h22; B = 8'hAB; #100;
A = 8'h22; B = 8'hAC; #100;
A = 8'h22; B = 8'hAD; #100;
A = 8'h22; B = 8'hAE; #100;
A = 8'h22; B = 8'hAF; #100;
A = 8'h22; B = 8'hB0; #100;
A = 8'h22; B = 8'hB1; #100;
A = 8'h22; B = 8'hB2; #100;
A = 8'h22; B = 8'hB3; #100;
A = 8'h22; B = 8'hB4; #100;
A = 8'h22; B = 8'hB5; #100;
A = 8'h22; B = 8'hB6; #100;
A = 8'h22; B = 8'hB7; #100;
A = 8'h22; B = 8'hB8; #100;
A = 8'h22; B = 8'hB9; #100;
A = 8'h22; B = 8'hBA; #100;
A = 8'h22; B = 8'hBB; #100;
A = 8'h22; B = 8'hBC; #100;
A = 8'h22; B = 8'hBD; #100;
A = 8'h22; B = 8'hBE; #100;
A = 8'h22; B = 8'hBF; #100;
A = 8'h22; B = 8'hC0; #100;
A = 8'h22; B = 8'hC1; #100;
A = 8'h22; B = 8'hC2; #100;
A = 8'h22; B = 8'hC3; #100;
A = 8'h22; B = 8'hC4; #100;
A = 8'h22; B = 8'hC5; #100;
A = 8'h22; B = 8'hC6; #100;
A = 8'h22; B = 8'hC7; #100;
A = 8'h22; B = 8'hC8; #100;
A = 8'h22; B = 8'hC9; #100;
A = 8'h22; B = 8'hCA; #100;
A = 8'h22; B = 8'hCB; #100;
A = 8'h22; B = 8'hCC; #100;
A = 8'h22; B = 8'hCD; #100;
A = 8'h22; B = 8'hCE; #100;
A = 8'h22; B = 8'hCF; #100;
A = 8'h22; B = 8'hD0; #100;
A = 8'h22; B = 8'hD1; #100;
A = 8'h22; B = 8'hD2; #100;
A = 8'h22; B = 8'hD3; #100;
A = 8'h22; B = 8'hD4; #100;
A = 8'h22; B = 8'hD5; #100;
A = 8'h22; B = 8'hD6; #100;
A = 8'h22; B = 8'hD7; #100;
A = 8'h22; B = 8'hD8; #100;
A = 8'h22; B = 8'hD9; #100;
A = 8'h22; B = 8'hDA; #100;
A = 8'h22; B = 8'hDB; #100;
A = 8'h22; B = 8'hDC; #100;
A = 8'h22; B = 8'hDD; #100;
A = 8'h22; B = 8'hDE; #100;
A = 8'h22; B = 8'hDF; #100;
A = 8'h22; B = 8'hE0; #100;
A = 8'h22; B = 8'hE1; #100;
A = 8'h22; B = 8'hE2; #100;
A = 8'h22; B = 8'hE3; #100;
A = 8'h22; B = 8'hE4; #100;
A = 8'h22; B = 8'hE5; #100;
A = 8'h22; B = 8'hE6; #100;
A = 8'h22; B = 8'hE7; #100;
A = 8'h22; B = 8'hE8; #100;
A = 8'h22; B = 8'hE9; #100;
A = 8'h22; B = 8'hEA; #100;
A = 8'h22; B = 8'hEB; #100;
A = 8'h22; B = 8'hEC; #100;
A = 8'h22; B = 8'hED; #100;
A = 8'h22; B = 8'hEE; #100;
A = 8'h22; B = 8'hEF; #100;
A = 8'h22; B = 8'hF0; #100;
A = 8'h22; B = 8'hF1; #100;
A = 8'h22; B = 8'hF2; #100;
A = 8'h22; B = 8'hF3; #100;
A = 8'h22; B = 8'hF4; #100;
A = 8'h22; B = 8'hF5; #100;
A = 8'h22; B = 8'hF6; #100;
A = 8'h22; B = 8'hF7; #100;
A = 8'h22; B = 8'hF8; #100;
A = 8'h22; B = 8'hF9; #100;
A = 8'h22; B = 8'hFA; #100;
A = 8'h22; B = 8'hFB; #100;
A = 8'h22; B = 8'hFC; #100;
A = 8'h22; B = 8'hFD; #100;
A = 8'h22; B = 8'hFE; #100;
A = 8'h22; B = 8'hFF; #100;
A = 8'h23; B = 8'h0; #100;
A = 8'h23; B = 8'h1; #100;
A = 8'h23; B = 8'h2; #100;
A = 8'h23; B = 8'h3; #100;
A = 8'h23; B = 8'h4; #100;
A = 8'h23; B = 8'h5; #100;
A = 8'h23; B = 8'h6; #100;
A = 8'h23; B = 8'h7; #100;
A = 8'h23; B = 8'h8; #100;
A = 8'h23; B = 8'h9; #100;
A = 8'h23; B = 8'hA; #100;
A = 8'h23; B = 8'hB; #100;
A = 8'h23; B = 8'hC; #100;
A = 8'h23; B = 8'hD; #100;
A = 8'h23; B = 8'hE; #100;
A = 8'h23; B = 8'hF; #100;
A = 8'h23; B = 8'h10; #100;
A = 8'h23; B = 8'h11; #100;
A = 8'h23; B = 8'h12; #100;
A = 8'h23; B = 8'h13; #100;
A = 8'h23; B = 8'h14; #100;
A = 8'h23; B = 8'h15; #100;
A = 8'h23; B = 8'h16; #100;
A = 8'h23; B = 8'h17; #100;
A = 8'h23; B = 8'h18; #100;
A = 8'h23; B = 8'h19; #100;
A = 8'h23; B = 8'h1A; #100;
A = 8'h23; B = 8'h1B; #100;
A = 8'h23; B = 8'h1C; #100;
A = 8'h23; B = 8'h1D; #100;
A = 8'h23; B = 8'h1E; #100;
A = 8'h23; B = 8'h1F; #100;
A = 8'h23; B = 8'h20; #100;
A = 8'h23; B = 8'h21; #100;
A = 8'h23; B = 8'h22; #100;
A = 8'h23; B = 8'h23; #100;
A = 8'h23; B = 8'h24; #100;
A = 8'h23; B = 8'h25; #100;
A = 8'h23; B = 8'h26; #100;
A = 8'h23; B = 8'h27; #100;
A = 8'h23; B = 8'h28; #100;
A = 8'h23; B = 8'h29; #100;
A = 8'h23; B = 8'h2A; #100;
A = 8'h23; B = 8'h2B; #100;
A = 8'h23; B = 8'h2C; #100;
A = 8'h23; B = 8'h2D; #100;
A = 8'h23; B = 8'h2E; #100;
A = 8'h23; B = 8'h2F; #100;
A = 8'h23; B = 8'h30; #100;
A = 8'h23; B = 8'h31; #100;
A = 8'h23; B = 8'h32; #100;
A = 8'h23; B = 8'h33; #100;
A = 8'h23; B = 8'h34; #100;
A = 8'h23; B = 8'h35; #100;
A = 8'h23; B = 8'h36; #100;
A = 8'h23; B = 8'h37; #100;
A = 8'h23; B = 8'h38; #100;
A = 8'h23; B = 8'h39; #100;
A = 8'h23; B = 8'h3A; #100;
A = 8'h23; B = 8'h3B; #100;
A = 8'h23; B = 8'h3C; #100;
A = 8'h23; B = 8'h3D; #100;
A = 8'h23; B = 8'h3E; #100;
A = 8'h23; B = 8'h3F; #100;
A = 8'h23; B = 8'h40; #100;
A = 8'h23; B = 8'h41; #100;
A = 8'h23; B = 8'h42; #100;
A = 8'h23; B = 8'h43; #100;
A = 8'h23; B = 8'h44; #100;
A = 8'h23; B = 8'h45; #100;
A = 8'h23; B = 8'h46; #100;
A = 8'h23; B = 8'h47; #100;
A = 8'h23; B = 8'h48; #100;
A = 8'h23; B = 8'h49; #100;
A = 8'h23; B = 8'h4A; #100;
A = 8'h23; B = 8'h4B; #100;
A = 8'h23; B = 8'h4C; #100;
A = 8'h23; B = 8'h4D; #100;
A = 8'h23; B = 8'h4E; #100;
A = 8'h23; B = 8'h4F; #100;
A = 8'h23; B = 8'h50; #100;
A = 8'h23; B = 8'h51; #100;
A = 8'h23; B = 8'h52; #100;
A = 8'h23; B = 8'h53; #100;
A = 8'h23; B = 8'h54; #100;
A = 8'h23; B = 8'h55; #100;
A = 8'h23; B = 8'h56; #100;
A = 8'h23; B = 8'h57; #100;
A = 8'h23; B = 8'h58; #100;
A = 8'h23; B = 8'h59; #100;
A = 8'h23; B = 8'h5A; #100;
A = 8'h23; B = 8'h5B; #100;
A = 8'h23; B = 8'h5C; #100;
A = 8'h23; B = 8'h5D; #100;
A = 8'h23; B = 8'h5E; #100;
A = 8'h23; B = 8'h5F; #100;
A = 8'h23; B = 8'h60; #100;
A = 8'h23; B = 8'h61; #100;
A = 8'h23; B = 8'h62; #100;
A = 8'h23; B = 8'h63; #100;
A = 8'h23; B = 8'h64; #100;
A = 8'h23; B = 8'h65; #100;
A = 8'h23; B = 8'h66; #100;
A = 8'h23; B = 8'h67; #100;
A = 8'h23; B = 8'h68; #100;
A = 8'h23; B = 8'h69; #100;
A = 8'h23; B = 8'h6A; #100;
A = 8'h23; B = 8'h6B; #100;
A = 8'h23; B = 8'h6C; #100;
A = 8'h23; B = 8'h6D; #100;
A = 8'h23; B = 8'h6E; #100;
A = 8'h23; B = 8'h6F; #100;
A = 8'h23; B = 8'h70; #100;
A = 8'h23; B = 8'h71; #100;
A = 8'h23; B = 8'h72; #100;
A = 8'h23; B = 8'h73; #100;
A = 8'h23; B = 8'h74; #100;
A = 8'h23; B = 8'h75; #100;
A = 8'h23; B = 8'h76; #100;
A = 8'h23; B = 8'h77; #100;
A = 8'h23; B = 8'h78; #100;
A = 8'h23; B = 8'h79; #100;
A = 8'h23; B = 8'h7A; #100;
A = 8'h23; B = 8'h7B; #100;
A = 8'h23; B = 8'h7C; #100;
A = 8'h23; B = 8'h7D; #100;
A = 8'h23; B = 8'h7E; #100;
A = 8'h23; B = 8'h7F; #100;
A = 8'h23; B = 8'h80; #100;
A = 8'h23; B = 8'h81; #100;
A = 8'h23; B = 8'h82; #100;
A = 8'h23; B = 8'h83; #100;
A = 8'h23; B = 8'h84; #100;
A = 8'h23; B = 8'h85; #100;
A = 8'h23; B = 8'h86; #100;
A = 8'h23; B = 8'h87; #100;
A = 8'h23; B = 8'h88; #100;
A = 8'h23; B = 8'h89; #100;
A = 8'h23; B = 8'h8A; #100;
A = 8'h23; B = 8'h8B; #100;
A = 8'h23; B = 8'h8C; #100;
A = 8'h23; B = 8'h8D; #100;
A = 8'h23; B = 8'h8E; #100;
A = 8'h23; B = 8'h8F; #100;
A = 8'h23; B = 8'h90; #100;
A = 8'h23; B = 8'h91; #100;
A = 8'h23; B = 8'h92; #100;
A = 8'h23; B = 8'h93; #100;
A = 8'h23; B = 8'h94; #100;
A = 8'h23; B = 8'h95; #100;
A = 8'h23; B = 8'h96; #100;
A = 8'h23; B = 8'h97; #100;
A = 8'h23; B = 8'h98; #100;
A = 8'h23; B = 8'h99; #100;
A = 8'h23; B = 8'h9A; #100;
A = 8'h23; B = 8'h9B; #100;
A = 8'h23; B = 8'h9C; #100;
A = 8'h23; B = 8'h9D; #100;
A = 8'h23; B = 8'h9E; #100;
A = 8'h23; B = 8'h9F; #100;
A = 8'h23; B = 8'hA0; #100;
A = 8'h23; B = 8'hA1; #100;
A = 8'h23; B = 8'hA2; #100;
A = 8'h23; B = 8'hA3; #100;
A = 8'h23; B = 8'hA4; #100;
A = 8'h23; B = 8'hA5; #100;
A = 8'h23; B = 8'hA6; #100;
A = 8'h23; B = 8'hA7; #100;
A = 8'h23; B = 8'hA8; #100;
A = 8'h23; B = 8'hA9; #100;
A = 8'h23; B = 8'hAA; #100;
A = 8'h23; B = 8'hAB; #100;
A = 8'h23; B = 8'hAC; #100;
A = 8'h23; B = 8'hAD; #100;
A = 8'h23; B = 8'hAE; #100;
A = 8'h23; B = 8'hAF; #100;
A = 8'h23; B = 8'hB0; #100;
A = 8'h23; B = 8'hB1; #100;
A = 8'h23; B = 8'hB2; #100;
A = 8'h23; B = 8'hB3; #100;
A = 8'h23; B = 8'hB4; #100;
A = 8'h23; B = 8'hB5; #100;
A = 8'h23; B = 8'hB6; #100;
A = 8'h23; B = 8'hB7; #100;
A = 8'h23; B = 8'hB8; #100;
A = 8'h23; B = 8'hB9; #100;
A = 8'h23; B = 8'hBA; #100;
A = 8'h23; B = 8'hBB; #100;
A = 8'h23; B = 8'hBC; #100;
A = 8'h23; B = 8'hBD; #100;
A = 8'h23; B = 8'hBE; #100;
A = 8'h23; B = 8'hBF; #100;
A = 8'h23; B = 8'hC0; #100;
A = 8'h23; B = 8'hC1; #100;
A = 8'h23; B = 8'hC2; #100;
A = 8'h23; B = 8'hC3; #100;
A = 8'h23; B = 8'hC4; #100;
A = 8'h23; B = 8'hC5; #100;
A = 8'h23; B = 8'hC6; #100;
A = 8'h23; B = 8'hC7; #100;
A = 8'h23; B = 8'hC8; #100;
A = 8'h23; B = 8'hC9; #100;
A = 8'h23; B = 8'hCA; #100;
A = 8'h23; B = 8'hCB; #100;
A = 8'h23; B = 8'hCC; #100;
A = 8'h23; B = 8'hCD; #100;
A = 8'h23; B = 8'hCE; #100;
A = 8'h23; B = 8'hCF; #100;
A = 8'h23; B = 8'hD0; #100;
A = 8'h23; B = 8'hD1; #100;
A = 8'h23; B = 8'hD2; #100;
A = 8'h23; B = 8'hD3; #100;
A = 8'h23; B = 8'hD4; #100;
A = 8'h23; B = 8'hD5; #100;
A = 8'h23; B = 8'hD6; #100;
A = 8'h23; B = 8'hD7; #100;
A = 8'h23; B = 8'hD8; #100;
A = 8'h23; B = 8'hD9; #100;
A = 8'h23; B = 8'hDA; #100;
A = 8'h23; B = 8'hDB; #100;
A = 8'h23; B = 8'hDC; #100;
A = 8'h23; B = 8'hDD; #100;
A = 8'h23; B = 8'hDE; #100;
A = 8'h23; B = 8'hDF; #100;
A = 8'h23; B = 8'hE0; #100;
A = 8'h23; B = 8'hE1; #100;
A = 8'h23; B = 8'hE2; #100;
A = 8'h23; B = 8'hE3; #100;
A = 8'h23; B = 8'hE4; #100;
A = 8'h23; B = 8'hE5; #100;
A = 8'h23; B = 8'hE6; #100;
A = 8'h23; B = 8'hE7; #100;
A = 8'h23; B = 8'hE8; #100;
A = 8'h23; B = 8'hE9; #100;
A = 8'h23; B = 8'hEA; #100;
A = 8'h23; B = 8'hEB; #100;
A = 8'h23; B = 8'hEC; #100;
A = 8'h23; B = 8'hED; #100;
A = 8'h23; B = 8'hEE; #100;
A = 8'h23; B = 8'hEF; #100;
A = 8'h23; B = 8'hF0; #100;
A = 8'h23; B = 8'hF1; #100;
A = 8'h23; B = 8'hF2; #100;
A = 8'h23; B = 8'hF3; #100;
A = 8'h23; B = 8'hF4; #100;
A = 8'h23; B = 8'hF5; #100;
A = 8'h23; B = 8'hF6; #100;
A = 8'h23; B = 8'hF7; #100;
A = 8'h23; B = 8'hF8; #100;
A = 8'h23; B = 8'hF9; #100;
A = 8'h23; B = 8'hFA; #100;
A = 8'h23; B = 8'hFB; #100;
A = 8'h23; B = 8'hFC; #100;
A = 8'h23; B = 8'hFD; #100;
A = 8'h23; B = 8'hFE; #100;
A = 8'h23; B = 8'hFF; #100;
A = 8'h24; B = 8'h0; #100;
A = 8'h24; B = 8'h1; #100;
A = 8'h24; B = 8'h2; #100;
A = 8'h24; B = 8'h3; #100;
A = 8'h24; B = 8'h4; #100;
A = 8'h24; B = 8'h5; #100;
A = 8'h24; B = 8'h6; #100;
A = 8'h24; B = 8'h7; #100;
A = 8'h24; B = 8'h8; #100;
A = 8'h24; B = 8'h9; #100;
A = 8'h24; B = 8'hA; #100;
A = 8'h24; B = 8'hB; #100;
A = 8'h24; B = 8'hC; #100;
A = 8'h24; B = 8'hD; #100;
A = 8'h24; B = 8'hE; #100;
A = 8'h24; B = 8'hF; #100;
A = 8'h24; B = 8'h10; #100;
A = 8'h24; B = 8'h11; #100;
A = 8'h24; B = 8'h12; #100;
A = 8'h24; B = 8'h13; #100;
A = 8'h24; B = 8'h14; #100;
A = 8'h24; B = 8'h15; #100;
A = 8'h24; B = 8'h16; #100;
A = 8'h24; B = 8'h17; #100;
A = 8'h24; B = 8'h18; #100;
A = 8'h24; B = 8'h19; #100;
A = 8'h24; B = 8'h1A; #100;
A = 8'h24; B = 8'h1B; #100;
A = 8'h24; B = 8'h1C; #100;
A = 8'h24; B = 8'h1D; #100;
A = 8'h24; B = 8'h1E; #100;
A = 8'h24; B = 8'h1F; #100;
A = 8'h24; B = 8'h20; #100;
A = 8'h24; B = 8'h21; #100;
A = 8'h24; B = 8'h22; #100;
A = 8'h24; B = 8'h23; #100;
A = 8'h24; B = 8'h24; #100;
A = 8'h24; B = 8'h25; #100;
A = 8'h24; B = 8'h26; #100;
A = 8'h24; B = 8'h27; #100;
A = 8'h24; B = 8'h28; #100;
A = 8'h24; B = 8'h29; #100;
A = 8'h24; B = 8'h2A; #100;
A = 8'h24; B = 8'h2B; #100;
A = 8'h24; B = 8'h2C; #100;
A = 8'h24; B = 8'h2D; #100;
A = 8'h24; B = 8'h2E; #100;
A = 8'h24; B = 8'h2F; #100;
A = 8'h24; B = 8'h30; #100;
A = 8'h24; B = 8'h31; #100;
A = 8'h24; B = 8'h32; #100;
A = 8'h24; B = 8'h33; #100;
A = 8'h24; B = 8'h34; #100;
A = 8'h24; B = 8'h35; #100;
A = 8'h24; B = 8'h36; #100;
A = 8'h24; B = 8'h37; #100;
A = 8'h24; B = 8'h38; #100;
A = 8'h24; B = 8'h39; #100;
A = 8'h24; B = 8'h3A; #100;
A = 8'h24; B = 8'h3B; #100;
A = 8'h24; B = 8'h3C; #100;
A = 8'h24; B = 8'h3D; #100;
A = 8'h24; B = 8'h3E; #100;
A = 8'h24; B = 8'h3F; #100;
A = 8'h24; B = 8'h40; #100;
A = 8'h24; B = 8'h41; #100;
A = 8'h24; B = 8'h42; #100;
A = 8'h24; B = 8'h43; #100;
A = 8'h24; B = 8'h44; #100;
A = 8'h24; B = 8'h45; #100;
A = 8'h24; B = 8'h46; #100;
A = 8'h24; B = 8'h47; #100;
A = 8'h24; B = 8'h48; #100;
A = 8'h24; B = 8'h49; #100;
A = 8'h24; B = 8'h4A; #100;
A = 8'h24; B = 8'h4B; #100;
A = 8'h24; B = 8'h4C; #100;
A = 8'h24; B = 8'h4D; #100;
A = 8'h24; B = 8'h4E; #100;
A = 8'h24; B = 8'h4F; #100;
A = 8'h24; B = 8'h50; #100;
A = 8'h24; B = 8'h51; #100;
A = 8'h24; B = 8'h52; #100;
A = 8'h24; B = 8'h53; #100;
A = 8'h24; B = 8'h54; #100;
A = 8'h24; B = 8'h55; #100;
A = 8'h24; B = 8'h56; #100;
A = 8'h24; B = 8'h57; #100;
A = 8'h24; B = 8'h58; #100;
A = 8'h24; B = 8'h59; #100;
A = 8'h24; B = 8'h5A; #100;
A = 8'h24; B = 8'h5B; #100;
A = 8'h24; B = 8'h5C; #100;
A = 8'h24; B = 8'h5D; #100;
A = 8'h24; B = 8'h5E; #100;
A = 8'h24; B = 8'h5F; #100;
A = 8'h24; B = 8'h60; #100;
A = 8'h24; B = 8'h61; #100;
A = 8'h24; B = 8'h62; #100;
A = 8'h24; B = 8'h63; #100;
A = 8'h24; B = 8'h64; #100;
A = 8'h24; B = 8'h65; #100;
A = 8'h24; B = 8'h66; #100;
A = 8'h24; B = 8'h67; #100;
A = 8'h24; B = 8'h68; #100;
A = 8'h24; B = 8'h69; #100;
A = 8'h24; B = 8'h6A; #100;
A = 8'h24; B = 8'h6B; #100;
A = 8'h24; B = 8'h6C; #100;
A = 8'h24; B = 8'h6D; #100;
A = 8'h24; B = 8'h6E; #100;
A = 8'h24; B = 8'h6F; #100;
A = 8'h24; B = 8'h70; #100;
A = 8'h24; B = 8'h71; #100;
A = 8'h24; B = 8'h72; #100;
A = 8'h24; B = 8'h73; #100;
A = 8'h24; B = 8'h74; #100;
A = 8'h24; B = 8'h75; #100;
A = 8'h24; B = 8'h76; #100;
A = 8'h24; B = 8'h77; #100;
A = 8'h24; B = 8'h78; #100;
A = 8'h24; B = 8'h79; #100;
A = 8'h24; B = 8'h7A; #100;
A = 8'h24; B = 8'h7B; #100;
A = 8'h24; B = 8'h7C; #100;
A = 8'h24; B = 8'h7D; #100;
A = 8'h24; B = 8'h7E; #100;
A = 8'h24; B = 8'h7F; #100;
A = 8'h24; B = 8'h80; #100;
A = 8'h24; B = 8'h81; #100;
A = 8'h24; B = 8'h82; #100;
A = 8'h24; B = 8'h83; #100;
A = 8'h24; B = 8'h84; #100;
A = 8'h24; B = 8'h85; #100;
A = 8'h24; B = 8'h86; #100;
A = 8'h24; B = 8'h87; #100;
A = 8'h24; B = 8'h88; #100;
A = 8'h24; B = 8'h89; #100;
A = 8'h24; B = 8'h8A; #100;
A = 8'h24; B = 8'h8B; #100;
A = 8'h24; B = 8'h8C; #100;
A = 8'h24; B = 8'h8D; #100;
A = 8'h24; B = 8'h8E; #100;
A = 8'h24; B = 8'h8F; #100;
A = 8'h24; B = 8'h90; #100;
A = 8'h24; B = 8'h91; #100;
A = 8'h24; B = 8'h92; #100;
A = 8'h24; B = 8'h93; #100;
A = 8'h24; B = 8'h94; #100;
A = 8'h24; B = 8'h95; #100;
A = 8'h24; B = 8'h96; #100;
A = 8'h24; B = 8'h97; #100;
A = 8'h24; B = 8'h98; #100;
A = 8'h24; B = 8'h99; #100;
A = 8'h24; B = 8'h9A; #100;
A = 8'h24; B = 8'h9B; #100;
A = 8'h24; B = 8'h9C; #100;
A = 8'h24; B = 8'h9D; #100;
A = 8'h24; B = 8'h9E; #100;
A = 8'h24; B = 8'h9F; #100;
A = 8'h24; B = 8'hA0; #100;
A = 8'h24; B = 8'hA1; #100;
A = 8'h24; B = 8'hA2; #100;
A = 8'h24; B = 8'hA3; #100;
A = 8'h24; B = 8'hA4; #100;
A = 8'h24; B = 8'hA5; #100;
A = 8'h24; B = 8'hA6; #100;
A = 8'h24; B = 8'hA7; #100;
A = 8'h24; B = 8'hA8; #100;
A = 8'h24; B = 8'hA9; #100;
A = 8'h24; B = 8'hAA; #100;
A = 8'h24; B = 8'hAB; #100;
A = 8'h24; B = 8'hAC; #100;
A = 8'h24; B = 8'hAD; #100;
A = 8'h24; B = 8'hAE; #100;
A = 8'h24; B = 8'hAF; #100;
A = 8'h24; B = 8'hB0; #100;
A = 8'h24; B = 8'hB1; #100;
A = 8'h24; B = 8'hB2; #100;
A = 8'h24; B = 8'hB3; #100;
A = 8'h24; B = 8'hB4; #100;
A = 8'h24; B = 8'hB5; #100;
A = 8'h24; B = 8'hB6; #100;
A = 8'h24; B = 8'hB7; #100;
A = 8'h24; B = 8'hB8; #100;
A = 8'h24; B = 8'hB9; #100;
A = 8'h24; B = 8'hBA; #100;
A = 8'h24; B = 8'hBB; #100;
A = 8'h24; B = 8'hBC; #100;
A = 8'h24; B = 8'hBD; #100;
A = 8'h24; B = 8'hBE; #100;
A = 8'h24; B = 8'hBF; #100;
A = 8'h24; B = 8'hC0; #100;
A = 8'h24; B = 8'hC1; #100;
A = 8'h24; B = 8'hC2; #100;
A = 8'h24; B = 8'hC3; #100;
A = 8'h24; B = 8'hC4; #100;
A = 8'h24; B = 8'hC5; #100;
A = 8'h24; B = 8'hC6; #100;
A = 8'h24; B = 8'hC7; #100;
A = 8'h24; B = 8'hC8; #100;
A = 8'h24; B = 8'hC9; #100;
A = 8'h24; B = 8'hCA; #100;
A = 8'h24; B = 8'hCB; #100;
A = 8'h24; B = 8'hCC; #100;
A = 8'h24; B = 8'hCD; #100;
A = 8'h24; B = 8'hCE; #100;
A = 8'h24; B = 8'hCF; #100;
A = 8'h24; B = 8'hD0; #100;
A = 8'h24; B = 8'hD1; #100;
A = 8'h24; B = 8'hD2; #100;
A = 8'h24; B = 8'hD3; #100;
A = 8'h24; B = 8'hD4; #100;
A = 8'h24; B = 8'hD5; #100;
A = 8'h24; B = 8'hD6; #100;
A = 8'h24; B = 8'hD7; #100;
A = 8'h24; B = 8'hD8; #100;
A = 8'h24; B = 8'hD9; #100;
A = 8'h24; B = 8'hDA; #100;
A = 8'h24; B = 8'hDB; #100;
A = 8'h24; B = 8'hDC; #100;
A = 8'h24; B = 8'hDD; #100;
A = 8'h24; B = 8'hDE; #100;
A = 8'h24; B = 8'hDF; #100;
A = 8'h24; B = 8'hE0; #100;
A = 8'h24; B = 8'hE1; #100;
A = 8'h24; B = 8'hE2; #100;
A = 8'h24; B = 8'hE3; #100;
A = 8'h24; B = 8'hE4; #100;
A = 8'h24; B = 8'hE5; #100;
A = 8'h24; B = 8'hE6; #100;
A = 8'h24; B = 8'hE7; #100;
A = 8'h24; B = 8'hE8; #100;
A = 8'h24; B = 8'hE9; #100;
A = 8'h24; B = 8'hEA; #100;
A = 8'h24; B = 8'hEB; #100;
A = 8'h24; B = 8'hEC; #100;
A = 8'h24; B = 8'hED; #100;
A = 8'h24; B = 8'hEE; #100;
A = 8'h24; B = 8'hEF; #100;
A = 8'h24; B = 8'hF0; #100;
A = 8'h24; B = 8'hF1; #100;
A = 8'h24; B = 8'hF2; #100;
A = 8'h24; B = 8'hF3; #100;
A = 8'h24; B = 8'hF4; #100;
A = 8'h24; B = 8'hF5; #100;
A = 8'h24; B = 8'hF6; #100;
A = 8'h24; B = 8'hF7; #100;
A = 8'h24; B = 8'hF8; #100;
A = 8'h24; B = 8'hF9; #100;
A = 8'h24; B = 8'hFA; #100;
A = 8'h24; B = 8'hFB; #100;
A = 8'h24; B = 8'hFC; #100;
A = 8'h24; B = 8'hFD; #100;
A = 8'h24; B = 8'hFE; #100;
A = 8'h24; B = 8'hFF; #100;
A = 8'h25; B = 8'h0; #100;
A = 8'h25; B = 8'h1; #100;
A = 8'h25; B = 8'h2; #100;
A = 8'h25; B = 8'h3; #100;
A = 8'h25; B = 8'h4; #100;
A = 8'h25; B = 8'h5; #100;
A = 8'h25; B = 8'h6; #100;
A = 8'h25; B = 8'h7; #100;
A = 8'h25; B = 8'h8; #100;
A = 8'h25; B = 8'h9; #100;
A = 8'h25; B = 8'hA; #100;
A = 8'h25; B = 8'hB; #100;
A = 8'h25; B = 8'hC; #100;
A = 8'h25; B = 8'hD; #100;
A = 8'h25; B = 8'hE; #100;
A = 8'h25; B = 8'hF; #100;
A = 8'h25; B = 8'h10; #100;
A = 8'h25; B = 8'h11; #100;
A = 8'h25; B = 8'h12; #100;
A = 8'h25; B = 8'h13; #100;
A = 8'h25; B = 8'h14; #100;
A = 8'h25; B = 8'h15; #100;
A = 8'h25; B = 8'h16; #100;
A = 8'h25; B = 8'h17; #100;
A = 8'h25; B = 8'h18; #100;
A = 8'h25; B = 8'h19; #100;
A = 8'h25; B = 8'h1A; #100;
A = 8'h25; B = 8'h1B; #100;
A = 8'h25; B = 8'h1C; #100;
A = 8'h25; B = 8'h1D; #100;
A = 8'h25; B = 8'h1E; #100;
A = 8'h25; B = 8'h1F; #100;
A = 8'h25; B = 8'h20; #100;
A = 8'h25; B = 8'h21; #100;
A = 8'h25; B = 8'h22; #100;
A = 8'h25; B = 8'h23; #100;
A = 8'h25; B = 8'h24; #100;
A = 8'h25; B = 8'h25; #100;
A = 8'h25; B = 8'h26; #100;
A = 8'h25; B = 8'h27; #100;
A = 8'h25; B = 8'h28; #100;
A = 8'h25; B = 8'h29; #100;
A = 8'h25; B = 8'h2A; #100;
A = 8'h25; B = 8'h2B; #100;
A = 8'h25; B = 8'h2C; #100;
A = 8'h25; B = 8'h2D; #100;
A = 8'h25; B = 8'h2E; #100;
A = 8'h25; B = 8'h2F; #100;
A = 8'h25; B = 8'h30; #100;
A = 8'h25; B = 8'h31; #100;
A = 8'h25; B = 8'h32; #100;
A = 8'h25; B = 8'h33; #100;
A = 8'h25; B = 8'h34; #100;
A = 8'h25; B = 8'h35; #100;
A = 8'h25; B = 8'h36; #100;
A = 8'h25; B = 8'h37; #100;
A = 8'h25; B = 8'h38; #100;
A = 8'h25; B = 8'h39; #100;
A = 8'h25; B = 8'h3A; #100;
A = 8'h25; B = 8'h3B; #100;
A = 8'h25; B = 8'h3C; #100;
A = 8'h25; B = 8'h3D; #100;
A = 8'h25; B = 8'h3E; #100;
A = 8'h25; B = 8'h3F; #100;
A = 8'h25; B = 8'h40; #100;
A = 8'h25; B = 8'h41; #100;
A = 8'h25; B = 8'h42; #100;
A = 8'h25; B = 8'h43; #100;
A = 8'h25; B = 8'h44; #100;
A = 8'h25; B = 8'h45; #100;
A = 8'h25; B = 8'h46; #100;
A = 8'h25; B = 8'h47; #100;
A = 8'h25; B = 8'h48; #100;
A = 8'h25; B = 8'h49; #100;
A = 8'h25; B = 8'h4A; #100;
A = 8'h25; B = 8'h4B; #100;
A = 8'h25; B = 8'h4C; #100;
A = 8'h25; B = 8'h4D; #100;
A = 8'h25; B = 8'h4E; #100;
A = 8'h25; B = 8'h4F; #100;
A = 8'h25; B = 8'h50; #100;
A = 8'h25; B = 8'h51; #100;
A = 8'h25; B = 8'h52; #100;
A = 8'h25; B = 8'h53; #100;
A = 8'h25; B = 8'h54; #100;
A = 8'h25; B = 8'h55; #100;
A = 8'h25; B = 8'h56; #100;
A = 8'h25; B = 8'h57; #100;
A = 8'h25; B = 8'h58; #100;
A = 8'h25; B = 8'h59; #100;
A = 8'h25; B = 8'h5A; #100;
A = 8'h25; B = 8'h5B; #100;
A = 8'h25; B = 8'h5C; #100;
A = 8'h25; B = 8'h5D; #100;
A = 8'h25; B = 8'h5E; #100;
A = 8'h25; B = 8'h5F; #100;
A = 8'h25; B = 8'h60; #100;
A = 8'h25; B = 8'h61; #100;
A = 8'h25; B = 8'h62; #100;
A = 8'h25; B = 8'h63; #100;
A = 8'h25; B = 8'h64; #100;
A = 8'h25; B = 8'h65; #100;
A = 8'h25; B = 8'h66; #100;
A = 8'h25; B = 8'h67; #100;
A = 8'h25; B = 8'h68; #100;
A = 8'h25; B = 8'h69; #100;
A = 8'h25; B = 8'h6A; #100;
A = 8'h25; B = 8'h6B; #100;
A = 8'h25; B = 8'h6C; #100;
A = 8'h25; B = 8'h6D; #100;
A = 8'h25; B = 8'h6E; #100;
A = 8'h25; B = 8'h6F; #100;
A = 8'h25; B = 8'h70; #100;
A = 8'h25; B = 8'h71; #100;
A = 8'h25; B = 8'h72; #100;
A = 8'h25; B = 8'h73; #100;
A = 8'h25; B = 8'h74; #100;
A = 8'h25; B = 8'h75; #100;
A = 8'h25; B = 8'h76; #100;
A = 8'h25; B = 8'h77; #100;
A = 8'h25; B = 8'h78; #100;
A = 8'h25; B = 8'h79; #100;
A = 8'h25; B = 8'h7A; #100;
A = 8'h25; B = 8'h7B; #100;
A = 8'h25; B = 8'h7C; #100;
A = 8'h25; B = 8'h7D; #100;
A = 8'h25; B = 8'h7E; #100;
A = 8'h25; B = 8'h7F; #100;
A = 8'h25; B = 8'h80; #100;
A = 8'h25; B = 8'h81; #100;
A = 8'h25; B = 8'h82; #100;
A = 8'h25; B = 8'h83; #100;
A = 8'h25; B = 8'h84; #100;
A = 8'h25; B = 8'h85; #100;
A = 8'h25; B = 8'h86; #100;
A = 8'h25; B = 8'h87; #100;
A = 8'h25; B = 8'h88; #100;
A = 8'h25; B = 8'h89; #100;
A = 8'h25; B = 8'h8A; #100;
A = 8'h25; B = 8'h8B; #100;
A = 8'h25; B = 8'h8C; #100;
A = 8'h25; B = 8'h8D; #100;
A = 8'h25; B = 8'h8E; #100;
A = 8'h25; B = 8'h8F; #100;
A = 8'h25; B = 8'h90; #100;
A = 8'h25; B = 8'h91; #100;
A = 8'h25; B = 8'h92; #100;
A = 8'h25; B = 8'h93; #100;
A = 8'h25; B = 8'h94; #100;
A = 8'h25; B = 8'h95; #100;
A = 8'h25; B = 8'h96; #100;
A = 8'h25; B = 8'h97; #100;
A = 8'h25; B = 8'h98; #100;
A = 8'h25; B = 8'h99; #100;
A = 8'h25; B = 8'h9A; #100;
A = 8'h25; B = 8'h9B; #100;
A = 8'h25; B = 8'h9C; #100;
A = 8'h25; B = 8'h9D; #100;
A = 8'h25; B = 8'h9E; #100;
A = 8'h25; B = 8'h9F; #100;
A = 8'h25; B = 8'hA0; #100;
A = 8'h25; B = 8'hA1; #100;
A = 8'h25; B = 8'hA2; #100;
A = 8'h25; B = 8'hA3; #100;
A = 8'h25; B = 8'hA4; #100;
A = 8'h25; B = 8'hA5; #100;
A = 8'h25; B = 8'hA6; #100;
A = 8'h25; B = 8'hA7; #100;
A = 8'h25; B = 8'hA8; #100;
A = 8'h25; B = 8'hA9; #100;
A = 8'h25; B = 8'hAA; #100;
A = 8'h25; B = 8'hAB; #100;
A = 8'h25; B = 8'hAC; #100;
A = 8'h25; B = 8'hAD; #100;
A = 8'h25; B = 8'hAE; #100;
A = 8'h25; B = 8'hAF; #100;
A = 8'h25; B = 8'hB0; #100;
A = 8'h25; B = 8'hB1; #100;
A = 8'h25; B = 8'hB2; #100;
A = 8'h25; B = 8'hB3; #100;
A = 8'h25; B = 8'hB4; #100;
A = 8'h25; B = 8'hB5; #100;
A = 8'h25; B = 8'hB6; #100;
A = 8'h25; B = 8'hB7; #100;
A = 8'h25; B = 8'hB8; #100;
A = 8'h25; B = 8'hB9; #100;
A = 8'h25; B = 8'hBA; #100;
A = 8'h25; B = 8'hBB; #100;
A = 8'h25; B = 8'hBC; #100;
A = 8'h25; B = 8'hBD; #100;
A = 8'h25; B = 8'hBE; #100;
A = 8'h25; B = 8'hBF; #100;
A = 8'h25; B = 8'hC0; #100;
A = 8'h25; B = 8'hC1; #100;
A = 8'h25; B = 8'hC2; #100;
A = 8'h25; B = 8'hC3; #100;
A = 8'h25; B = 8'hC4; #100;
A = 8'h25; B = 8'hC5; #100;
A = 8'h25; B = 8'hC6; #100;
A = 8'h25; B = 8'hC7; #100;
A = 8'h25; B = 8'hC8; #100;
A = 8'h25; B = 8'hC9; #100;
A = 8'h25; B = 8'hCA; #100;
A = 8'h25; B = 8'hCB; #100;
A = 8'h25; B = 8'hCC; #100;
A = 8'h25; B = 8'hCD; #100;
A = 8'h25; B = 8'hCE; #100;
A = 8'h25; B = 8'hCF; #100;
A = 8'h25; B = 8'hD0; #100;
A = 8'h25; B = 8'hD1; #100;
A = 8'h25; B = 8'hD2; #100;
A = 8'h25; B = 8'hD3; #100;
A = 8'h25; B = 8'hD4; #100;
A = 8'h25; B = 8'hD5; #100;
A = 8'h25; B = 8'hD6; #100;
A = 8'h25; B = 8'hD7; #100;
A = 8'h25; B = 8'hD8; #100;
A = 8'h25; B = 8'hD9; #100;
A = 8'h25; B = 8'hDA; #100;
A = 8'h25; B = 8'hDB; #100;
A = 8'h25; B = 8'hDC; #100;
A = 8'h25; B = 8'hDD; #100;
A = 8'h25; B = 8'hDE; #100;
A = 8'h25; B = 8'hDF; #100;
A = 8'h25; B = 8'hE0; #100;
A = 8'h25; B = 8'hE1; #100;
A = 8'h25; B = 8'hE2; #100;
A = 8'h25; B = 8'hE3; #100;
A = 8'h25; B = 8'hE4; #100;
A = 8'h25; B = 8'hE5; #100;
A = 8'h25; B = 8'hE6; #100;
A = 8'h25; B = 8'hE7; #100;
A = 8'h25; B = 8'hE8; #100;
A = 8'h25; B = 8'hE9; #100;
A = 8'h25; B = 8'hEA; #100;
A = 8'h25; B = 8'hEB; #100;
A = 8'h25; B = 8'hEC; #100;
A = 8'h25; B = 8'hED; #100;
A = 8'h25; B = 8'hEE; #100;
A = 8'h25; B = 8'hEF; #100;
A = 8'h25; B = 8'hF0; #100;
A = 8'h25; B = 8'hF1; #100;
A = 8'h25; B = 8'hF2; #100;
A = 8'h25; B = 8'hF3; #100;
A = 8'h25; B = 8'hF4; #100;
A = 8'h25; B = 8'hF5; #100;
A = 8'h25; B = 8'hF6; #100;
A = 8'h25; B = 8'hF7; #100;
A = 8'h25; B = 8'hF8; #100;
A = 8'h25; B = 8'hF9; #100;
A = 8'h25; B = 8'hFA; #100;
A = 8'h25; B = 8'hFB; #100;
A = 8'h25; B = 8'hFC; #100;
A = 8'h25; B = 8'hFD; #100;
A = 8'h25; B = 8'hFE; #100;
A = 8'h25; B = 8'hFF; #100;
A = 8'h26; B = 8'h0; #100;
A = 8'h26; B = 8'h1; #100;
A = 8'h26; B = 8'h2; #100;
A = 8'h26; B = 8'h3; #100;
A = 8'h26; B = 8'h4; #100;
A = 8'h26; B = 8'h5; #100;
A = 8'h26; B = 8'h6; #100;
A = 8'h26; B = 8'h7; #100;
A = 8'h26; B = 8'h8; #100;
A = 8'h26; B = 8'h9; #100;
A = 8'h26; B = 8'hA; #100;
A = 8'h26; B = 8'hB; #100;
A = 8'h26; B = 8'hC; #100;
A = 8'h26; B = 8'hD; #100;
A = 8'h26; B = 8'hE; #100;
A = 8'h26; B = 8'hF; #100;
A = 8'h26; B = 8'h10; #100;
A = 8'h26; B = 8'h11; #100;
A = 8'h26; B = 8'h12; #100;
A = 8'h26; B = 8'h13; #100;
A = 8'h26; B = 8'h14; #100;
A = 8'h26; B = 8'h15; #100;
A = 8'h26; B = 8'h16; #100;
A = 8'h26; B = 8'h17; #100;
A = 8'h26; B = 8'h18; #100;
A = 8'h26; B = 8'h19; #100;
A = 8'h26; B = 8'h1A; #100;
A = 8'h26; B = 8'h1B; #100;
A = 8'h26; B = 8'h1C; #100;
A = 8'h26; B = 8'h1D; #100;
A = 8'h26; B = 8'h1E; #100;
A = 8'h26; B = 8'h1F; #100;
A = 8'h26; B = 8'h20; #100;
A = 8'h26; B = 8'h21; #100;
A = 8'h26; B = 8'h22; #100;
A = 8'h26; B = 8'h23; #100;
A = 8'h26; B = 8'h24; #100;
A = 8'h26; B = 8'h25; #100;
A = 8'h26; B = 8'h26; #100;
A = 8'h26; B = 8'h27; #100;
A = 8'h26; B = 8'h28; #100;
A = 8'h26; B = 8'h29; #100;
A = 8'h26; B = 8'h2A; #100;
A = 8'h26; B = 8'h2B; #100;
A = 8'h26; B = 8'h2C; #100;
A = 8'h26; B = 8'h2D; #100;
A = 8'h26; B = 8'h2E; #100;
A = 8'h26; B = 8'h2F; #100;
A = 8'h26; B = 8'h30; #100;
A = 8'h26; B = 8'h31; #100;
A = 8'h26; B = 8'h32; #100;
A = 8'h26; B = 8'h33; #100;
A = 8'h26; B = 8'h34; #100;
A = 8'h26; B = 8'h35; #100;
A = 8'h26; B = 8'h36; #100;
A = 8'h26; B = 8'h37; #100;
A = 8'h26; B = 8'h38; #100;
A = 8'h26; B = 8'h39; #100;
A = 8'h26; B = 8'h3A; #100;
A = 8'h26; B = 8'h3B; #100;
A = 8'h26; B = 8'h3C; #100;
A = 8'h26; B = 8'h3D; #100;
A = 8'h26; B = 8'h3E; #100;
A = 8'h26; B = 8'h3F; #100;
A = 8'h26; B = 8'h40; #100;
A = 8'h26; B = 8'h41; #100;
A = 8'h26; B = 8'h42; #100;
A = 8'h26; B = 8'h43; #100;
A = 8'h26; B = 8'h44; #100;
A = 8'h26; B = 8'h45; #100;
A = 8'h26; B = 8'h46; #100;
A = 8'h26; B = 8'h47; #100;
A = 8'h26; B = 8'h48; #100;
A = 8'h26; B = 8'h49; #100;
A = 8'h26; B = 8'h4A; #100;
A = 8'h26; B = 8'h4B; #100;
A = 8'h26; B = 8'h4C; #100;
A = 8'h26; B = 8'h4D; #100;
A = 8'h26; B = 8'h4E; #100;
A = 8'h26; B = 8'h4F; #100;
A = 8'h26; B = 8'h50; #100;
A = 8'h26; B = 8'h51; #100;
A = 8'h26; B = 8'h52; #100;
A = 8'h26; B = 8'h53; #100;
A = 8'h26; B = 8'h54; #100;
A = 8'h26; B = 8'h55; #100;
A = 8'h26; B = 8'h56; #100;
A = 8'h26; B = 8'h57; #100;
A = 8'h26; B = 8'h58; #100;
A = 8'h26; B = 8'h59; #100;
A = 8'h26; B = 8'h5A; #100;
A = 8'h26; B = 8'h5B; #100;
A = 8'h26; B = 8'h5C; #100;
A = 8'h26; B = 8'h5D; #100;
A = 8'h26; B = 8'h5E; #100;
A = 8'h26; B = 8'h5F; #100;
A = 8'h26; B = 8'h60; #100;
A = 8'h26; B = 8'h61; #100;
A = 8'h26; B = 8'h62; #100;
A = 8'h26; B = 8'h63; #100;
A = 8'h26; B = 8'h64; #100;
A = 8'h26; B = 8'h65; #100;
A = 8'h26; B = 8'h66; #100;
A = 8'h26; B = 8'h67; #100;
A = 8'h26; B = 8'h68; #100;
A = 8'h26; B = 8'h69; #100;
A = 8'h26; B = 8'h6A; #100;
A = 8'h26; B = 8'h6B; #100;
A = 8'h26; B = 8'h6C; #100;
A = 8'h26; B = 8'h6D; #100;
A = 8'h26; B = 8'h6E; #100;
A = 8'h26; B = 8'h6F; #100;
A = 8'h26; B = 8'h70; #100;
A = 8'h26; B = 8'h71; #100;
A = 8'h26; B = 8'h72; #100;
A = 8'h26; B = 8'h73; #100;
A = 8'h26; B = 8'h74; #100;
A = 8'h26; B = 8'h75; #100;
A = 8'h26; B = 8'h76; #100;
A = 8'h26; B = 8'h77; #100;
A = 8'h26; B = 8'h78; #100;
A = 8'h26; B = 8'h79; #100;
A = 8'h26; B = 8'h7A; #100;
A = 8'h26; B = 8'h7B; #100;
A = 8'h26; B = 8'h7C; #100;
A = 8'h26; B = 8'h7D; #100;
A = 8'h26; B = 8'h7E; #100;
A = 8'h26; B = 8'h7F; #100;
A = 8'h26; B = 8'h80; #100;
A = 8'h26; B = 8'h81; #100;
A = 8'h26; B = 8'h82; #100;
A = 8'h26; B = 8'h83; #100;
A = 8'h26; B = 8'h84; #100;
A = 8'h26; B = 8'h85; #100;
A = 8'h26; B = 8'h86; #100;
A = 8'h26; B = 8'h87; #100;
A = 8'h26; B = 8'h88; #100;
A = 8'h26; B = 8'h89; #100;
A = 8'h26; B = 8'h8A; #100;
A = 8'h26; B = 8'h8B; #100;
A = 8'h26; B = 8'h8C; #100;
A = 8'h26; B = 8'h8D; #100;
A = 8'h26; B = 8'h8E; #100;
A = 8'h26; B = 8'h8F; #100;
A = 8'h26; B = 8'h90; #100;
A = 8'h26; B = 8'h91; #100;
A = 8'h26; B = 8'h92; #100;
A = 8'h26; B = 8'h93; #100;
A = 8'h26; B = 8'h94; #100;
A = 8'h26; B = 8'h95; #100;
A = 8'h26; B = 8'h96; #100;
A = 8'h26; B = 8'h97; #100;
A = 8'h26; B = 8'h98; #100;
A = 8'h26; B = 8'h99; #100;
A = 8'h26; B = 8'h9A; #100;
A = 8'h26; B = 8'h9B; #100;
A = 8'h26; B = 8'h9C; #100;
A = 8'h26; B = 8'h9D; #100;
A = 8'h26; B = 8'h9E; #100;
A = 8'h26; B = 8'h9F; #100;
A = 8'h26; B = 8'hA0; #100;
A = 8'h26; B = 8'hA1; #100;
A = 8'h26; B = 8'hA2; #100;
A = 8'h26; B = 8'hA3; #100;
A = 8'h26; B = 8'hA4; #100;
A = 8'h26; B = 8'hA5; #100;
A = 8'h26; B = 8'hA6; #100;
A = 8'h26; B = 8'hA7; #100;
A = 8'h26; B = 8'hA8; #100;
A = 8'h26; B = 8'hA9; #100;
A = 8'h26; B = 8'hAA; #100;
A = 8'h26; B = 8'hAB; #100;
A = 8'h26; B = 8'hAC; #100;
A = 8'h26; B = 8'hAD; #100;
A = 8'h26; B = 8'hAE; #100;
A = 8'h26; B = 8'hAF; #100;
A = 8'h26; B = 8'hB0; #100;
A = 8'h26; B = 8'hB1; #100;
A = 8'h26; B = 8'hB2; #100;
A = 8'h26; B = 8'hB3; #100;
A = 8'h26; B = 8'hB4; #100;
A = 8'h26; B = 8'hB5; #100;
A = 8'h26; B = 8'hB6; #100;
A = 8'h26; B = 8'hB7; #100;
A = 8'h26; B = 8'hB8; #100;
A = 8'h26; B = 8'hB9; #100;
A = 8'h26; B = 8'hBA; #100;
A = 8'h26; B = 8'hBB; #100;
A = 8'h26; B = 8'hBC; #100;
A = 8'h26; B = 8'hBD; #100;
A = 8'h26; B = 8'hBE; #100;
A = 8'h26; B = 8'hBF; #100;
A = 8'h26; B = 8'hC0; #100;
A = 8'h26; B = 8'hC1; #100;
A = 8'h26; B = 8'hC2; #100;
A = 8'h26; B = 8'hC3; #100;
A = 8'h26; B = 8'hC4; #100;
A = 8'h26; B = 8'hC5; #100;
A = 8'h26; B = 8'hC6; #100;
A = 8'h26; B = 8'hC7; #100;
A = 8'h26; B = 8'hC8; #100;
A = 8'h26; B = 8'hC9; #100;
A = 8'h26; B = 8'hCA; #100;
A = 8'h26; B = 8'hCB; #100;
A = 8'h26; B = 8'hCC; #100;
A = 8'h26; B = 8'hCD; #100;
A = 8'h26; B = 8'hCE; #100;
A = 8'h26; B = 8'hCF; #100;
A = 8'h26; B = 8'hD0; #100;
A = 8'h26; B = 8'hD1; #100;
A = 8'h26; B = 8'hD2; #100;
A = 8'h26; B = 8'hD3; #100;
A = 8'h26; B = 8'hD4; #100;
A = 8'h26; B = 8'hD5; #100;
A = 8'h26; B = 8'hD6; #100;
A = 8'h26; B = 8'hD7; #100;
A = 8'h26; B = 8'hD8; #100;
A = 8'h26; B = 8'hD9; #100;
A = 8'h26; B = 8'hDA; #100;
A = 8'h26; B = 8'hDB; #100;
A = 8'h26; B = 8'hDC; #100;
A = 8'h26; B = 8'hDD; #100;
A = 8'h26; B = 8'hDE; #100;
A = 8'h26; B = 8'hDF; #100;
A = 8'h26; B = 8'hE0; #100;
A = 8'h26; B = 8'hE1; #100;
A = 8'h26; B = 8'hE2; #100;
A = 8'h26; B = 8'hE3; #100;
A = 8'h26; B = 8'hE4; #100;
A = 8'h26; B = 8'hE5; #100;
A = 8'h26; B = 8'hE6; #100;
A = 8'h26; B = 8'hE7; #100;
A = 8'h26; B = 8'hE8; #100;
A = 8'h26; B = 8'hE9; #100;
A = 8'h26; B = 8'hEA; #100;
A = 8'h26; B = 8'hEB; #100;
A = 8'h26; B = 8'hEC; #100;
A = 8'h26; B = 8'hED; #100;
A = 8'h26; B = 8'hEE; #100;
A = 8'h26; B = 8'hEF; #100;
A = 8'h26; B = 8'hF0; #100;
A = 8'h26; B = 8'hF1; #100;
A = 8'h26; B = 8'hF2; #100;
A = 8'h26; B = 8'hF3; #100;
A = 8'h26; B = 8'hF4; #100;
A = 8'h26; B = 8'hF5; #100;
A = 8'h26; B = 8'hF6; #100;
A = 8'h26; B = 8'hF7; #100;
A = 8'h26; B = 8'hF8; #100;
A = 8'h26; B = 8'hF9; #100;
A = 8'h26; B = 8'hFA; #100;
A = 8'h26; B = 8'hFB; #100;
A = 8'h26; B = 8'hFC; #100;
A = 8'h26; B = 8'hFD; #100;
A = 8'h26; B = 8'hFE; #100;
A = 8'h26; B = 8'hFF; #100;
A = 8'h27; B = 8'h0; #100;
A = 8'h27; B = 8'h1; #100;
A = 8'h27; B = 8'h2; #100;
A = 8'h27; B = 8'h3; #100;
A = 8'h27; B = 8'h4; #100;
A = 8'h27; B = 8'h5; #100;
A = 8'h27; B = 8'h6; #100;
A = 8'h27; B = 8'h7; #100;
A = 8'h27; B = 8'h8; #100;
A = 8'h27; B = 8'h9; #100;
A = 8'h27; B = 8'hA; #100;
A = 8'h27; B = 8'hB; #100;
A = 8'h27; B = 8'hC; #100;
A = 8'h27; B = 8'hD; #100;
A = 8'h27; B = 8'hE; #100;
A = 8'h27; B = 8'hF; #100;
A = 8'h27; B = 8'h10; #100;
A = 8'h27; B = 8'h11; #100;
A = 8'h27; B = 8'h12; #100;
A = 8'h27; B = 8'h13; #100;
A = 8'h27; B = 8'h14; #100;
A = 8'h27; B = 8'h15; #100;
A = 8'h27; B = 8'h16; #100;
A = 8'h27; B = 8'h17; #100;
A = 8'h27; B = 8'h18; #100;
A = 8'h27; B = 8'h19; #100;
A = 8'h27; B = 8'h1A; #100;
A = 8'h27; B = 8'h1B; #100;
A = 8'h27; B = 8'h1C; #100;
A = 8'h27; B = 8'h1D; #100;
A = 8'h27; B = 8'h1E; #100;
A = 8'h27; B = 8'h1F; #100;
A = 8'h27; B = 8'h20; #100;
A = 8'h27; B = 8'h21; #100;
A = 8'h27; B = 8'h22; #100;
A = 8'h27; B = 8'h23; #100;
A = 8'h27; B = 8'h24; #100;
A = 8'h27; B = 8'h25; #100;
A = 8'h27; B = 8'h26; #100;
A = 8'h27; B = 8'h27; #100;
A = 8'h27; B = 8'h28; #100;
A = 8'h27; B = 8'h29; #100;
A = 8'h27; B = 8'h2A; #100;
A = 8'h27; B = 8'h2B; #100;
A = 8'h27; B = 8'h2C; #100;
A = 8'h27; B = 8'h2D; #100;
A = 8'h27; B = 8'h2E; #100;
A = 8'h27; B = 8'h2F; #100;
A = 8'h27; B = 8'h30; #100;
A = 8'h27; B = 8'h31; #100;
A = 8'h27; B = 8'h32; #100;
A = 8'h27; B = 8'h33; #100;
A = 8'h27; B = 8'h34; #100;
A = 8'h27; B = 8'h35; #100;
A = 8'h27; B = 8'h36; #100;
A = 8'h27; B = 8'h37; #100;
A = 8'h27; B = 8'h38; #100;
A = 8'h27; B = 8'h39; #100;
A = 8'h27; B = 8'h3A; #100;
A = 8'h27; B = 8'h3B; #100;
A = 8'h27; B = 8'h3C; #100;
A = 8'h27; B = 8'h3D; #100;
A = 8'h27; B = 8'h3E; #100;
A = 8'h27; B = 8'h3F; #100;
A = 8'h27; B = 8'h40; #100;
A = 8'h27; B = 8'h41; #100;
A = 8'h27; B = 8'h42; #100;
A = 8'h27; B = 8'h43; #100;
A = 8'h27; B = 8'h44; #100;
A = 8'h27; B = 8'h45; #100;
A = 8'h27; B = 8'h46; #100;
A = 8'h27; B = 8'h47; #100;
A = 8'h27; B = 8'h48; #100;
A = 8'h27; B = 8'h49; #100;
A = 8'h27; B = 8'h4A; #100;
A = 8'h27; B = 8'h4B; #100;
A = 8'h27; B = 8'h4C; #100;
A = 8'h27; B = 8'h4D; #100;
A = 8'h27; B = 8'h4E; #100;
A = 8'h27; B = 8'h4F; #100;
A = 8'h27; B = 8'h50; #100;
A = 8'h27; B = 8'h51; #100;
A = 8'h27; B = 8'h52; #100;
A = 8'h27; B = 8'h53; #100;
A = 8'h27; B = 8'h54; #100;
A = 8'h27; B = 8'h55; #100;
A = 8'h27; B = 8'h56; #100;
A = 8'h27; B = 8'h57; #100;
A = 8'h27; B = 8'h58; #100;
A = 8'h27; B = 8'h59; #100;
A = 8'h27; B = 8'h5A; #100;
A = 8'h27; B = 8'h5B; #100;
A = 8'h27; B = 8'h5C; #100;
A = 8'h27; B = 8'h5D; #100;
A = 8'h27; B = 8'h5E; #100;
A = 8'h27; B = 8'h5F; #100;
A = 8'h27; B = 8'h60; #100;
A = 8'h27; B = 8'h61; #100;
A = 8'h27; B = 8'h62; #100;
A = 8'h27; B = 8'h63; #100;
A = 8'h27; B = 8'h64; #100;
A = 8'h27; B = 8'h65; #100;
A = 8'h27; B = 8'h66; #100;
A = 8'h27; B = 8'h67; #100;
A = 8'h27; B = 8'h68; #100;
A = 8'h27; B = 8'h69; #100;
A = 8'h27; B = 8'h6A; #100;
A = 8'h27; B = 8'h6B; #100;
A = 8'h27; B = 8'h6C; #100;
A = 8'h27; B = 8'h6D; #100;
A = 8'h27; B = 8'h6E; #100;
A = 8'h27; B = 8'h6F; #100;
A = 8'h27; B = 8'h70; #100;
A = 8'h27; B = 8'h71; #100;
A = 8'h27; B = 8'h72; #100;
A = 8'h27; B = 8'h73; #100;
A = 8'h27; B = 8'h74; #100;
A = 8'h27; B = 8'h75; #100;
A = 8'h27; B = 8'h76; #100;
A = 8'h27; B = 8'h77; #100;
A = 8'h27; B = 8'h78; #100;
A = 8'h27; B = 8'h79; #100;
A = 8'h27; B = 8'h7A; #100;
A = 8'h27; B = 8'h7B; #100;
A = 8'h27; B = 8'h7C; #100;
A = 8'h27; B = 8'h7D; #100;
A = 8'h27; B = 8'h7E; #100;
A = 8'h27; B = 8'h7F; #100;
A = 8'h27; B = 8'h80; #100;
A = 8'h27; B = 8'h81; #100;
A = 8'h27; B = 8'h82; #100;
A = 8'h27; B = 8'h83; #100;
A = 8'h27; B = 8'h84; #100;
A = 8'h27; B = 8'h85; #100;
A = 8'h27; B = 8'h86; #100;
A = 8'h27; B = 8'h87; #100;
A = 8'h27; B = 8'h88; #100;
A = 8'h27; B = 8'h89; #100;
A = 8'h27; B = 8'h8A; #100;
A = 8'h27; B = 8'h8B; #100;
A = 8'h27; B = 8'h8C; #100;
A = 8'h27; B = 8'h8D; #100;
A = 8'h27; B = 8'h8E; #100;
A = 8'h27; B = 8'h8F; #100;
A = 8'h27; B = 8'h90; #100;
A = 8'h27; B = 8'h91; #100;
A = 8'h27; B = 8'h92; #100;
A = 8'h27; B = 8'h93; #100;
A = 8'h27; B = 8'h94; #100;
A = 8'h27; B = 8'h95; #100;
A = 8'h27; B = 8'h96; #100;
A = 8'h27; B = 8'h97; #100;
A = 8'h27; B = 8'h98; #100;
A = 8'h27; B = 8'h99; #100;
A = 8'h27; B = 8'h9A; #100;
A = 8'h27; B = 8'h9B; #100;
A = 8'h27; B = 8'h9C; #100;
A = 8'h27; B = 8'h9D; #100;
A = 8'h27; B = 8'h9E; #100;
A = 8'h27; B = 8'h9F; #100;
A = 8'h27; B = 8'hA0; #100;
A = 8'h27; B = 8'hA1; #100;
A = 8'h27; B = 8'hA2; #100;
A = 8'h27; B = 8'hA3; #100;
A = 8'h27; B = 8'hA4; #100;
A = 8'h27; B = 8'hA5; #100;
A = 8'h27; B = 8'hA6; #100;
A = 8'h27; B = 8'hA7; #100;
A = 8'h27; B = 8'hA8; #100;
A = 8'h27; B = 8'hA9; #100;
A = 8'h27; B = 8'hAA; #100;
A = 8'h27; B = 8'hAB; #100;
A = 8'h27; B = 8'hAC; #100;
A = 8'h27; B = 8'hAD; #100;
A = 8'h27; B = 8'hAE; #100;
A = 8'h27; B = 8'hAF; #100;
A = 8'h27; B = 8'hB0; #100;
A = 8'h27; B = 8'hB1; #100;
A = 8'h27; B = 8'hB2; #100;
A = 8'h27; B = 8'hB3; #100;
A = 8'h27; B = 8'hB4; #100;
A = 8'h27; B = 8'hB5; #100;
A = 8'h27; B = 8'hB6; #100;
A = 8'h27; B = 8'hB7; #100;
A = 8'h27; B = 8'hB8; #100;
A = 8'h27; B = 8'hB9; #100;
A = 8'h27; B = 8'hBA; #100;
A = 8'h27; B = 8'hBB; #100;
A = 8'h27; B = 8'hBC; #100;
A = 8'h27; B = 8'hBD; #100;
A = 8'h27; B = 8'hBE; #100;
A = 8'h27; B = 8'hBF; #100;
A = 8'h27; B = 8'hC0; #100;
A = 8'h27; B = 8'hC1; #100;
A = 8'h27; B = 8'hC2; #100;
A = 8'h27; B = 8'hC3; #100;
A = 8'h27; B = 8'hC4; #100;
A = 8'h27; B = 8'hC5; #100;
A = 8'h27; B = 8'hC6; #100;
A = 8'h27; B = 8'hC7; #100;
A = 8'h27; B = 8'hC8; #100;
A = 8'h27; B = 8'hC9; #100;
A = 8'h27; B = 8'hCA; #100;
A = 8'h27; B = 8'hCB; #100;
A = 8'h27; B = 8'hCC; #100;
A = 8'h27; B = 8'hCD; #100;
A = 8'h27; B = 8'hCE; #100;
A = 8'h27; B = 8'hCF; #100;
A = 8'h27; B = 8'hD0; #100;
A = 8'h27; B = 8'hD1; #100;
A = 8'h27; B = 8'hD2; #100;
A = 8'h27; B = 8'hD3; #100;
A = 8'h27; B = 8'hD4; #100;
A = 8'h27; B = 8'hD5; #100;
A = 8'h27; B = 8'hD6; #100;
A = 8'h27; B = 8'hD7; #100;
A = 8'h27; B = 8'hD8; #100;
A = 8'h27; B = 8'hD9; #100;
A = 8'h27; B = 8'hDA; #100;
A = 8'h27; B = 8'hDB; #100;
A = 8'h27; B = 8'hDC; #100;
A = 8'h27; B = 8'hDD; #100;
A = 8'h27; B = 8'hDE; #100;
A = 8'h27; B = 8'hDF; #100;
A = 8'h27; B = 8'hE0; #100;
A = 8'h27; B = 8'hE1; #100;
A = 8'h27; B = 8'hE2; #100;
A = 8'h27; B = 8'hE3; #100;
A = 8'h27; B = 8'hE4; #100;
A = 8'h27; B = 8'hE5; #100;
A = 8'h27; B = 8'hE6; #100;
A = 8'h27; B = 8'hE7; #100;
A = 8'h27; B = 8'hE8; #100;
A = 8'h27; B = 8'hE9; #100;
A = 8'h27; B = 8'hEA; #100;
A = 8'h27; B = 8'hEB; #100;
A = 8'h27; B = 8'hEC; #100;
A = 8'h27; B = 8'hED; #100;
A = 8'h27; B = 8'hEE; #100;
A = 8'h27; B = 8'hEF; #100;
A = 8'h27; B = 8'hF0; #100;
A = 8'h27; B = 8'hF1; #100;
A = 8'h27; B = 8'hF2; #100;
A = 8'h27; B = 8'hF3; #100;
A = 8'h27; B = 8'hF4; #100;
A = 8'h27; B = 8'hF5; #100;
A = 8'h27; B = 8'hF6; #100;
A = 8'h27; B = 8'hF7; #100;
A = 8'h27; B = 8'hF8; #100;
A = 8'h27; B = 8'hF9; #100;
A = 8'h27; B = 8'hFA; #100;
A = 8'h27; B = 8'hFB; #100;
A = 8'h27; B = 8'hFC; #100;
A = 8'h27; B = 8'hFD; #100;
A = 8'h27; B = 8'hFE; #100;
A = 8'h27; B = 8'hFF; #100;
A = 8'h28; B = 8'h0; #100;
A = 8'h28; B = 8'h1; #100;
A = 8'h28; B = 8'h2; #100;
A = 8'h28; B = 8'h3; #100;
A = 8'h28; B = 8'h4; #100;
A = 8'h28; B = 8'h5; #100;
A = 8'h28; B = 8'h6; #100;
A = 8'h28; B = 8'h7; #100;
A = 8'h28; B = 8'h8; #100;
A = 8'h28; B = 8'h9; #100;
A = 8'h28; B = 8'hA; #100;
A = 8'h28; B = 8'hB; #100;
A = 8'h28; B = 8'hC; #100;
A = 8'h28; B = 8'hD; #100;
A = 8'h28; B = 8'hE; #100;
A = 8'h28; B = 8'hF; #100;
A = 8'h28; B = 8'h10; #100;
A = 8'h28; B = 8'h11; #100;
A = 8'h28; B = 8'h12; #100;
A = 8'h28; B = 8'h13; #100;
A = 8'h28; B = 8'h14; #100;
A = 8'h28; B = 8'h15; #100;
A = 8'h28; B = 8'h16; #100;
A = 8'h28; B = 8'h17; #100;
A = 8'h28; B = 8'h18; #100;
A = 8'h28; B = 8'h19; #100;
A = 8'h28; B = 8'h1A; #100;
A = 8'h28; B = 8'h1B; #100;
A = 8'h28; B = 8'h1C; #100;
A = 8'h28; B = 8'h1D; #100;
A = 8'h28; B = 8'h1E; #100;
A = 8'h28; B = 8'h1F; #100;
A = 8'h28; B = 8'h20; #100;
A = 8'h28; B = 8'h21; #100;
A = 8'h28; B = 8'h22; #100;
A = 8'h28; B = 8'h23; #100;
A = 8'h28; B = 8'h24; #100;
A = 8'h28; B = 8'h25; #100;
A = 8'h28; B = 8'h26; #100;
A = 8'h28; B = 8'h27; #100;
A = 8'h28; B = 8'h28; #100;
A = 8'h28; B = 8'h29; #100;
A = 8'h28; B = 8'h2A; #100;
A = 8'h28; B = 8'h2B; #100;
A = 8'h28; B = 8'h2C; #100;
A = 8'h28; B = 8'h2D; #100;
A = 8'h28; B = 8'h2E; #100;
A = 8'h28; B = 8'h2F; #100;
A = 8'h28; B = 8'h30; #100;
A = 8'h28; B = 8'h31; #100;
A = 8'h28; B = 8'h32; #100;
A = 8'h28; B = 8'h33; #100;
A = 8'h28; B = 8'h34; #100;
A = 8'h28; B = 8'h35; #100;
A = 8'h28; B = 8'h36; #100;
A = 8'h28; B = 8'h37; #100;
A = 8'h28; B = 8'h38; #100;
A = 8'h28; B = 8'h39; #100;
A = 8'h28; B = 8'h3A; #100;
A = 8'h28; B = 8'h3B; #100;
A = 8'h28; B = 8'h3C; #100;
A = 8'h28; B = 8'h3D; #100;
A = 8'h28; B = 8'h3E; #100;
A = 8'h28; B = 8'h3F; #100;
A = 8'h28; B = 8'h40; #100;
A = 8'h28; B = 8'h41; #100;
A = 8'h28; B = 8'h42; #100;
A = 8'h28; B = 8'h43; #100;
A = 8'h28; B = 8'h44; #100;
A = 8'h28; B = 8'h45; #100;
A = 8'h28; B = 8'h46; #100;
A = 8'h28; B = 8'h47; #100;
A = 8'h28; B = 8'h48; #100;
A = 8'h28; B = 8'h49; #100;
A = 8'h28; B = 8'h4A; #100;
A = 8'h28; B = 8'h4B; #100;
A = 8'h28; B = 8'h4C; #100;
A = 8'h28; B = 8'h4D; #100;
A = 8'h28; B = 8'h4E; #100;
A = 8'h28; B = 8'h4F; #100;
A = 8'h28; B = 8'h50; #100;
A = 8'h28; B = 8'h51; #100;
A = 8'h28; B = 8'h52; #100;
A = 8'h28; B = 8'h53; #100;
A = 8'h28; B = 8'h54; #100;
A = 8'h28; B = 8'h55; #100;
A = 8'h28; B = 8'h56; #100;
A = 8'h28; B = 8'h57; #100;
A = 8'h28; B = 8'h58; #100;
A = 8'h28; B = 8'h59; #100;
A = 8'h28; B = 8'h5A; #100;
A = 8'h28; B = 8'h5B; #100;
A = 8'h28; B = 8'h5C; #100;
A = 8'h28; B = 8'h5D; #100;
A = 8'h28; B = 8'h5E; #100;
A = 8'h28; B = 8'h5F; #100;
A = 8'h28; B = 8'h60; #100;
A = 8'h28; B = 8'h61; #100;
A = 8'h28; B = 8'h62; #100;
A = 8'h28; B = 8'h63; #100;
A = 8'h28; B = 8'h64; #100;
A = 8'h28; B = 8'h65; #100;
A = 8'h28; B = 8'h66; #100;
A = 8'h28; B = 8'h67; #100;
A = 8'h28; B = 8'h68; #100;
A = 8'h28; B = 8'h69; #100;
A = 8'h28; B = 8'h6A; #100;
A = 8'h28; B = 8'h6B; #100;
A = 8'h28; B = 8'h6C; #100;
A = 8'h28; B = 8'h6D; #100;
A = 8'h28; B = 8'h6E; #100;
A = 8'h28; B = 8'h6F; #100;
A = 8'h28; B = 8'h70; #100;
A = 8'h28; B = 8'h71; #100;
A = 8'h28; B = 8'h72; #100;
A = 8'h28; B = 8'h73; #100;
A = 8'h28; B = 8'h74; #100;
A = 8'h28; B = 8'h75; #100;
A = 8'h28; B = 8'h76; #100;
A = 8'h28; B = 8'h77; #100;
A = 8'h28; B = 8'h78; #100;
A = 8'h28; B = 8'h79; #100;
A = 8'h28; B = 8'h7A; #100;
A = 8'h28; B = 8'h7B; #100;
A = 8'h28; B = 8'h7C; #100;
A = 8'h28; B = 8'h7D; #100;
A = 8'h28; B = 8'h7E; #100;
A = 8'h28; B = 8'h7F; #100;
A = 8'h28; B = 8'h80; #100;
A = 8'h28; B = 8'h81; #100;
A = 8'h28; B = 8'h82; #100;
A = 8'h28; B = 8'h83; #100;
A = 8'h28; B = 8'h84; #100;
A = 8'h28; B = 8'h85; #100;
A = 8'h28; B = 8'h86; #100;
A = 8'h28; B = 8'h87; #100;
A = 8'h28; B = 8'h88; #100;
A = 8'h28; B = 8'h89; #100;
A = 8'h28; B = 8'h8A; #100;
A = 8'h28; B = 8'h8B; #100;
A = 8'h28; B = 8'h8C; #100;
A = 8'h28; B = 8'h8D; #100;
A = 8'h28; B = 8'h8E; #100;
A = 8'h28; B = 8'h8F; #100;
A = 8'h28; B = 8'h90; #100;
A = 8'h28; B = 8'h91; #100;
A = 8'h28; B = 8'h92; #100;
A = 8'h28; B = 8'h93; #100;
A = 8'h28; B = 8'h94; #100;
A = 8'h28; B = 8'h95; #100;
A = 8'h28; B = 8'h96; #100;
A = 8'h28; B = 8'h97; #100;
A = 8'h28; B = 8'h98; #100;
A = 8'h28; B = 8'h99; #100;
A = 8'h28; B = 8'h9A; #100;
A = 8'h28; B = 8'h9B; #100;
A = 8'h28; B = 8'h9C; #100;
A = 8'h28; B = 8'h9D; #100;
A = 8'h28; B = 8'h9E; #100;
A = 8'h28; B = 8'h9F; #100;
A = 8'h28; B = 8'hA0; #100;
A = 8'h28; B = 8'hA1; #100;
A = 8'h28; B = 8'hA2; #100;
A = 8'h28; B = 8'hA3; #100;
A = 8'h28; B = 8'hA4; #100;
A = 8'h28; B = 8'hA5; #100;
A = 8'h28; B = 8'hA6; #100;
A = 8'h28; B = 8'hA7; #100;
A = 8'h28; B = 8'hA8; #100;
A = 8'h28; B = 8'hA9; #100;
A = 8'h28; B = 8'hAA; #100;
A = 8'h28; B = 8'hAB; #100;
A = 8'h28; B = 8'hAC; #100;
A = 8'h28; B = 8'hAD; #100;
A = 8'h28; B = 8'hAE; #100;
A = 8'h28; B = 8'hAF; #100;
A = 8'h28; B = 8'hB0; #100;
A = 8'h28; B = 8'hB1; #100;
A = 8'h28; B = 8'hB2; #100;
A = 8'h28; B = 8'hB3; #100;
A = 8'h28; B = 8'hB4; #100;
A = 8'h28; B = 8'hB5; #100;
A = 8'h28; B = 8'hB6; #100;
A = 8'h28; B = 8'hB7; #100;
A = 8'h28; B = 8'hB8; #100;
A = 8'h28; B = 8'hB9; #100;
A = 8'h28; B = 8'hBA; #100;
A = 8'h28; B = 8'hBB; #100;
A = 8'h28; B = 8'hBC; #100;
A = 8'h28; B = 8'hBD; #100;
A = 8'h28; B = 8'hBE; #100;
A = 8'h28; B = 8'hBF; #100;
A = 8'h28; B = 8'hC0; #100;
A = 8'h28; B = 8'hC1; #100;
A = 8'h28; B = 8'hC2; #100;
A = 8'h28; B = 8'hC3; #100;
A = 8'h28; B = 8'hC4; #100;
A = 8'h28; B = 8'hC5; #100;
A = 8'h28; B = 8'hC6; #100;
A = 8'h28; B = 8'hC7; #100;
A = 8'h28; B = 8'hC8; #100;
A = 8'h28; B = 8'hC9; #100;
A = 8'h28; B = 8'hCA; #100;
A = 8'h28; B = 8'hCB; #100;
A = 8'h28; B = 8'hCC; #100;
A = 8'h28; B = 8'hCD; #100;
A = 8'h28; B = 8'hCE; #100;
A = 8'h28; B = 8'hCF; #100;
A = 8'h28; B = 8'hD0; #100;
A = 8'h28; B = 8'hD1; #100;
A = 8'h28; B = 8'hD2; #100;
A = 8'h28; B = 8'hD3; #100;
A = 8'h28; B = 8'hD4; #100;
A = 8'h28; B = 8'hD5; #100;
A = 8'h28; B = 8'hD6; #100;
A = 8'h28; B = 8'hD7; #100;
A = 8'h28; B = 8'hD8; #100;
A = 8'h28; B = 8'hD9; #100;
A = 8'h28; B = 8'hDA; #100;
A = 8'h28; B = 8'hDB; #100;
A = 8'h28; B = 8'hDC; #100;
A = 8'h28; B = 8'hDD; #100;
A = 8'h28; B = 8'hDE; #100;
A = 8'h28; B = 8'hDF; #100;
A = 8'h28; B = 8'hE0; #100;
A = 8'h28; B = 8'hE1; #100;
A = 8'h28; B = 8'hE2; #100;
A = 8'h28; B = 8'hE3; #100;
A = 8'h28; B = 8'hE4; #100;
A = 8'h28; B = 8'hE5; #100;
A = 8'h28; B = 8'hE6; #100;
A = 8'h28; B = 8'hE7; #100;
A = 8'h28; B = 8'hE8; #100;
A = 8'h28; B = 8'hE9; #100;
A = 8'h28; B = 8'hEA; #100;
A = 8'h28; B = 8'hEB; #100;
A = 8'h28; B = 8'hEC; #100;
A = 8'h28; B = 8'hED; #100;
A = 8'h28; B = 8'hEE; #100;
A = 8'h28; B = 8'hEF; #100;
A = 8'h28; B = 8'hF0; #100;
A = 8'h28; B = 8'hF1; #100;
A = 8'h28; B = 8'hF2; #100;
A = 8'h28; B = 8'hF3; #100;
A = 8'h28; B = 8'hF4; #100;
A = 8'h28; B = 8'hF5; #100;
A = 8'h28; B = 8'hF6; #100;
A = 8'h28; B = 8'hF7; #100;
A = 8'h28; B = 8'hF8; #100;
A = 8'h28; B = 8'hF9; #100;
A = 8'h28; B = 8'hFA; #100;
A = 8'h28; B = 8'hFB; #100;
A = 8'h28; B = 8'hFC; #100;
A = 8'h28; B = 8'hFD; #100;
A = 8'h28; B = 8'hFE; #100;
A = 8'h28; B = 8'hFF; #100;
A = 8'h29; B = 8'h0; #100;
A = 8'h29; B = 8'h1; #100;
A = 8'h29; B = 8'h2; #100;
A = 8'h29; B = 8'h3; #100;
A = 8'h29; B = 8'h4; #100;
A = 8'h29; B = 8'h5; #100;
A = 8'h29; B = 8'h6; #100;
A = 8'h29; B = 8'h7; #100;
A = 8'h29; B = 8'h8; #100;
A = 8'h29; B = 8'h9; #100;
A = 8'h29; B = 8'hA; #100;
A = 8'h29; B = 8'hB; #100;
A = 8'h29; B = 8'hC; #100;
A = 8'h29; B = 8'hD; #100;
A = 8'h29; B = 8'hE; #100;
A = 8'h29; B = 8'hF; #100;
A = 8'h29; B = 8'h10; #100;
A = 8'h29; B = 8'h11; #100;
A = 8'h29; B = 8'h12; #100;
A = 8'h29; B = 8'h13; #100;
A = 8'h29; B = 8'h14; #100;
A = 8'h29; B = 8'h15; #100;
A = 8'h29; B = 8'h16; #100;
A = 8'h29; B = 8'h17; #100;
A = 8'h29; B = 8'h18; #100;
A = 8'h29; B = 8'h19; #100;
A = 8'h29; B = 8'h1A; #100;
A = 8'h29; B = 8'h1B; #100;
A = 8'h29; B = 8'h1C; #100;
A = 8'h29; B = 8'h1D; #100;
A = 8'h29; B = 8'h1E; #100;
A = 8'h29; B = 8'h1F; #100;
A = 8'h29; B = 8'h20; #100;
A = 8'h29; B = 8'h21; #100;
A = 8'h29; B = 8'h22; #100;
A = 8'h29; B = 8'h23; #100;
A = 8'h29; B = 8'h24; #100;
A = 8'h29; B = 8'h25; #100;
A = 8'h29; B = 8'h26; #100;
A = 8'h29; B = 8'h27; #100;
A = 8'h29; B = 8'h28; #100;
A = 8'h29; B = 8'h29; #100;
A = 8'h29; B = 8'h2A; #100;
A = 8'h29; B = 8'h2B; #100;
A = 8'h29; B = 8'h2C; #100;
A = 8'h29; B = 8'h2D; #100;
A = 8'h29; B = 8'h2E; #100;
A = 8'h29; B = 8'h2F; #100;
A = 8'h29; B = 8'h30; #100;
A = 8'h29; B = 8'h31; #100;
A = 8'h29; B = 8'h32; #100;
A = 8'h29; B = 8'h33; #100;
A = 8'h29; B = 8'h34; #100;
A = 8'h29; B = 8'h35; #100;
A = 8'h29; B = 8'h36; #100;
A = 8'h29; B = 8'h37; #100;
A = 8'h29; B = 8'h38; #100;
A = 8'h29; B = 8'h39; #100;
A = 8'h29; B = 8'h3A; #100;
A = 8'h29; B = 8'h3B; #100;
A = 8'h29; B = 8'h3C; #100;
A = 8'h29; B = 8'h3D; #100;
A = 8'h29; B = 8'h3E; #100;
A = 8'h29; B = 8'h3F; #100;
A = 8'h29; B = 8'h40; #100;
A = 8'h29; B = 8'h41; #100;
A = 8'h29; B = 8'h42; #100;
A = 8'h29; B = 8'h43; #100;
A = 8'h29; B = 8'h44; #100;
A = 8'h29; B = 8'h45; #100;
A = 8'h29; B = 8'h46; #100;
A = 8'h29; B = 8'h47; #100;
A = 8'h29; B = 8'h48; #100;
A = 8'h29; B = 8'h49; #100;
A = 8'h29; B = 8'h4A; #100;
A = 8'h29; B = 8'h4B; #100;
A = 8'h29; B = 8'h4C; #100;
A = 8'h29; B = 8'h4D; #100;
A = 8'h29; B = 8'h4E; #100;
A = 8'h29; B = 8'h4F; #100;
A = 8'h29; B = 8'h50; #100;
A = 8'h29; B = 8'h51; #100;
A = 8'h29; B = 8'h52; #100;
A = 8'h29; B = 8'h53; #100;
A = 8'h29; B = 8'h54; #100;
A = 8'h29; B = 8'h55; #100;
A = 8'h29; B = 8'h56; #100;
A = 8'h29; B = 8'h57; #100;
A = 8'h29; B = 8'h58; #100;
A = 8'h29; B = 8'h59; #100;
A = 8'h29; B = 8'h5A; #100;
A = 8'h29; B = 8'h5B; #100;
A = 8'h29; B = 8'h5C; #100;
A = 8'h29; B = 8'h5D; #100;
A = 8'h29; B = 8'h5E; #100;
A = 8'h29; B = 8'h5F; #100;
A = 8'h29; B = 8'h60; #100;
A = 8'h29; B = 8'h61; #100;
A = 8'h29; B = 8'h62; #100;
A = 8'h29; B = 8'h63; #100;
A = 8'h29; B = 8'h64; #100;
A = 8'h29; B = 8'h65; #100;
A = 8'h29; B = 8'h66; #100;
A = 8'h29; B = 8'h67; #100;
A = 8'h29; B = 8'h68; #100;
A = 8'h29; B = 8'h69; #100;
A = 8'h29; B = 8'h6A; #100;
A = 8'h29; B = 8'h6B; #100;
A = 8'h29; B = 8'h6C; #100;
A = 8'h29; B = 8'h6D; #100;
A = 8'h29; B = 8'h6E; #100;
A = 8'h29; B = 8'h6F; #100;
A = 8'h29; B = 8'h70; #100;
A = 8'h29; B = 8'h71; #100;
A = 8'h29; B = 8'h72; #100;
A = 8'h29; B = 8'h73; #100;
A = 8'h29; B = 8'h74; #100;
A = 8'h29; B = 8'h75; #100;
A = 8'h29; B = 8'h76; #100;
A = 8'h29; B = 8'h77; #100;
A = 8'h29; B = 8'h78; #100;
A = 8'h29; B = 8'h79; #100;
A = 8'h29; B = 8'h7A; #100;
A = 8'h29; B = 8'h7B; #100;
A = 8'h29; B = 8'h7C; #100;
A = 8'h29; B = 8'h7D; #100;
A = 8'h29; B = 8'h7E; #100;
A = 8'h29; B = 8'h7F; #100;
A = 8'h29; B = 8'h80; #100;
A = 8'h29; B = 8'h81; #100;
A = 8'h29; B = 8'h82; #100;
A = 8'h29; B = 8'h83; #100;
A = 8'h29; B = 8'h84; #100;
A = 8'h29; B = 8'h85; #100;
A = 8'h29; B = 8'h86; #100;
A = 8'h29; B = 8'h87; #100;
A = 8'h29; B = 8'h88; #100;
A = 8'h29; B = 8'h89; #100;
A = 8'h29; B = 8'h8A; #100;
A = 8'h29; B = 8'h8B; #100;
A = 8'h29; B = 8'h8C; #100;
A = 8'h29; B = 8'h8D; #100;
A = 8'h29; B = 8'h8E; #100;
A = 8'h29; B = 8'h8F; #100;
A = 8'h29; B = 8'h90; #100;
A = 8'h29; B = 8'h91; #100;
A = 8'h29; B = 8'h92; #100;
A = 8'h29; B = 8'h93; #100;
A = 8'h29; B = 8'h94; #100;
A = 8'h29; B = 8'h95; #100;
A = 8'h29; B = 8'h96; #100;
A = 8'h29; B = 8'h97; #100;
A = 8'h29; B = 8'h98; #100;
A = 8'h29; B = 8'h99; #100;
A = 8'h29; B = 8'h9A; #100;
A = 8'h29; B = 8'h9B; #100;
A = 8'h29; B = 8'h9C; #100;
A = 8'h29; B = 8'h9D; #100;
A = 8'h29; B = 8'h9E; #100;
A = 8'h29; B = 8'h9F; #100;
A = 8'h29; B = 8'hA0; #100;
A = 8'h29; B = 8'hA1; #100;
A = 8'h29; B = 8'hA2; #100;
A = 8'h29; B = 8'hA3; #100;
A = 8'h29; B = 8'hA4; #100;
A = 8'h29; B = 8'hA5; #100;
A = 8'h29; B = 8'hA6; #100;
A = 8'h29; B = 8'hA7; #100;
A = 8'h29; B = 8'hA8; #100;
A = 8'h29; B = 8'hA9; #100;
A = 8'h29; B = 8'hAA; #100;
A = 8'h29; B = 8'hAB; #100;
A = 8'h29; B = 8'hAC; #100;
A = 8'h29; B = 8'hAD; #100;
A = 8'h29; B = 8'hAE; #100;
A = 8'h29; B = 8'hAF; #100;
A = 8'h29; B = 8'hB0; #100;
A = 8'h29; B = 8'hB1; #100;
A = 8'h29; B = 8'hB2; #100;
A = 8'h29; B = 8'hB3; #100;
A = 8'h29; B = 8'hB4; #100;
A = 8'h29; B = 8'hB5; #100;
A = 8'h29; B = 8'hB6; #100;
A = 8'h29; B = 8'hB7; #100;
A = 8'h29; B = 8'hB8; #100;
A = 8'h29; B = 8'hB9; #100;
A = 8'h29; B = 8'hBA; #100;
A = 8'h29; B = 8'hBB; #100;
A = 8'h29; B = 8'hBC; #100;
A = 8'h29; B = 8'hBD; #100;
A = 8'h29; B = 8'hBE; #100;
A = 8'h29; B = 8'hBF; #100;
A = 8'h29; B = 8'hC0; #100;
A = 8'h29; B = 8'hC1; #100;
A = 8'h29; B = 8'hC2; #100;
A = 8'h29; B = 8'hC3; #100;
A = 8'h29; B = 8'hC4; #100;
A = 8'h29; B = 8'hC5; #100;
A = 8'h29; B = 8'hC6; #100;
A = 8'h29; B = 8'hC7; #100;
A = 8'h29; B = 8'hC8; #100;
A = 8'h29; B = 8'hC9; #100;
A = 8'h29; B = 8'hCA; #100;
A = 8'h29; B = 8'hCB; #100;
A = 8'h29; B = 8'hCC; #100;
A = 8'h29; B = 8'hCD; #100;
A = 8'h29; B = 8'hCE; #100;
A = 8'h29; B = 8'hCF; #100;
A = 8'h29; B = 8'hD0; #100;
A = 8'h29; B = 8'hD1; #100;
A = 8'h29; B = 8'hD2; #100;
A = 8'h29; B = 8'hD3; #100;
A = 8'h29; B = 8'hD4; #100;
A = 8'h29; B = 8'hD5; #100;
A = 8'h29; B = 8'hD6; #100;
A = 8'h29; B = 8'hD7; #100;
A = 8'h29; B = 8'hD8; #100;
A = 8'h29; B = 8'hD9; #100;
A = 8'h29; B = 8'hDA; #100;
A = 8'h29; B = 8'hDB; #100;
A = 8'h29; B = 8'hDC; #100;
A = 8'h29; B = 8'hDD; #100;
A = 8'h29; B = 8'hDE; #100;
A = 8'h29; B = 8'hDF; #100;
A = 8'h29; B = 8'hE0; #100;
A = 8'h29; B = 8'hE1; #100;
A = 8'h29; B = 8'hE2; #100;
A = 8'h29; B = 8'hE3; #100;
A = 8'h29; B = 8'hE4; #100;
A = 8'h29; B = 8'hE5; #100;
A = 8'h29; B = 8'hE6; #100;
A = 8'h29; B = 8'hE7; #100;
A = 8'h29; B = 8'hE8; #100;
A = 8'h29; B = 8'hE9; #100;
A = 8'h29; B = 8'hEA; #100;
A = 8'h29; B = 8'hEB; #100;
A = 8'h29; B = 8'hEC; #100;
A = 8'h29; B = 8'hED; #100;
A = 8'h29; B = 8'hEE; #100;
A = 8'h29; B = 8'hEF; #100;
A = 8'h29; B = 8'hF0; #100;
A = 8'h29; B = 8'hF1; #100;
A = 8'h29; B = 8'hF2; #100;
A = 8'h29; B = 8'hF3; #100;
A = 8'h29; B = 8'hF4; #100;
A = 8'h29; B = 8'hF5; #100;
A = 8'h29; B = 8'hF6; #100;
A = 8'h29; B = 8'hF7; #100;
A = 8'h29; B = 8'hF8; #100;
A = 8'h29; B = 8'hF9; #100;
A = 8'h29; B = 8'hFA; #100;
A = 8'h29; B = 8'hFB; #100;
A = 8'h29; B = 8'hFC; #100;
A = 8'h29; B = 8'hFD; #100;
A = 8'h29; B = 8'hFE; #100;
A = 8'h29; B = 8'hFF; #100;
A = 8'h2A; B = 8'h0; #100;
A = 8'h2A; B = 8'h1; #100;
A = 8'h2A; B = 8'h2; #100;
A = 8'h2A; B = 8'h3; #100;
A = 8'h2A; B = 8'h4; #100;
A = 8'h2A; B = 8'h5; #100;
A = 8'h2A; B = 8'h6; #100;
A = 8'h2A; B = 8'h7; #100;
A = 8'h2A; B = 8'h8; #100;
A = 8'h2A; B = 8'h9; #100;
A = 8'h2A; B = 8'hA; #100;
A = 8'h2A; B = 8'hB; #100;
A = 8'h2A; B = 8'hC; #100;
A = 8'h2A; B = 8'hD; #100;
A = 8'h2A; B = 8'hE; #100;
A = 8'h2A; B = 8'hF; #100;
A = 8'h2A; B = 8'h10; #100;
A = 8'h2A; B = 8'h11; #100;
A = 8'h2A; B = 8'h12; #100;
A = 8'h2A; B = 8'h13; #100;
A = 8'h2A; B = 8'h14; #100;
A = 8'h2A; B = 8'h15; #100;
A = 8'h2A; B = 8'h16; #100;
A = 8'h2A; B = 8'h17; #100;
A = 8'h2A; B = 8'h18; #100;
A = 8'h2A; B = 8'h19; #100;
A = 8'h2A; B = 8'h1A; #100;
A = 8'h2A; B = 8'h1B; #100;
A = 8'h2A; B = 8'h1C; #100;
A = 8'h2A; B = 8'h1D; #100;
A = 8'h2A; B = 8'h1E; #100;
A = 8'h2A; B = 8'h1F; #100;
A = 8'h2A; B = 8'h20; #100;
A = 8'h2A; B = 8'h21; #100;
A = 8'h2A; B = 8'h22; #100;
A = 8'h2A; B = 8'h23; #100;
A = 8'h2A; B = 8'h24; #100;
A = 8'h2A; B = 8'h25; #100;
A = 8'h2A; B = 8'h26; #100;
A = 8'h2A; B = 8'h27; #100;
A = 8'h2A; B = 8'h28; #100;
A = 8'h2A; B = 8'h29; #100;
A = 8'h2A; B = 8'h2A; #100;
A = 8'h2A; B = 8'h2B; #100;
A = 8'h2A; B = 8'h2C; #100;
A = 8'h2A; B = 8'h2D; #100;
A = 8'h2A; B = 8'h2E; #100;
A = 8'h2A; B = 8'h2F; #100;
A = 8'h2A; B = 8'h30; #100;
A = 8'h2A; B = 8'h31; #100;
A = 8'h2A; B = 8'h32; #100;
A = 8'h2A; B = 8'h33; #100;
A = 8'h2A; B = 8'h34; #100;
A = 8'h2A; B = 8'h35; #100;
A = 8'h2A; B = 8'h36; #100;
A = 8'h2A; B = 8'h37; #100;
A = 8'h2A; B = 8'h38; #100;
A = 8'h2A; B = 8'h39; #100;
A = 8'h2A; B = 8'h3A; #100;
A = 8'h2A; B = 8'h3B; #100;
A = 8'h2A; B = 8'h3C; #100;
A = 8'h2A; B = 8'h3D; #100;
A = 8'h2A; B = 8'h3E; #100;
A = 8'h2A; B = 8'h3F; #100;
A = 8'h2A; B = 8'h40; #100;
A = 8'h2A; B = 8'h41; #100;
A = 8'h2A; B = 8'h42; #100;
A = 8'h2A; B = 8'h43; #100;
A = 8'h2A; B = 8'h44; #100;
A = 8'h2A; B = 8'h45; #100;
A = 8'h2A; B = 8'h46; #100;
A = 8'h2A; B = 8'h47; #100;
A = 8'h2A; B = 8'h48; #100;
A = 8'h2A; B = 8'h49; #100;
A = 8'h2A; B = 8'h4A; #100;
A = 8'h2A; B = 8'h4B; #100;
A = 8'h2A; B = 8'h4C; #100;
A = 8'h2A; B = 8'h4D; #100;
A = 8'h2A; B = 8'h4E; #100;
A = 8'h2A; B = 8'h4F; #100;
A = 8'h2A; B = 8'h50; #100;
A = 8'h2A; B = 8'h51; #100;
A = 8'h2A; B = 8'h52; #100;
A = 8'h2A; B = 8'h53; #100;
A = 8'h2A; B = 8'h54; #100;
A = 8'h2A; B = 8'h55; #100;
A = 8'h2A; B = 8'h56; #100;
A = 8'h2A; B = 8'h57; #100;
A = 8'h2A; B = 8'h58; #100;
A = 8'h2A; B = 8'h59; #100;
A = 8'h2A; B = 8'h5A; #100;
A = 8'h2A; B = 8'h5B; #100;
A = 8'h2A; B = 8'h5C; #100;
A = 8'h2A; B = 8'h5D; #100;
A = 8'h2A; B = 8'h5E; #100;
A = 8'h2A; B = 8'h5F; #100;
A = 8'h2A; B = 8'h60; #100;
A = 8'h2A; B = 8'h61; #100;
A = 8'h2A; B = 8'h62; #100;
A = 8'h2A; B = 8'h63; #100;
A = 8'h2A; B = 8'h64; #100;
A = 8'h2A; B = 8'h65; #100;
A = 8'h2A; B = 8'h66; #100;
A = 8'h2A; B = 8'h67; #100;
A = 8'h2A; B = 8'h68; #100;
A = 8'h2A; B = 8'h69; #100;
A = 8'h2A; B = 8'h6A; #100;
A = 8'h2A; B = 8'h6B; #100;
A = 8'h2A; B = 8'h6C; #100;
A = 8'h2A; B = 8'h6D; #100;
A = 8'h2A; B = 8'h6E; #100;
A = 8'h2A; B = 8'h6F; #100;
A = 8'h2A; B = 8'h70; #100;
A = 8'h2A; B = 8'h71; #100;
A = 8'h2A; B = 8'h72; #100;
A = 8'h2A; B = 8'h73; #100;
A = 8'h2A; B = 8'h74; #100;
A = 8'h2A; B = 8'h75; #100;
A = 8'h2A; B = 8'h76; #100;
A = 8'h2A; B = 8'h77; #100;
A = 8'h2A; B = 8'h78; #100;
A = 8'h2A; B = 8'h79; #100;
A = 8'h2A; B = 8'h7A; #100;
A = 8'h2A; B = 8'h7B; #100;
A = 8'h2A; B = 8'h7C; #100;
A = 8'h2A; B = 8'h7D; #100;
A = 8'h2A; B = 8'h7E; #100;
A = 8'h2A; B = 8'h7F; #100;
A = 8'h2A; B = 8'h80; #100;
A = 8'h2A; B = 8'h81; #100;
A = 8'h2A; B = 8'h82; #100;
A = 8'h2A; B = 8'h83; #100;
A = 8'h2A; B = 8'h84; #100;
A = 8'h2A; B = 8'h85; #100;
A = 8'h2A; B = 8'h86; #100;
A = 8'h2A; B = 8'h87; #100;
A = 8'h2A; B = 8'h88; #100;
A = 8'h2A; B = 8'h89; #100;
A = 8'h2A; B = 8'h8A; #100;
A = 8'h2A; B = 8'h8B; #100;
A = 8'h2A; B = 8'h8C; #100;
A = 8'h2A; B = 8'h8D; #100;
A = 8'h2A; B = 8'h8E; #100;
A = 8'h2A; B = 8'h8F; #100;
A = 8'h2A; B = 8'h90; #100;
A = 8'h2A; B = 8'h91; #100;
A = 8'h2A; B = 8'h92; #100;
A = 8'h2A; B = 8'h93; #100;
A = 8'h2A; B = 8'h94; #100;
A = 8'h2A; B = 8'h95; #100;
A = 8'h2A; B = 8'h96; #100;
A = 8'h2A; B = 8'h97; #100;
A = 8'h2A; B = 8'h98; #100;
A = 8'h2A; B = 8'h99; #100;
A = 8'h2A; B = 8'h9A; #100;
A = 8'h2A; B = 8'h9B; #100;
A = 8'h2A; B = 8'h9C; #100;
A = 8'h2A; B = 8'h9D; #100;
A = 8'h2A; B = 8'h9E; #100;
A = 8'h2A; B = 8'h9F; #100;
A = 8'h2A; B = 8'hA0; #100;
A = 8'h2A; B = 8'hA1; #100;
A = 8'h2A; B = 8'hA2; #100;
A = 8'h2A; B = 8'hA3; #100;
A = 8'h2A; B = 8'hA4; #100;
A = 8'h2A; B = 8'hA5; #100;
A = 8'h2A; B = 8'hA6; #100;
A = 8'h2A; B = 8'hA7; #100;
A = 8'h2A; B = 8'hA8; #100;
A = 8'h2A; B = 8'hA9; #100;
A = 8'h2A; B = 8'hAA; #100;
A = 8'h2A; B = 8'hAB; #100;
A = 8'h2A; B = 8'hAC; #100;
A = 8'h2A; B = 8'hAD; #100;
A = 8'h2A; B = 8'hAE; #100;
A = 8'h2A; B = 8'hAF; #100;
A = 8'h2A; B = 8'hB0; #100;
A = 8'h2A; B = 8'hB1; #100;
A = 8'h2A; B = 8'hB2; #100;
A = 8'h2A; B = 8'hB3; #100;
A = 8'h2A; B = 8'hB4; #100;
A = 8'h2A; B = 8'hB5; #100;
A = 8'h2A; B = 8'hB6; #100;
A = 8'h2A; B = 8'hB7; #100;
A = 8'h2A; B = 8'hB8; #100;
A = 8'h2A; B = 8'hB9; #100;
A = 8'h2A; B = 8'hBA; #100;
A = 8'h2A; B = 8'hBB; #100;
A = 8'h2A; B = 8'hBC; #100;
A = 8'h2A; B = 8'hBD; #100;
A = 8'h2A; B = 8'hBE; #100;
A = 8'h2A; B = 8'hBF; #100;
A = 8'h2A; B = 8'hC0; #100;
A = 8'h2A; B = 8'hC1; #100;
A = 8'h2A; B = 8'hC2; #100;
A = 8'h2A; B = 8'hC3; #100;
A = 8'h2A; B = 8'hC4; #100;
A = 8'h2A; B = 8'hC5; #100;
A = 8'h2A; B = 8'hC6; #100;
A = 8'h2A; B = 8'hC7; #100;
A = 8'h2A; B = 8'hC8; #100;
A = 8'h2A; B = 8'hC9; #100;
A = 8'h2A; B = 8'hCA; #100;
A = 8'h2A; B = 8'hCB; #100;
A = 8'h2A; B = 8'hCC; #100;
A = 8'h2A; B = 8'hCD; #100;
A = 8'h2A; B = 8'hCE; #100;
A = 8'h2A; B = 8'hCF; #100;
A = 8'h2A; B = 8'hD0; #100;
A = 8'h2A; B = 8'hD1; #100;
A = 8'h2A; B = 8'hD2; #100;
A = 8'h2A; B = 8'hD3; #100;
A = 8'h2A; B = 8'hD4; #100;
A = 8'h2A; B = 8'hD5; #100;
A = 8'h2A; B = 8'hD6; #100;
A = 8'h2A; B = 8'hD7; #100;
A = 8'h2A; B = 8'hD8; #100;
A = 8'h2A; B = 8'hD9; #100;
A = 8'h2A; B = 8'hDA; #100;
A = 8'h2A; B = 8'hDB; #100;
A = 8'h2A; B = 8'hDC; #100;
A = 8'h2A; B = 8'hDD; #100;
A = 8'h2A; B = 8'hDE; #100;
A = 8'h2A; B = 8'hDF; #100;
A = 8'h2A; B = 8'hE0; #100;
A = 8'h2A; B = 8'hE1; #100;
A = 8'h2A; B = 8'hE2; #100;
A = 8'h2A; B = 8'hE3; #100;
A = 8'h2A; B = 8'hE4; #100;
A = 8'h2A; B = 8'hE5; #100;
A = 8'h2A; B = 8'hE6; #100;
A = 8'h2A; B = 8'hE7; #100;
A = 8'h2A; B = 8'hE8; #100;
A = 8'h2A; B = 8'hE9; #100;
A = 8'h2A; B = 8'hEA; #100;
A = 8'h2A; B = 8'hEB; #100;
A = 8'h2A; B = 8'hEC; #100;
A = 8'h2A; B = 8'hED; #100;
A = 8'h2A; B = 8'hEE; #100;
A = 8'h2A; B = 8'hEF; #100;
A = 8'h2A; B = 8'hF0; #100;
A = 8'h2A; B = 8'hF1; #100;
A = 8'h2A; B = 8'hF2; #100;
A = 8'h2A; B = 8'hF3; #100;
A = 8'h2A; B = 8'hF4; #100;
A = 8'h2A; B = 8'hF5; #100;
A = 8'h2A; B = 8'hF6; #100;
A = 8'h2A; B = 8'hF7; #100;
A = 8'h2A; B = 8'hF8; #100;
A = 8'h2A; B = 8'hF9; #100;
A = 8'h2A; B = 8'hFA; #100;
A = 8'h2A; B = 8'hFB; #100;
A = 8'h2A; B = 8'hFC; #100;
A = 8'h2A; B = 8'hFD; #100;
A = 8'h2A; B = 8'hFE; #100;
A = 8'h2A; B = 8'hFF; #100;
A = 8'h2B; B = 8'h0; #100;
A = 8'h2B; B = 8'h1; #100;
A = 8'h2B; B = 8'h2; #100;
A = 8'h2B; B = 8'h3; #100;
A = 8'h2B; B = 8'h4; #100;
A = 8'h2B; B = 8'h5; #100;
A = 8'h2B; B = 8'h6; #100;
A = 8'h2B; B = 8'h7; #100;
A = 8'h2B; B = 8'h8; #100;
A = 8'h2B; B = 8'h9; #100;
A = 8'h2B; B = 8'hA; #100;
A = 8'h2B; B = 8'hB; #100;
A = 8'h2B; B = 8'hC; #100;
A = 8'h2B; B = 8'hD; #100;
A = 8'h2B; B = 8'hE; #100;
A = 8'h2B; B = 8'hF; #100;
A = 8'h2B; B = 8'h10; #100;
A = 8'h2B; B = 8'h11; #100;
A = 8'h2B; B = 8'h12; #100;
A = 8'h2B; B = 8'h13; #100;
A = 8'h2B; B = 8'h14; #100;
A = 8'h2B; B = 8'h15; #100;
A = 8'h2B; B = 8'h16; #100;
A = 8'h2B; B = 8'h17; #100;
A = 8'h2B; B = 8'h18; #100;
A = 8'h2B; B = 8'h19; #100;
A = 8'h2B; B = 8'h1A; #100;
A = 8'h2B; B = 8'h1B; #100;
A = 8'h2B; B = 8'h1C; #100;
A = 8'h2B; B = 8'h1D; #100;
A = 8'h2B; B = 8'h1E; #100;
A = 8'h2B; B = 8'h1F; #100;
A = 8'h2B; B = 8'h20; #100;
A = 8'h2B; B = 8'h21; #100;
A = 8'h2B; B = 8'h22; #100;
A = 8'h2B; B = 8'h23; #100;
A = 8'h2B; B = 8'h24; #100;
A = 8'h2B; B = 8'h25; #100;
A = 8'h2B; B = 8'h26; #100;
A = 8'h2B; B = 8'h27; #100;
A = 8'h2B; B = 8'h28; #100;
A = 8'h2B; B = 8'h29; #100;
A = 8'h2B; B = 8'h2A; #100;
A = 8'h2B; B = 8'h2B; #100;
A = 8'h2B; B = 8'h2C; #100;
A = 8'h2B; B = 8'h2D; #100;
A = 8'h2B; B = 8'h2E; #100;
A = 8'h2B; B = 8'h2F; #100;
A = 8'h2B; B = 8'h30; #100;
A = 8'h2B; B = 8'h31; #100;
A = 8'h2B; B = 8'h32; #100;
A = 8'h2B; B = 8'h33; #100;
A = 8'h2B; B = 8'h34; #100;
A = 8'h2B; B = 8'h35; #100;
A = 8'h2B; B = 8'h36; #100;
A = 8'h2B; B = 8'h37; #100;
A = 8'h2B; B = 8'h38; #100;
A = 8'h2B; B = 8'h39; #100;
A = 8'h2B; B = 8'h3A; #100;
A = 8'h2B; B = 8'h3B; #100;
A = 8'h2B; B = 8'h3C; #100;
A = 8'h2B; B = 8'h3D; #100;
A = 8'h2B; B = 8'h3E; #100;
A = 8'h2B; B = 8'h3F; #100;
A = 8'h2B; B = 8'h40; #100;
A = 8'h2B; B = 8'h41; #100;
A = 8'h2B; B = 8'h42; #100;
A = 8'h2B; B = 8'h43; #100;
A = 8'h2B; B = 8'h44; #100;
A = 8'h2B; B = 8'h45; #100;
A = 8'h2B; B = 8'h46; #100;
A = 8'h2B; B = 8'h47; #100;
A = 8'h2B; B = 8'h48; #100;
A = 8'h2B; B = 8'h49; #100;
A = 8'h2B; B = 8'h4A; #100;
A = 8'h2B; B = 8'h4B; #100;
A = 8'h2B; B = 8'h4C; #100;
A = 8'h2B; B = 8'h4D; #100;
A = 8'h2B; B = 8'h4E; #100;
A = 8'h2B; B = 8'h4F; #100;
A = 8'h2B; B = 8'h50; #100;
A = 8'h2B; B = 8'h51; #100;
A = 8'h2B; B = 8'h52; #100;
A = 8'h2B; B = 8'h53; #100;
A = 8'h2B; B = 8'h54; #100;
A = 8'h2B; B = 8'h55; #100;
A = 8'h2B; B = 8'h56; #100;
A = 8'h2B; B = 8'h57; #100;
A = 8'h2B; B = 8'h58; #100;
A = 8'h2B; B = 8'h59; #100;
A = 8'h2B; B = 8'h5A; #100;
A = 8'h2B; B = 8'h5B; #100;
A = 8'h2B; B = 8'h5C; #100;
A = 8'h2B; B = 8'h5D; #100;
A = 8'h2B; B = 8'h5E; #100;
A = 8'h2B; B = 8'h5F; #100;
A = 8'h2B; B = 8'h60; #100;
A = 8'h2B; B = 8'h61; #100;
A = 8'h2B; B = 8'h62; #100;
A = 8'h2B; B = 8'h63; #100;
A = 8'h2B; B = 8'h64; #100;
A = 8'h2B; B = 8'h65; #100;
A = 8'h2B; B = 8'h66; #100;
A = 8'h2B; B = 8'h67; #100;
A = 8'h2B; B = 8'h68; #100;
A = 8'h2B; B = 8'h69; #100;
A = 8'h2B; B = 8'h6A; #100;
A = 8'h2B; B = 8'h6B; #100;
A = 8'h2B; B = 8'h6C; #100;
A = 8'h2B; B = 8'h6D; #100;
A = 8'h2B; B = 8'h6E; #100;
A = 8'h2B; B = 8'h6F; #100;
A = 8'h2B; B = 8'h70; #100;
A = 8'h2B; B = 8'h71; #100;
A = 8'h2B; B = 8'h72; #100;
A = 8'h2B; B = 8'h73; #100;
A = 8'h2B; B = 8'h74; #100;
A = 8'h2B; B = 8'h75; #100;
A = 8'h2B; B = 8'h76; #100;
A = 8'h2B; B = 8'h77; #100;
A = 8'h2B; B = 8'h78; #100;
A = 8'h2B; B = 8'h79; #100;
A = 8'h2B; B = 8'h7A; #100;
A = 8'h2B; B = 8'h7B; #100;
A = 8'h2B; B = 8'h7C; #100;
A = 8'h2B; B = 8'h7D; #100;
A = 8'h2B; B = 8'h7E; #100;
A = 8'h2B; B = 8'h7F; #100;
A = 8'h2B; B = 8'h80; #100;
A = 8'h2B; B = 8'h81; #100;
A = 8'h2B; B = 8'h82; #100;
A = 8'h2B; B = 8'h83; #100;
A = 8'h2B; B = 8'h84; #100;
A = 8'h2B; B = 8'h85; #100;
A = 8'h2B; B = 8'h86; #100;
A = 8'h2B; B = 8'h87; #100;
A = 8'h2B; B = 8'h88; #100;
A = 8'h2B; B = 8'h89; #100;
A = 8'h2B; B = 8'h8A; #100;
A = 8'h2B; B = 8'h8B; #100;
A = 8'h2B; B = 8'h8C; #100;
A = 8'h2B; B = 8'h8D; #100;
A = 8'h2B; B = 8'h8E; #100;
A = 8'h2B; B = 8'h8F; #100;
A = 8'h2B; B = 8'h90; #100;
A = 8'h2B; B = 8'h91; #100;
A = 8'h2B; B = 8'h92; #100;
A = 8'h2B; B = 8'h93; #100;
A = 8'h2B; B = 8'h94; #100;
A = 8'h2B; B = 8'h95; #100;
A = 8'h2B; B = 8'h96; #100;
A = 8'h2B; B = 8'h97; #100;
A = 8'h2B; B = 8'h98; #100;
A = 8'h2B; B = 8'h99; #100;
A = 8'h2B; B = 8'h9A; #100;
A = 8'h2B; B = 8'h9B; #100;
A = 8'h2B; B = 8'h9C; #100;
A = 8'h2B; B = 8'h9D; #100;
A = 8'h2B; B = 8'h9E; #100;
A = 8'h2B; B = 8'h9F; #100;
A = 8'h2B; B = 8'hA0; #100;
A = 8'h2B; B = 8'hA1; #100;
A = 8'h2B; B = 8'hA2; #100;
A = 8'h2B; B = 8'hA3; #100;
A = 8'h2B; B = 8'hA4; #100;
A = 8'h2B; B = 8'hA5; #100;
A = 8'h2B; B = 8'hA6; #100;
A = 8'h2B; B = 8'hA7; #100;
A = 8'h2B; B = 8'hA8; #100;
A = 8'h2B; B = 8'hA9; #100;
A = 8'h2B; B = 8'hAA; #100;
A = 8'h2B; B = 8'hAB; #100;
A = 8'h2B; B = 8'hAC; #100;
A = 8'h2B; B = 8'hAD; #100;
A = 8'h2B; B = 8'hAE; #100;
A = 8'h2B; B = 8'hAF; #100;
A = 8'h2B; B = 8'hB0; #100;
A = 8'h2B; B = 8'hB1; #100;
A = 8'h2B; B = 8'hB2; #100;
A = 8'h2B; B = 8'hB3; #100;
A = 8'h2B; B = 8'hB4; #100;
A = 8'h2B; B = 8'hB5; #100;
A = 8'h2B; B = 8'hB6; #100;
A = 8'h2B; B = 8'hB7; #100;
A = 8'h2B; B = 8'hB8; #100;
A = 8'h2B; B = 8'hB9; #100;
A = 8'h2B; B = 8'hBA; #100;
A = 8'h2B; B = 8'hBB; #100;
A = 8'h2B; B = 8'hBC; #100;
A = 8'h2B; B = 8'hBD; #100;
A = 8'h2B; B = 8'hBE; #100;
A = 8'h2B; B = 8'hBF; #100;
A = 8'h2B; B = 8'hC0; #100;
A = 8'h2B; B = 8'hC1; #100;
A = 8'h2B; B = 8'hC2; #100;
A = 8'h2B; B = 8'hC3; #100;
A = 8'h2B; B = 8'hC4; #100;
A = 8'h2B; B = 8'hC5; #100;
A = 8'h2B; B = 8'hC6; #100;
A = 8'h2B; B = 8'hC7; #100;
A = 8'h2B; B = 8'hC8; #100;
A = 8'h2B; B = 8'hC9; #100;
A = 8'h2B; B = 8'hCA; #100;
A = 8'h2B; B = 8'hCB; #100;
A = 8'h2B; B = 8'hCC; #100;
A = 8'h2B; B = 8'hCD; #100;
A = 8'h2B; B = 8'hCE; #100;
A = 8'h2B; B = 8'hCF; #100;
A = 8'h2B; B = 8'hD0; #100;
A = 8'h2B; B = 8'hD1; #100;
A = 8'h2B; B = 8'hD2; #100;
A = 8'h2B; B = 8'hD3; #100;
A = 8'h2B; B = 8'hD4; #100;
A = 8'h2B; B = 8'hD5; #100;
A = 8'h2B; B = 8'hD6; #100;
A = 8'h2B; B = 8'hD7; #100;
A = 8'h2B; B = 8'hD8; #100;
A = 8'h2B; B = 8'hD9; #100;
A = 8'h2B; B = 8'hDA; #100;
A = 8'h2B; B = 8'hDB; #100;
A = 8'h2B; B = 8'hDC; #100;
A = 8'h2B; B = 8'hDD; #100;
A = 8'h2B; B = 8'hDE; #100;
A = 8'h2B; B = 8'hDF; #100;
A = 8'h2B; B = 8'hE0; #100;
A = 8'h2B; B = 8'hE1; #100;
A = 8'h2B; B = 8'hE2; #100;
A = 8'h2B; B = 8'hE3; #100;
A = 8'h2B; B = 8'hE4; #100;
A = 8'h2B; B = 8'hE5; #100;
A = 8'h2B; B = 8'hE6; #100;
A = 8'h2B; B = 8'hE7; #100;
A = 8'h2B; B = 8'hE8; #100;
A = 8'h2B; B = 8'hE9; #100;
A = 8'h2B; B = 8'hEA; #100;
A = 8'h2B; B = 8'hEB; #100;
A = 8'h2B; B = 8'hEC; #100;
A = 8'h2B; B = 8'hED; #100;
A = 8'h2B; B = 8'hEE; #100;
A = 8'h2B; B = 8'hEF; #100;
A = 8'h2B; B = 8'hF0; #100;
A = 8'h2B; B = 8'hF1; #100;
A = 8'h2B; B = 8'hF2; #100;
A = 8'h2B; B = 8'hF3; #100;
A = 8'h2B; B = 8'hF4; #100;
A = 8'h2B; B = 8'hF5; #100;
A = 8'h2B; B = 8'hF6; #100;
A = 8'h2B; B = 8'hF7; #100;
A = 8'h2B; B = 8'hF8; #100;
A = 8'h2B; B = 8'hF9; #100;
A = 8'h2B; B = 8'hFA; #100;
A = 8'h2B; B = 8'hFB; #100;
A = 8'h2B; B = 8'hFC; #100;
A = 8'h2B; B = 8'hFD; #100;
A = 8'h2B; B = 8'hFE; #100;
A = 8'h2B; B = 8'hFF; #100;
A = 8'h2C; B = 8'h0; #100;
A = 8'h2C; B = 8'h1; #100;
A = 8'h2C; B = 8'h2; #100;
A = 8'h2C; B = 8'h3; #100;
A = 8'h2C; B = 8'h4; #100;
A = 8'h2C; B = 8'h5; #100;
A = 8'h2C; B = 8'h6; #100;
A = 8'h2C; B = 8'h7; #100;
A = 8'h2C; B = 8'h8; #100;
A = 8'h2C; B = 8'h9; #100;
A = 8'h2C; B = 8'hA; #100;
A = 8'h2C; B = 8'hB; #100;
A = 8'h2C; B = 8'hC; #100;
A = 8'h2C; B = 8'hD; #100;
A = 8'h2C; B = 8'hE; #100;
A = 8'h2C; B = 8'hF; #100;
A = 8'h2C; B = 8'h10; #100;
A = 8'h2C; B = 8'h11; #100;
A = 8'h2C; B = 8'h12; #100;
A = 8'h2C; B = 8'h13; #100;
A = 8'h2C; B = 8'h14; #100;
A = 8'h2C; B = 8'h15; #100;
A = 8'h2C; B = 8'h16; #100;
A = 8'h2C; B = 8'h17; #100;
A = 8'h2C; B = 8'h18; #100;
A = 8'h2C; B = 8'h19; #100;
A = 8'h2C; B = 8'h1A; #100;
A = 8'h2C; B = 8'h1B; #100;
A = 8'h2C; B = 8'h1C; #100;
A = 8'h2C; B = 8'h1D; #100;
A = 8'h2C; B = 8'h1E; #100;
A = 8'h2C; B = 8'h1F; #100;
A = 8'h2C; B = 8'h20; #100;
A = 8'h2C; B = 8'h21; #100;
A = 8'h2C; B = 8'h22; #100;
A = 8'h2C; B = 8'h23; #100;
A = 8'h2C; B = 8'h24; #100;
A = 8'h2C; B = 8'h25; #100;
A = 8'h2C; B = 8'h26; #100;
A = 8'h2C; B = 8'h27; #100;
A = 8'h2C; B = 8'h28; #100;
A = 8'h2C; B = 8'h29; #100;
A = 8'h2C; B = 8'h2A; #100;
A = 8'h2C; B = 8'h2B; #100;
A = 8'h2C; B = 8'h2C; #100;
A = 8'h2C; B = 8'h2D; #100;
A = 8'h2C; B = 8'h2E; #100;
A = 8'h2C; B = 8'h2F; #100;
A = 8'h2C; B = 8'h30; #100;
A = 8'h2C; B = 8'h31; #100;
A = 8'h2C; B = 8'h32; #100;
A = 8'h2C; B = 8'h33; #100;
A = 8'h2C; B = 8'h34; #100;
A = 8'h2C; B = 8'h35; #100;
A = 8'h2C; B = 8'h36; #100;
A = 8'h2C; B = 8'h37; #100;
A = 8'h2C; B = 8'h38; #100;
A = 8'h2C; B = 8'h39; #100;
A = 8'h2C; B = 8'h3A; #100;
A = 8'h2C; B = 8'h3B; #100;
A = 8'h2C; B = 8'h3C; #100;
A = 8'h2C; B = 8'h3D; #100;
A = 8'h2C; B = 8'h3E; #100;
A = 8'h2C; B = 8'h3F; #100;
A = 8'h2C; B = 8'h40; #100;
A = 8'h2C; B = 8'h41; #100;
A = 8'h2C; B = 8'h42; #100;
A = 8'h2C; B = 8'h43; #100;
A = 8'h2C; B = 8'h44; #100;
A = 8'h2C; B = 8'h45; #100;
A = 8'h2C; B = 8'h46; #100;
A = 8'h2C; B = 8'h47; #100;
A = 8'h2C; B = 8'h48; #100;
A = 8'h2C; B = 8'h49; #100;
A = 8'h2C; B = 8'h4A; #100;
A = 8'h2C; B = 8'h4B; #100;
A = 8'h2C; B = 8'h4C; #100;
A = 8'h2C; B = 8'h4D; #100;
A = 8'h2C; B = 8'h4E; #100;
A = 8'h2C; B = 8'h4F; #100;
A = 8'h2C; B = 8'h50; #100;
A = 8'h2C; B = 8'h51; #100;
A = 8'h2C; B = 8'h52; #100;
A = 8'h2C; B = 8'h53; #100;
A = 8'h2C; B = 8'h54; #100;
A = 8'h2C; B = 8'h55; #100;
A = 8'h2C; B = 8'h56; #100;
A = 8'h2C; B = 8'h57; #100;
A = 8'h2C; B = 8'h58; #100;
A = 8'h2C; B = 8'h59; #100;
A = 8'h2C; B = 8'h5A; #100;
A = 8'h2C; B = 8'h5B; #100;
A = 8'h2C; B = 8'h5C; #100;
A = 8'h2C; B = 8'h5D; #100;
A = 8'h2C; B = 8'h5E; #100;
A = 8'h2C; B = 8'h5F; #100;
A = 8'h2C; B = 8'h60; #100;
A = 8'h2C; B = 8'h61; #100;
A = 8'h2C; B = 8'h62; #100;
A = 8'h2C; B = 8'h63; #100;
A = 8'h2C; B = 8'h64; #100;
A = 8'h2C; B = 8'h65; #100;
A = 8'h2C; B = 8'h66; #100;
A = 8'h2C; B = 8'h67; #100;
A = 8'h2C; B = 8'h68; #100;
A = 8'h2C; B = 8'h69; #100;
A = 8'h2C; B = 8'h6A; #100;
A = 8'h2C; B = 8'h6B; #100;
A = 8'h2C; B = 8'h6C; #100;
A = 8'h2C; B = 8'h6D; #100;
A = 8'h2C; B = 8'h6E; #100;
A = 8'h2C; B = 8'h6F; #100;
A = 8'h2C; B = 8'h70; #100;
A = 8'h2C; B = 8'h71; #100;
A = 8'h2C; B = 8'h72; #100;
A = 8'h2C; B = 8'h73; #100;
A = 8'h2C; B = 8'h74; #100;
A = 8'h2C; B = 8'h75; #100;
A = 8'h2C; B = 8'h76; #100;
A = 8'h2C; B = 8'h77; #100;
A = 8'h2C; B = 8'h78; #100;
A = 8'h2C; B = 8'h79; #100;
A = 8'h2C; B = 8'h7A; #100;
A = 8'h2C; B = 8'h7B; #100;
A = 8'h2C; B = 8'h7C; #100;
A = 8'h2C; B = 8'h7D; #100;
A = 8'h2C; B = 8'h7E; #100;
A = 8'h2C; B = 8'h7F; #100;
A = 8'h2C; B = 8'h80; #100;
A = 8'h2C; B = 8'h81; #100;
A = 8'h2C; B = 8'h82; #100;
A = 8'h2C; B = 8'h83; #100;
A = 8'h2C; B = 8'h84; #100;
A = 8'h2C; B = 8'h85; #100;
A = 8'h2C; B = 8'h86; #100;
A = 8'h2C; B = 8'h87; #100;
A = 8'h2C; B = 8'h88; #100;
A = 8'h2C; B = 8'h89; #100;
A = 8'h2C; B = 8'h8A; #100;
A = 8'h2C; B = 8'h8B; #100;
A = 8'h2C; B = 8'h8C; #100;
A = 8'h2C; B = 8'h8D; #100;
A = 8'h2C; B = 8'h8E; #100;
A = 8'h2C; B = 8'h8F; #100;
A = 8'h2C; B = 8'h90; #100;
A = 8'h2C; B = 8'h91; #100;
A = 8'h2C; B = 8'h92; #100;
A = 8'h2C; B = 8'h93; #100;
A = 8'h2C; B = 8'h94; #100;
A = 8'h2C; B = 8'h95; #100;
A = 8'h2C; B = 8'h96; #100;
A = 8'h2C; B = 8'h97; #100;
A = 8'h2C; B = 8'h98; #100;
A = 8'h2C; B = 8'h99; #100;
A = 8'h2C; B = 8'h9A; #100;
A = 8'h2C; B = 8'h9B; #100;
A = 8'h2C; B = 8'h9C; #100;
A = 8'h2C; B = 8'h9D; #100;
A = 8'h2C; B = 8'h9E; #100;
A = 8'h2C; B = 8'h9F; #100;
A = 8'h2C; B = 8'hA0; #100;
A = 8'h2C; B = 8'hA1; #100;
A = 8'h2C; B = 8'hA2; #100;
A = 8'h2C; B = 8'hA3; #100;
A = 8'h2C; B = 8'hA4; #100;
A = 8'h2C; B = 8'hA5; #100;
A = 8'h2C; B = 8'hA6; #100;
A = 8'h2C; B = 8'hA7; #100;
A = 8'h2C; B = 8'hA8; #100;
A = 8'h2C; B = 8'hA9; #100;
A = 8'h2C; B = 8'hAA; #100;
A = 8'h2C; B = 8'hAB; #100;
A = 8'h2C; B = 8'hAC; #100;
A = 8'h2C; B = 8'hAD; #100;
A = 8'h2C; B = 8'hAE; #100;
A = 8'h2C; B = 8'hAF; #100;
A = 8'h2C; B = 8'hB0; #100;
A = 8'h2C; B = 8'hB1; #100;
A = 8'h2C; B = 8'hB2; #100;
A = 8'h2C; B = 8'hB3; #100;
A = 8'h2C; B = 8'hB4; #100;
A = 8'h2C; B = 8'hB5; #100;
A = 8'h2C; B = 8'hB6; #100;
A = 8'h2C; B = 8'hB7; #100;
A = 8'h2C; B = 8'hB8; #100;
A = 8'h2C; B = 8'hB9; #100;
A = 8'h2C; B = 8'hBA; #100;
A = 8'h2C; B = 8'hBB; #100;
A = 8'h2C; B = 8'hBC; #100;
A = 8'h2C; B = 8'hBD; #100;
A = 8'h2C; B = 8'hBE; #100;
A = 8'h2C; B = 8'hBF; #100;
A = 8'h2C; B = 8'hC0; #100;
A = 8'h2C; B = 8'hC1; #100;
A = 8'h2C; B = 8'hC2; #100;
A = 8'h2C; B = 8'hC3; #100;
A = 8'h2C; B = 8'hC4; #100;
A = 8'h2C; B = 8'hC5; #100;
A = 8'h2C; B = 8'hC6; #100;
A = 8'h2C; B = 8'hC7; #100;
A = 8'h2C; B = 8'hC8; #100;
A = 8'h2C; B = 8'hC9; #100;
A = 8'h2C; B = 8'hCA; #100;
A = 8'h2C; B = 8'hCB; #100;
A = 8'h2C; B = 8'hCC; #100;
A = 8'h2C; B = 8'hCD; #100;
A = 8'h2C; B = 8'hCE; #100;
A = 8'h2C; B = 8'hCF; #100;
A = 8'h2C; B = 8'hD0; #100;
A = 8'h2C; B = 8'hD1; #100;
A = 8'h2C; B = 8'hD2; #100;
A = 8'h2C; B = 8'hD3; #100;
A = 8'h2C; B = 8'hD4; #100;
A = 8'h2C; B = 8'hD5; #100;
A = 8'h2C; B = 8'hD6; #100;
A = 8'h2C; B = 8'hD7; #100;
A = 8'h2C; B = 8'hD8; #100;
A = 8'h2C; B = 8'hD9; #100;
A = 8'h2C; B = 8'hDA; #100;
A = 8'h2C; B = 8'hDB; #100;
A = 8'h2C; B = 8'hDC; #100;
A = 8'h2C; B = 8'hDD; #100;
A = 8'h2C; B = 8'hDE; #100;
A = 8'h2C; B = 8'hDF; #100;
A = 8'h2C; B = 8'hE0; #100;
A = 8'h2C; B = 8'hE1; #100;
A = 8'h2C; B = 8'hE2; #100;
A = 8'h2C; B = 8'hE3; #100;
A = 8'h2C; B = 8'hE4; #100;
A = 8'h2C; B = 8'hE5; #100;
A = 8'h2C; B = 8'hE6; #100;
A = 8'h2C; B = 8'hE7; #100;
A = 8'h2C; B = 8'hE8; #100;
A = 8'h2C; B = 8'hE9; #100;
A = 8'h2C; B = 8'hEA; #100;
A = 8'h2C; B = 8'hEB; #100;
A = 8'h2C; B = 8'hEC; #100;
A = 8'h2C; B = 8'hED; #100;
A = 8'h2C; B = 8'hEE; #100;
A = 8'h2C; B = 8'hEF; #100;
A = 8'h2C; B = 8'hF0; #100;
A = 8'h2C; B = 8'hF1; #100;
A = 8'h2C; B = 8'hF2; #100;
A = 8'h2C; B = 8'hF3; #100;
A = 8'h2C; B = 8'hF4; #100;
A = 8'h2C; B = 8'hF5; #100;
A = 8'h2C; B = 8'hF6; #100;
A = 8'h2C; B = 8'hF7; #100;
A = 8'h2C; B = 8'hF8; #100;
A = 8'h2C; B = 8'hF9; #100;
A = 8'h2C; B = 8'hFA; #100;
A = 8'h2C; B = 8'hFB; #100;
A = 8'h2C; B = 8'hFC; #100;
A = 8'h2C; B = 8'hFD; #100;
A = 8'h2C; B = 8'hFE; #100;
A = 8'h2C; B = 8'hFF; #100;
A = 8'h2D; B = 8'h0; #100;
A = 8'h2D; B = 8'h1; #100;
A = 8'h2D; B = 8'h2; #100;
A = 8'h2D; B = 8'h3; #100;
A = 8'h2D; B = 8'h4; #100;
A = 8'h2D; B = 8'h5; #100;
A = 8'h2D; B = 8'h6; #100;
A = 8'h2D; B = 8'h7; #100;
A = 8'h2D; B = 8'h8; #100;
A = 8'h2D; B = 8'h9; #100;
A = 8'h2D; B = 8'hA; #100;
A = 8'h2D; B = 8'hB; #100;
A = 8'h2D; B = 8'hC; #100;
A = 8'h2D; B = 8'hD; #100;
A = 8'h2D; B = 8'hE; #100;
A = 8'h2D; B = 8'hF; #100;
A = 8'h2D; B = 8'h10; #100;
A = 8'h2D; B = 8'h11; #100;
A = 8'h2D; B = 8'h12; #100;
A = 8'h2D; B = 8'h13; #100;
A = 8'h2D; B = 8'h14; #100;
A = 8'h2D; B = 8'h15; #100;
A = 8'h2D; B = 8'h16; #100;
A = 8'h2D; B = 8'h17; #100;
A = 8'h2D; B = 8'h18; #100;
A = 8'h2D; B = 8'h19; #100;
A = 8'h2D; B = 8'h1A; #100;
A = 8'h2D; B = 8'h1B; #100;
A = 8'h2D; B = 8'h1C; #100;
A = 8'h2D; B = 8'h1D; #100;
A = 8'h2D; B = 8'h1E; #100;
A = 8'h2D; B = 8'h1F; #100;
A = 8'h2D; B = 8'h20; #100;
A = 8'h2D; B = 8'h21; #100;
A = 8'h2D; B = 8'h22; #100;
A = 8'h2D; B = 8'h23; #100;
A = 8'h2D; B = 8'h24; #100;
A = 8'h2D; B = 8'h25; #100;
A = 8'h2D; B = 8'h26; #100;
A = 8'h2D; B = 8'h27; #100;
A = 8'h2D; B = 8'h28; #100;
A = 8'h2D; B = 8'h29; #100;
A = 8'h2D; B = 8'h2A; #100;
A = 8'h2D; B = 8'h2B; #100;
A = 8'h2D; B = 8'h2C; #100;
A = 8'h2D; B = 8'h2D; #100;
A = 8'h2D; B = 8'h2E; #100;
A = 8'h2D; B = 8'h2F; #100;
A = 8'h2D; B = 8'h30; #100;
A = 8'h2D; B = 8'h31; #100;
A = 8'h2D; B = 8'h32; #100;
A = 8'h2D; B = 8'h33; #100;
A = 8'h2D; B = 8'h34; #100;
A = 8'h2D; B = 8'h35; #100;
A = 8'h2D; B = 8'h36; #100;
A = 8'h2D; B = 8'h37; #100;
A = 8'h2D; B = 8'h38; #100;
A = 8'h2D; B = 8'h39; #100;
A = 8'h2D; B = 8'h3A; #100;
A = 8'h2D; B = 8'h3B; #100;
A = 8'h2D; B = 8'h3C; #100;
A = 8'h2D; B = 8'h3D; #100;
A = 8'h2D; B = 8'h3E; #100;
A = 8'h2D; B = 8'h3F; #100;
A = 8'h2D; B = 8'h40; #100;
A = 8'h2D; B = 8'h41; #100;
A = 8'h2D; B = 8'h42; #100;
A = 8'h2D; B = 8'h43; #100;
A = 8'h2D; B = 8'h44; #100;
A = 8'h2D; B = 8'h45; #100;
A = 8'h2D; B = 8'h46; #100;
A = 8'h2D; B = 8'h47; #100;
A = 8'h2D; B = 8'h48; #100;
A = 8'h2D; B = 8'h49; #100;
A = 8'h2D; B = 8'h4A; #100;
A = 8'h2D; B = 8'h4B; #100;
A = 8'h2D; B = 8'h4C; #100;
A = 8'h2D; B = 8'h4D; #100;
A = 8'h2D; B = 8'h4E; #100;
A = 8'h2D; B = 8'h4F; #100;
A = 8'h2D; B = 8'h50; #100;
A = 8'h2D; B = 8'h51; #100;
A = 8'h2D; B = 8'h52; #100;
A = 8'h2D; B = 8'h53; #100;
A = 8'h2D; B = 8'h54; #100;
A = 8'h2D; B = 8'h55; #100;
A = 8'h2D; B = 8'h56; #100;
A = 8'h2D; B = 8'h57; #100;
A = 8'h2D; B = 8'h58; #100;
A = 8'h2D; B = 8'h59; #100;
A = 8'h2D; B = 8'h5A; #100;
A = 8'h2D; B = 8'h5B; #100;
A = 8'h2D; B = 8'h5C; #100;
A = 8'h2D; B = 8'h5D; #100;
A = 8'h2D; B = 8'h5E; #100;
A = 8'h2D; B = 8'h5F; #100;
A = 8'h2D; B = 8'h60; #100;
A = 8'h2D; B = 8'h61; #100;
A = 8'h2D; B = 8'h62; #100;
A = 8'h2D; B = 8'h63; #100;
A = 8'h2D; B = 8'h64; #100;
A = 8'h2D; B = 8'h65; #100;
A = 8'h2D; B = 8'h66; #100;
A = 8'h2D; B = 8'h67; #100;
A = 8'h2D; B = 8'h68; #100;
A = 8'h2D; B = 8'h69; #100;
A = 8'h2D; B = 8'h6A; #100;
A = 8'h2D; B = 8'h6B; #100;
A = 8'h2D; B = 8'h6C; #100;
A = 8'h2D; B = 8'h6D; #100;
A = 8'h2D; B = 8'h6E; #100;
A = 8'h2D; B = 8'h6F; #100;
A = 8'h2D; B = 8'h70; #100;
A = 8'h2D; B = 8'h71; #100;
A = 8'h2D; B = 8'h72; #100;
A = 8'h2D; B = 8'h73; #100;
A = 8'h2D; B = 8'h74; #100;
A = 8'h2D; B = 8'h75; #100;
A = 8'h2D; B = 8'h76; #100;
A = 8'h2D; B = 8'h77; #100;
A = 8'h2D; B = 8'h78; #100;
A = 8'h2D; B = 8'h79; #100;
A = 8'h2D; B = 8'h7A; #100;
A = 8'h2D; B = 8'h7B; #100;
A = 8'h2D; B = 8'h7C; #100;
A = 8'h2D; B = 8'h7D; #100;
A = 8'h2D; B = 8'h7E; #100;
A = 8'h2D; B = 8'h7F; #100;
A = 8'h2D; B = 8'h80; #100;
A = 8'h2D; B = 8'h81; #100;
A = 8'h2D; B = 8'h82; #100;
A = 8'h2D; B = 8'h83; #100;
A = 8'h2D; B = 8'h84; #100;
A = 8'h2D; B = 8'h85; #100;
A = 8'h2D; B = 8'h86; #100;
A = 8'h2D; B = 8'h87; #100;
A = 8'h2D; B = 8'h88; #100;
A = 8'h2D; B = 8'h89; #100;
A = 8'h2D; B = 8'h8A; #100;
A = 8'h2D; B = 8'h8B; #100;
A = 8'h2D; B = 8'h8C; #100;
A = 8'h2D; B = 8'h8D; #100;
A = 8'h2D; B = 8'h8E; #100;
A = 8'h2D; B = 8'h8F; #100;
A = 8'h2D; B = 8'h90; #100;
A = 8'h2D; B = 8'h91; #100;
A = 8'h2D; B = 8'h92; #100;
A = 8'h2D; B = 8'h93; #100;
A = 8'h2D; B = 8'h94; #100;
A = 8'h2D; B = 8'h95; #100;
A = 8'h2D; B = 8'h96; #100;
A = 8'h2D; B = 8'h97; #100;
A = 8'h2D; B = 8'h98; #100;
A = 8'h2D; B = 8'h99; #100;
A = 8'h2D; B = 8'h9A; #100;
A = 8'h2D; B = 8'h9B; #100;
A = 8'h2D; B = 8'h9C; #100;
A = 8'h2D; B = 8'h9D; #100;
A = 8'h2D; B = 8'h9E; #100;
A = 8'h2D; B = 8'h9F; #100;
A = 8'h2D; B = 8'hA0; #100;
A = 8'h2D; B = 8'hA1; #100;
A = 8'h2D; B = 8'hA2; #100;
A = 8'h2D; B = 8'hA3; #100;
A = 8'h2D; B = 8'hA4; #100;
A = 8'h2D; B = 8'hA5; #100;
A = 8'h2D; B = 8'hA6; #100;
A = 8'h2D; B = 8'hA7; #100;
A = 8'h2D; B = 8'hA8; #100;
A = 8'h2D; B = 8'hA9; #100;
A = 8'h2D; B = 8'hAA; #100;
A = 8'h2D; B = 8'hAB; #100;
A = 8'h2D; B = 8'hAC; #100;
A = 8'h2D; B = 8'hAD; #100;
A = 8'h2D; B = 8'hAE; #100;
A = 8'h2D; B = 8'hAF; #100;
A = 8'h2D; B = 8'hB0; #100;
A = 8'h2D; B = 8'hB1; #100;
A = 8'h2D; B = 8'hB2; #100;
A = 8'h2D; B = 8'hB3; #100;
A = 8'h2D; B = 8'hB4; #100;
A = 8'h2D; B = 8'hB5; #100;
A = 8'h2D; B = 8'hB6; #100;
A = 8'h2D; B = 8'hB7; #100;
A = 8'h2D; B = 8'hB8; #100;
A = 8'h2D; B = 8'hB9; #100;
A = 8'h2D; B = 8'hBA; #100;
A = 8'h2D; B = 8'hBB; #100;
A = 8'h2D; B = 8'hBC; #100;
A = 8'h2D; B = 8'hBD; #100;
A = 8'h2D; B = 8'hBE; #100;
A = 8'h2D; B = 8'hBF; #100;
A = 8'h2D; B = 8'hC0; #100;
A = 8'h2D; B = 8'hC1; #100;
A = 8'h2D; B = 8'hC2; #100;
A = 8'h2D; B = 8'hC3; #100;
A = 8'h2D; B = 8'hC4; #100;
A = 8'h2D; B = 8'hC5; #100;
A = 8'h2D; B = 8'hC6; #100;
A = 8'h2D; B = 8'hC7; #100;
A = 8'h2D; B = 8'hC8; #100;
A = 8'h2D; B = 8'hC9; #100;
A = 8'h2D; B = 8'hCA; #100;
A = 8'h2D; B = 8'hCB; #100;
A = 8'h2D; B = 8'hCC; #100;
A = 8'h2D; B = 8'hCD; #100;
A = 8'h2D; B = 8'hCE; #100;
A = 8'h2D; B = 8'hCF; #100;
A = 8'h2D; B = 8'hD0; #100;
A = 8'h2D; B = 8'hD1; #100;
A = 8'h2D; B = 8'hD2; #100;
A = 8'h2D; B = 8'hD3; #100;
A = 8'h2D; B = 8'hD4; #100;
A = 8'h2D; B = 8'hD5; #100;
A = 8'h2D; B = 8'hD6; #100;
A = 8'h2D; B = 8'hD7; #100;
A = 8'h2D; B = 8'hD8; #100;
A = 8'h2D; B = 8'hD9; #100;
A = 8'h2D; B = 8'hDA; #100;
A = 8'h2D; B = 8'hDB; #100;
A = 8'h2D; B = 8'hDC; #100;
A = 8'h2D; B = 8'hDD; #100;
A = 8'h2D; B = 8'hDE; #100;
A = 8'h2D; B = 8'hDF; #100;
A = 8'h2D; B = 8'hE0; #100;
A = 8'h2D; B = 8'hE1; #100;
A = 8'h2D; B = 8'hE2; #100;
A = 8'h2D; B = 8'hE3; #100;
A = 8'h2D; B = 8'hE4; #100;
A = 8'h2D; B = 8'hE5; #100;
A = 8'h2D; B = 8'hE6; #100;
A = 8'h2D; B = 8'hE7; #100;
A = 8'h2D; B = 8'hE8; #100;
A = 8'h2D; B = 8'hE9; #100;
A = 8'h2D; B = 8'hEA; #100;
A = 8'h2D; B = 8'hEB; #100;
A = 8'h2D; B = 8'hEC; #100;
A = 8'h2D; B = 8'hED; #100;
A = 8'h2D; B = 8'hEE; #100;
A = 8'h2D; B = 8'hEF; #100;
A = 8'h2D; B = 8'hF0; #100;
A = 8'h2D; B = 8'hF1; #100;
A = 8'h2D; B = 8'hF2; #100;
A = 8'h2D; B = 8'hF3; #100;
A = 8'h2D; B = 8'hF4; #100;
A = 8'h2D; B = 8'hF5; #100;
A = 8'h2D; B = 8'hF6; #100;
A = 8'h2D; B = 8'hF7; #100;
A = 8'h2D; B = 8'hF8; #100;
A = 8'h2D; B = 8'hF9; #100;
A = 8'h2D; B = 8'hFA; #100;
A = 8'h2D; B = 8'hFB; #100;
A = 8'h2D; B = 8'hFC; #100;
A = 8'h2D; B = 8'hFD; #100;
A = 8'h2D; B = 8'hFE; #100;
A = 8'h2D; B = 8'hFF; #100;
A = 8'h2E; B = 8'h0; #100;
A = 8'h2E; B = 8'h1; #100;
A = 8'h2E; B = 8'h2; #100;
A = 8'h2E; B = 8'h3; #100;
A = 8'h2E; B = 8'h4; #100;
A = 8'h2E; B = 8'h5; #100;
A = 8'h2E; B = 8'h6; #100;
A = 8'h2E; B = 8'h7; #100;
A = 8'h2E; B = 8'h8; #100;
A = 8'h2E; B = 8'h9; #100;
A = 8'h2E; B = 8'hA; #100;
A = 8'h2E; B = 8'hB; #100;
A = 8'h2E; B = 8'hC; #100;
A = 8'h2E; B = 8'hD; #100;
A = 8'h2E; B = 8'hE; #100;
A = 8'h2E; B = 8'hF; #100;
A = 8'h2E; B = 8'h10; #100;
A = 8'h2E; B = 8'h11; #100;
A = 8'h2E; B = 8'h12; #100;
A = 8'h2E; B = 8'h13; #100;
A = 8'h2E; B = 8'h14; #100;
A = 8'h2E; B = 8'h15; #100;
A = 8'h2E; B = 8'h16; #100;
A = 8'h2E; B = 8'h17; #100;
A = 8'h2E; B = 8'h18; #100;
A = 8'h2E; B = 8'h19; #100;
A = 8'h2E; B = 8'h1A; #100;
A = 8'h2E; B = 8'h1B; #100;
A = 8'h2E; B = 8'h1C; #100;
A = 8'h2E; B = 8'h1D; #100;
A = 8'h2E; B = 8'h1E; #100;
A = 8'h2E; B = 8'h1F; #100;
A = 8'h2E; B = 8'h20; #100;
A = 8'h2E; B = 8'h21; #100;
A = 8'h2E; B = 8'h22; #100;
A = 8'h2E; B = 8'h23; #100;
A = 8'h2E; B = 8'h24; #100;
A = 8'h2E; B = 8'h25; #100;
A = 8'h2E; B = 8'h26; #100;
A = 8'h2E; B = 8'h27; #100;
A = 8'h2E; B = 8'h28; #100;
A = 8'h2E; B = 8'h29; #100;
A = 8'h2E; B = 8'h2A; #100;
A = 8'h2E; B = 8'h2B; #100;
A = 8'h2E; B = 8'h2C; #100;
A = 8'h2E; B = 8'h2D; #100;
A = 8'h2E; B = 8'h2E; #100;
A = 8'h2E; B = 8'h2F; #100;
A = 8'h2E; B = 8'h30; #100;
A = 8'h2E; B = 8'h31; #100;
A = 8'h2E; B = 8'h32; #100;
A = 8'h2E; B = 8'h33; #100;
A = 8'h2E; B = 8'h34; #100;
A = 8'h2E; B = 8'h35; #100;
A = 8'h2E; B = 8'h36; #100;
A = 8'h2E; B = 8'h37; #100;
A = 8'h2E; B = 8'h38; #100;
A = 8'h2E; B = 8'h39; #100;
A = 8'h2E; B = 8'h3A; #100;
A = 8'h2E; B = 8'h3B; #100;
A = 8'h2E; B = 8'h3C; #100;
A = 8'h2E; B = 8'h3D; #100;
A = 8'h2E; B = 8'h3E; #100;
A = 8'h2E; B = 8'h3F; #100;
A = 8'h2E; B = 8'h40; #100;
A = 8'h2E; B = 8'h41; #100;
A = 8'h2E; B = 8'h42; #100;
A = 8'h2E; B = 8'h43; #100;
A = 8'h2E; B = 8'h44; #100;
A = 8'h2E; B = 8'h45; #100;
A = 8'h2E; B = 8'h46; #100;
A = 8'h2E; B = 8'h47; #100;
A = 8'h2E; B = 8'h48; #100;
A = 8'h2E; B = 8'h49; #100;
A = 8'h2E; B = 8'h4A; #100;
A = 8'h2E; B = 8'h4B; #100;
A = 8'h2E; B = 8'h4C; #100;
A = 8'h2E; B = 8'h4D; #100;
A = 8'h2E; B = 8'h4E; #100;
A = 8'h2E; B = 8'h4F; #100;
A = 8'h2E; B = 8'h50; #100;
A = 8'h2E; B = 8'h51; #100;
A = 8'h2E; B = 8'h52; #100;
A = 8'h2E; B = 8'h53; #100;
A = 8'h2E; B = 8'h54; #100;
A = 8'h2E; B = 8'h55; #100;
A = 8'h2E; B = 8'h56; #100;
A = 8'h2E; B = 8'h57; #100;
A = 8'h2E; B = 8'h58; #100;
A = 8'h2E; B = 8'h59; #100;
A = 8'h2E; B = 8'h5A; #100;
A = 8'h2E; B = 8'h5B; #100;
A = 8'h2E; B = 8'h5C; #100;
A = 8'h2E; B = 8'h5D; #100;
A = 8'h2E; B = 8'h5E; #100;
A = 8'h2E; B = 8'h5F; #100;
A = 8'h2E; B = 8'h60; #100;
A = 8'h2E; B = 8'h61; #100;
A = 8'h2E; B = 8'h62; #100;
A = 8'h2E; B = 8'h63; #100;
A = 8'h2E; B = 8'h64; #100;
A = 8'h2E; B = 8'h65; #100;
A = 8'h2E; B = 8'h66; #100;
A = 8'h2E; B = 8'h67; #100;
A = 8'h2E; B = 8'h68; #100;
A = 8'h2E; B = 8'h69; #100;
A = 8'h2E; B = 8'h6A; #100;
A = 8'h2E; B = 8'h6B; #100;
A = 8'h2E; B = 8'h6C; #100;
A = 8'h2E; B = 8'h6D; #100;
A = 8'h2E; B = 8'h6E; #100;
A = 8'h2E; B = 8'h6F; #100;
A = 8'h2E; B = 8'h70; #100;
A = 8'h2E; B = 8'h71; #100;
A = 8'h2E; B = 8'h72; #100;
A = 8'h2E; B = 8'h73; #100;
A = 8'h2E; B = 8'h74; #100;
A = 8'h2E; B = 8'h75; #100;
A = 8'h2E; B = 8'h76; #100;
A = 8'h2E; B = 8'h77; #100;
A = 8'h2E; B = 8'h78; #100;
A = 8'h2E; B = 8'h79; #100;
A = 8'h2E; B = 8'h7A; #100;
A = 8'h2E; B = 8'h7B; #100;
A = 8'h2E; B = 8'h7C; #100;
A = 8'h2E; B = 8'h7D; #100;
A = 8'h2E; B = 8'h7E; #100;
A = 8'h2E; B = 8'h7F; #100;
A = 8'h2E; B = 8'h80; #100;
A = 8'h2E; B = 8'h81; #100;
A = 8'h2E; B = 8'h82; #100;
A = 8'h2E; B = 8'h83; #100;
A = 8'h2E; B = 8'h84; #100;
A = 8'h2E; B = 8'h85; #100;
A = 8'h2E; B = 8'h86; #100;
A = 8'h2E; B = 8'h87; #100;
A = 8'h2E; B = 8'h88; #100;
A = 8'h2E; B = 8'h89; #100;
A = 8'h2E; B = 8'h8A; #100;
A = 8'h2E; B = 8'h8B; #100;
A = 8'h2E; B = 8'h8C; #100;
A = 8'h2E; B = 8'h8D; #100;
A = 8'h2E; B = 8'h8E; #100;
A = 8'h2E; B = 8'h8F; #100;
A = 8'h2E; B = 8'h90; #100;
A = 8'h2E; B = 8'h91; #100;
A = 8'h2E; B = 8'h92; #100;
A = 8'h2E; B = 8'h93; #100;
A = 8'h2E; B = 8'h94; #100;
A = 8'h2E; B = 8'h95; #100;
A = 8'h2E; B = 8'h96; #100;
A = 8'h2E; B = 8'h97; #100;
A = 8'h2E; B = 8'h98; #100;
A = 8'h2E; B = 8'h99; #100;
A = 8'h2E; B = 8'h9A; #100;
A = 8'h2E; B = 8'h9B; #100;
A = 8'h2E; B = 8'h9C; #100;
A = 8'h2E; B = 8'h9D; #100;
A = 8'h2E; B = 8'h9E; #100;
A = 8'h2E; B = 8'h9F; #100;
A = 8'h2E; B = 8'hA0; #100;
A = 8'h2E; B = 8'hA1; #100;
A = 8'h2E; B = 8'hA2; #100;
A = 8'h2E; B = 8'hA3; #100;
A = 8'h2E; B = 8'hA4; #100;
A = 8'h2E; B = 8'hA5; #100;
A = 8'h2E; B = 8'hA6; #100;
A = 8'h2E; B = 8'hA7; #100;
A = 8'h2E; B = 8'hA8; #100;
A = 8'h2E; B = 8'hA9; #100;
A = 8'h2E; B = 8'hAA; #100;
A = 8'h2E; B = 8'hAB; #100;
A = 8'h2E; B = 8'hAC; #100;
A = 8'h2E; B = 8'hAD; #100;
A = 8'h2E; B = 8'hAE; #100;
A = 8'h2E; B = 8'hAF; #100;
A = 8'h2E; B = 8'hB0; #100;
A = 8'h2E; B = 8'hB1; #100;
A = 8'h2E; B = 8'hB2; #100;
A = 8'h2E; B = 8'hB3; #100;
A = 8'h2E; B = 8'hB4; #100;
A = 8'h2E; B = 8'hB5; #100;
A = 8'h2E; B = 8'hB6; #100;
A = 8'h2E; B = 8'hB7; #100;
A = 8'h2E; B = 8'hB8; #100;
A = 8'h2E; B = 8'hB9; #100;
A = 8'h2E; B = 8'hBA; #100;
A = 8'h2E; B = 8'hBB; #100;
A = 8'h2E; B = 8'hBC; #100;
A = 8'h2E; B = 8'hBD; #100;
A = 8'h2E; B = 8'hBE; #100;
A = 8'h2E; B = 8'hBF; #100;
A = 8'h2E; B = 8'hC0; #100;
A = 8'h2E; B = 8'hC1; #100;
A = 8'h2E; B = 8'hC2; #100;
A = 8'h2E; B = 8'hC3; #100;
A = 8'h2E; B = 8'hC4; #100;
A = 8'h2E; B = 8'hC5; #100;
A = 8'h2E; B = 8'hC6; #100;
A = 8'h2E; B = 8'hC7; #100;
A = 8'h2E; B = 8'hC8; #100;
A = 8'h2E; B = 8'hC9; #100;
A = 8'h2E; B = 8'hCA; #100;
A = 8'h2E; B = 8'hCB; #100;
A = 8'h2E; B = 8'hCC; #100;
A = 8'h2E; B = 8'hCD; #100;
A = 8'h2E; B = 8'hCE; #100;
A = 8'h2E; B = 8'hCF; #100;
A = 8'h2E; B = 8'hD0; #100;
A = 8'h2E; B = 8'hD1; #100;
A = 8'h2E; B = 8'hD2; #100;
A = 8'h2E; B = 8'hD3; #100;
A = 8'h2E; B = 8'hD4; #100;
A = 8'h2E; B = 8'hD5; #100;
A = 8'h2E; B = 8'hD6; #100;
A = 8'h2E; B = 8'hD7; #100;
A = 8'h2E; B = 8'hD8; #100;
A = 8'h2E; B = 8'hD9; #100;
A = 8'h2E; B = 8'hDA; #100;
A = 8'h2E; B = 8'hDB; #100;
A = 8'h2E; B = 8'hDC; #100;
A = 8'h2E; B = 8'hDD; #100;
A = 8'h2E; B = 8'hDE; #100;
A = 8'h2E; B = 8'hDF; #100;
A = 8'h2E; B = 8'hE0; #100;
A = 8'h2E; B = 8'hE1; #100;
A = 8'h2E; B = 8'hE2; #100;
A = 8'h2E; B = 8'hE3; #100;
A = 8'h2E; B = 8'hE4; #100;
A = 8'h2E; B = 8'hE5; #100;
A = 8'h2E; B = 8'hE6; #100;
A = 8'h2E; B = 8'hE7; #100;
A = 8'h2E; B = 8'hE8; #100;
A = 8'h2E; B = 8'hE9; #100;
A = 8'h2E; B = 8'hEA; #100;
A = 8'h2E; B = 8'hEB; #100;
A = 8'h2E; B = 8'hEC; #100;
A = 8'h2E; B = 8'hED; #100;
A = 8'h2E; B = 8'hEE; #100;
A = 8'h2E; B = 8'hEF; #100;
A = 8'h2E; B = 8'hF0; #100;
A = 8'h2E; B = 8'hF1; #100;
A = 8'h2E; B = 8'hF2; #100;
A = 8'h2E; B = 8'hF3; #100;
A = 8'h2E; B = 8'hF4; #100;
A = 8'h2E; B = 8'hF5; #100;
A = 8'h2E; B = 8'hF6; #100;
A = 8'h2E; B = 8'hF7; #100;
A = 8'h2E; B = 8'hF8; #100;
A = 8'h2E; B = 8'hF9; #100;
A = 8'h2E; B = 8'hFA; #100;
A = 8'h2E; B = 8'hFB; #100;
A = 8'h2E; B = 8'hFC; #100;
A = 8'h2E; B = 8'hFD; #100;
A = 8'h2E; B = 8'hFE; #100;
A = 8'h2E; B = 8'hFF; #100;
A = 8'h2F; B = 8'h0; #100;
A = 8'h2F; B = 8'h1; #100;
A = 8'h2F; B = 8'h2; #100;
A = 8'h2F; B = 8'h3; #100;
A = 8'h2F; B = 8'h4; #100;
A = 8'h2F; B = 8'h5; #100;
A = 8'h2F; B = 8'h6; #100;
A = 8'h2F; B = 8'h7; #100;
A = 8'h2F; B = 8'h8; #100;
A = 8'h2F; B = 8'h9; #100;
A = 8'h2F; B = 8'hA; #100;
A = 8'h2F; B = 8'hB; #100;
A = 8'h2F; B = 8'hC; #100;
A = 8'h2F; B = 8'hD; #100;
A = 8'h2F; B = 8'hE; #100;
A = 8'h2F; B = 8'hF; #100;
A = 8'h2F; B = 8'h10; #100;
A = 8'h2F; B = 8'h11; #100;
A = 8'h2F; B = 8'h12; #100;
A = 8'h2F; B = 8'h13; #100;
A = 8'h2F; B = 8'h14; #100;
A = 8'h2F; B = 8'h15; #100;
A = 8'h2F; B = 8'h16; #100;
A = 8'h2F; B = 8'h17; #100;
A = 8'h2F; B = 8'h18; #100;
A = 8'h2F; B = 8'h19; #100;
A = 8'h2F; B = 8'h1A; #100;
A = 8'h2F; B = 8'h1B; #100;
A = 8'h2F; B = 8'h1C; #100;
A = 8'h2F; B = 8'h1D; #100;
A = 8'h2F; B = 8'h1E; #100;
A = 8'h2F; B = 8'h1F; #100;
A = 8'h2F; B = 8'h20; #100;
A = 8'h2F; B = 8'h21; #100;
A = 8'h2F; B = 8'h22; #100;
A = 8'h2F; B = 8'h23; #100;
A = 8'h2F; B = 8'h24; #100;
A = 8'h2F; B = 8'h25; #100;
A = 8'h2F; B = 8'h26; #100;
A = 8'h2F; B = 8'h27; #100;
A = 8'h2F; B = 8'h28; #100;
A = 8'h2F; B = 8'h29; #100;
A = 8'h2F; B = 8'h2A; #100;
A = 8'h2F; B = 8'h2B; #100;
A = 8'h2F; B = 8'h2C; #100;
A = 8'h2F; B = 8'h2D; #100;
A = 8'h2F; B = 8'h2E; #100;
A = 8'h2F; B = 8'h2F; #100;
A = 8'h2F; B = 8'h30; #100;
A = 8'h2F; B = 8'h31; #100;
A = 8'h2F; B = 8'h32; #100;
A = 8'h2F; B = 8'h33; #100;
A = 8'h2F; B = 8'h34; #100;
A = 8'h2F; B = 8'h35; #100;
A = 8'h2F; B = 8'h36; #100;
A = 8'h2F; B = 8'h37; #100;
A = 8'h2F; B = 8'h38; #100;
A = 8'h2F; B = 8'h39; #100;
A = 8'h2F; B = 8'h3A; #100;
A = 8'h2F; B = 8'h3B; #100;
A = 8'h2F; B = 8'h3C; #100;
A = 8'h2F; B = 8'h3D; #100;
A = 8'h2F; B = 8'h3E; #100;
A = 8'h2F; B = 8'h3F; #100;
A = 8'h2F; B = 8'h40; #100;
A = 8'h2F; B = 8'h41; #100;
A = 8'h2F; B = 8'h42; #100;
A = 8'h2F; B = 8'h43; #100;
A = 8'h2F; B = 8'h44; #100;
A = 8'h2F; B = 8'h45; #100;
A = 8'h2F; B = 8'h46; #100;
A = 8'h2F; B = 8'h47; #100;
A = 8'h2F; B = 8'h48; #100;
A = 8'h2F; B = 8'h49; #100;
A = 8'h2F; B = 8'h4A; #100;
A = 8'h2F; B = 8'h4B; #100;
A = 8'h2F; B = 8'h4C; #100;
A = 8'h2F; B = 8'h4D; #100;
A = 8'h2F; B = 8'h4E; #100;
A = 8'h2F; B = 8'h4F; #100;
A = 8'h2F; B = 8'h50; #100;
A = 8'h2F; B = 8'h51; #100;
A = 8'h2F; B = 8'h52; #100;
A = 8'h2F; B = 8'h53; #100;
A = 8'h2F; B = 8'h54; #100;
A = 8'h2F; B = 8'h55; #100;
A = 8'h2F; B = 8'h56; #100;
A = 8'h2F; B = 8'h57; #100;
A = 8'h2F; B = 8'h58; #100;
A = 8'h2F; B = 8'h59; #100;
A = 8'h2F; B = 8'h5A; #100;
A = 8'h2F; B = 8'h5B; #100;
A = 8'h2F; B = 8'h5C; #100;
A = 8'h2F; B = 8'h5D; #100;
A = 8'h2F; B = 8'h5E; #100;
A = 8'h2F; B = 8'h5F; #100;
A = 8'h2F; B = 8'h60; #100;
A = 8'h2F; B = 8'h61; #100;
A = 8'h2F; B = 8'h62; #100;
A = 8'h2F; B = 8'h63; #100;
A = 8'h2F; B = 8'h64; #100;
A = 8'h2F; B = 8'h65; #100;
A = 8'h2F; B = 8'h66; #100;
A = 8'h2F; B = 8'h67; #100;
A = 8'h2F; B = 8'h68; #100;
A = 8'h2F; B = 8'h69; #100;
A = 8'h2F; B = 8'h6A; #100;
A = 8'h2F; B = 8'h6B; #100;
A = 8'h2F; B = 8'h6C; #100;
A = 8'h2F; B = 8'h6D; #100;
A = 8'h2F; B = 8'h6E; #100;
A = 8'h2F; B = 8'h6F; #100;
A = 8'h2F; B = 8'h70; #100;
A = 8'h2F; B = 8'h71; #100;
A = 8'h2F; B = 8'h72; #100;
A = 8'h2F; B = 8'h73; #100;
A = 8'h2F; B = 8'h74; #100;
A = 8'h2F; B = 8'h75; #100;
A = 8'h2F; B = 8'h76; #100;
A = 8'h2F; B = 8'h77; #100;
A = 8'h2F; B = 8'h78; #100;
A = 8'h2F; B = 8'h79; #100;
A = 8'h2F; B = 8'h7A; #100;
A = 8'h2F; B = 8'h7B; #100;
A = 8'h2F; B = 8'h7C; #100;
A = 8'h2F; B = 8'h7D; #100;
A = 8'h2F; B = 8'h7E; #100;
A = 8'h2F; B = 8'h7F; #100;
A = 8'h2F; B = 8'h80; #100;
A = 8'h2F; B = 8'h81; #100;
A = 8'h2F; B = 8'h82; #100;
A = 8'h2F; B = 8'h83; #100;
A = 8'h2F; B = 8'h84; #100;
A = 8'h2F; B = 8'h85; #100;
A = 8'h2F; B = 8'h86; #100;
A = 8'h2F; B = 8'h87; #100;
A = 8'h2F; B = 8'h88; #100;
A = 8'h2F; B = 8'h89; #100;
A = 8'h2F; B = 8'h8A; #100;
A = 8'h2F; B = 8'h8B; #100;
A = 8'h2F; B = 8'h8C; #100;
A = 8'h2F; B = 8'h8D; #100;
A = 8'h2F; B = 8'h8E; #100;
A = 8'h2F; B = 8'h8F; #100;
A = 8'h2F; B = 8'h90; #100;
A = 8'h2F; B = 8'h91; #100;
A = 8'h2F; B = 8'h92; #100;
A = 8'h2F; B = 8'h93; #100;
A = 8'h2F; B = 8'h94; #100;
A = 8'h2F; B = 8'h95; #100;
A = 8'h2F; B = 8'h96; #100;
A = 8'h2F; B = 8'h97; #100;
A = 8'h2F; B = 8'h98; #100;
A = 8'h2F; B = 8'h99; #100;
A = 8'h2F; B = 8'h9A; #100;
A = 8'h2F; B = 8'h9B; #100;
A = 8'h2F; B = 8'h9C; #100;
A = 8'h2F; B = 8'h9D; #100;
A = 8'h2F; B = 8'h9E; #100;
A = 8'h2F; B = 8'h9F; #100;
A = 8'h2F; B = 8'hA0; #100;
A = 8'h2F; B = 8'hA1; #100;
A = 8'h2F; B = 8'hA2; #100;
A = 8'h2F; B = 8'hA3; #100;
A = 8'h2F; B = 8'hA4; #100;
A = 8'h2F; B = 8'hA5; #100;
A = 8'h2F; B = 8'hA6; #100;
A = 8'h2F; B = 8'hA7; #100;
A = 8'h2F; B = 8'hA8; #100;
A = 8'h2F; B = 8'hA9; #100;
A = 8'h2F; B = 8'hAA; #100;
A = 8'h2F; B = 8'hAB; #100;
A = 8'h2F; B = 8'hAC; #100;
A = 8'h2F; B = 8'hAD; #100;
A = 8'h2F; B = 8'hAE; #100;
A = 8'h2F; B = 8'hAF; #100;
A = 8'h2F; B = 8'hB0; #100;
A = 8'h2F; B = 8'hB1; #100;
A = 8'h2F; B = 8'hB2; #100;
A = 8'h2F; B = 8'hB3; #100;
A = 8'h2F; B = 8'hB4; #100;
A = 8'h2F; B = 8'hB5; #100;
A = 8'h2F; B = 8'hB6; #100;
A = 8'h2F; B = 8'hB7; #100;
A = 8'h2F; B = 8'hB8; #100;
A = 8'h2F; B = 8'hB9; #100;
A = 8'h2F; B = 8'hBA; #100;
A = 8'h2F; B = 8'hBB; #100;
A = 8'h2F; B = 8'hBC; #100;
A = 8'h2F; B = 8'hBD; #100;
A = 8'h2F; B = 8'hBE; #100;
A = 8'h2F; B = 8'hBF; #100;
A = 8'h2F; B = 8'hC0; #100;
A = 8'h2F; B = 8'hC1; #100;
A = 8'h2F; B = 8'hC2; #100;
A = 8'h2F; B = 8'hC3; #100;
A = 8'h2F; B = 8'hC4; #100;
A = 8'h2F; B = 8'hC5; #100;
A = 8'h2F; B = 8'hC6; #100;
A = 8'h2F; B = 8'hC7; #100;
A = 8'h2F; B = 8'hC8; #100;
A = 8'h2F; B = 8'hC9; #100;
A = 8'h2F; B = 8'hCA; #100;
A = 8'h2F; B = 8'hCB; #100;
A = 8'h2F; B = 8'hCC; #100;
A = 8'h2F; B = 8'hCD; #100;
A = 8'h2F; B = 8'hCE; #100;
A = 8'h2F; B = 8'hCF; #100;
A = 8'h2F; B = 8'hD0; #100;
A = 8'h2F; B = 8'hD1; #100;
A = 8'h2F; B = 8'hD2; #100;
A = 8'h2F; B = 8'hD3; #100;
A = 8'h2F; B = 8'hD4; #100;
A = 8'h2F; B = 8'hD5; #100;
A = 8'h2F; B = 8'hD6; #100;
A = 8'h2F; B = 8'hD7; #100;
A = 8'h2F; B = 8'hD8; #100;
A = 8'h2F; B = 8'hD9; #100;
A = 8'h2F; B = 8'hDA; #100;
A = 8'h2F; B = 8'hDB; #100;
A = 8'h2F; B = 8'hDC; #100;
A = 8'h2F; B = 8'hDD; #100;
A = 8'h2F; B = 8'hDE; #100;
A = 8'h2F; B = 8'hDF; #100;
A = 8'h2F; B = 8'hE0; #100;
A = 8'h2F; B = 8'hE1; #100;
A = 8'h2F; B = 8'hE2; #100;
A = 8'h2F; B = 8'hE3; #100;
A = 8'h2F; B = 8'hE4; #100;
A = 8'h2F; B = 8'hE5; #100;
A = 8'h2F; B = 8'hE6; #100;
A = 8'h2F; B = 8'hE7; #100;
A = 8'h2F; B = 8'hE8; #100;
A = 8'h2F; B = 8'hE9; #100;
A = 8'h2F; B = 8'hEA; #100;
A = 8'h2F; B = 8'hEB; #100;
A = 8'h2F; B = 8'hEC; #100;
A = 8'h2F; B = 8'hED; #100;
A = 8'h2F; B = 8'hEE; #100;
A = 8'h2F; B = 8'hEF; #100;
A = 8'h2F; B = 8'hF0; #100;
A = 8'h2F; B = 8'hF1; #100;
A = 8'h2F; B = 8'hF2; #100;
A = 8'h2F; B = 8'hF3; #100;
A = 8'h2F; B = 8'hF4; #100;
A = 8'h2F; B = 8'hF5; #100;
A = 8'h2F; B = 8'hF6; #100;
A = 8'h2F; B = 8'hF7; #100;
A = 8'h2F; B = 8'hF8; #100;
A = 8'h2F; B = 8'hF9; #100;
A = 8'h2F; B = 8'hFA; #100;
A = 8'h2F; B = 8'hFB; #100;
A = 8'h2F; B = 8'hFC; #100;
A = 8'h2F; B = 8'hFD; #100;
A = 8'h2F; B = 8'hFE; #100;
A = 8'h2F; B = 8'hFF; #100;
A = 8'h30; B = 8'h0; #100;
A = 8'h30; B = 8'h1; #100;
A = 8'h30; B = 8'h2; #100;
A = 8'h30; B = 8'h3; #100;
A = 8'h30; B = 8'h4; #100;
A = 8'h30; B = 8'h5; #100;
A = 8'h30; B = 8'h6; #100;
A = 8'h30; B = 8'h7; #100;
A = 8'h30; B = 8'h8; #100;
A = 8'h30; B = 8'h9; #100;
A = 8'h30; B = 8'hA; #100;
A = 8'h30; B = 8'hB; #100;
A = 8'h30; B = 8'hC; #100;
A = 8'h30; B = 8'hD; #100;
A = 8'h30; B = 8'hE; #100;
A = 8'h30; B = 8'hF; #100;
A = 8'h30; B = 8'h10; #100;
A = 8'h30; B = 8'h11; #100;
A = 8'h30; B = 8'h12; #100;
A = 8'h30; B = 8'h13; #100;
A = 8'h30; B = 8'h14; #100;
A = 8'h30; B = 8'h15; #100;
A = 8'h30; B = 8'h16; #100;
A = 8'h30; B = 8'h17; #100;
A = 8'h30; B = 8'h18; #100;
A = 8'h30; B = 8'h19; #100;
A = 8'h30; B = 8'h1A; #100;
A = 8'h30; B = 8'h1B; #100;
A = 8'h30; B = 8'h1C; #100;
A = 8'h30; B = 8'h1D; #100;
A = 8'h30; B = 8'h1E; #100;
A = 8'h30; B = 8'h1F; #100;
A = 8'h30; B = 8'h20; #100;
A = 8'h30; B = 8'h21; #100;
A = 8'h30; B = 8'h22; #100;
A = 8'h30; B = 8'h23; #100;
A = 8'h30; B = 8'h24; #100;
A = 8'h30; B = 8'h25; #100;
A = 8'h30; B = 8'h26; #100;
A = 8'h30; B = 8'h27; #100;
A = 8'h30; B = 8'h28; #100;
A = 8'h30; B = 8'h29; #100;
A = 8'h30; B = 8'h2A; #100;
A = 8'h30; B = 8'h2B; #100;
A = 8'h30; B = 8'h2C; #100;
A = 8'h30; B = 8'h2D; #100;
A = 8'h30; B = 8'h2E; #100;
A = 8'h30; B = 8'h2F; #100;
A = 8'h30; B = 8'h30; #100;
A = 8'h30; B = 8'h31; #100;
A = 8'h30; B = 8'h32; #100;
A = 8'h30; B = 8'h33; #100;
A = 8'h30; B = 8'h34; #100;
A = 8'h30; B = 8'h35; #100;
A = 8'h30; B = 8'h36; #100;
A = 8'h30; B = 8'h37; #100;
A = 8'h30; B = 8'h38; #100;
A = 8'h30; B = 8'h39; #100;
A = 8'h30; B = 8'h3A; #100;
A = 8'h30; B = 8'h3B; #100;
A = 8'h30; B = 8'h3C; #100;
A = 8'h30; B = 8'h3D; #100;
A = 8'h30; B = 8'h3E; #100;
A = 8'h30; B = 8'h3F; #100;
A = 8'h30; B = 8'h40; #100;
A = 8'h30; B = 8'h41; #100;
A = 8'h30; B = 8'h42; #100;
A = 8'h30; B = 8'h43; #100;
A = 8'h30; B = 8'h44; #100;
A = 8'h30; B = 8'h45; #100;
A = 8'h30; B = 8'h46; #100;
A = 8'h30; B = 8'h47; #100;
A = 8'h30; B = 8'h48; #100;
A = 8'h30; B = 8'h49; #100;
A = 8'h30; B = 8'h4A; #100;
A = 8'h30; B = 8'h4B; #100;
A = 8'h30; B = 8'h4C; #100;
A = 8'h30; B = 8'h4D; #100;
A = 8'h30; B = 8'h4E; #100;
A = 8'h30; B = 8'h4F; #100;
A = 8'h30; B = 8'h50; #100;
A = 8'h30; B = 8'h51; #100;
A = 8'h30; B = 8'h52; #100;
A = 8'h30; B = 8'h53; #100;
A = 8'h30; B = 8'h54; #100;
A = 8'h30; B = 8'h55; #100;
A = 8'h30; B = 8'h56; #100;
A = 8'h30; B = 8'h57; #100;
A = 8'h30; B = 8'h58; #100;
A = 8'h30; B = 8'h59; #100;
A = 8'h30; B = 8'h5A; #100;
A = 8'h30; B = 8'h5B; #100;
A = 8'h30; B = 8'h5C; #100;
A = 8'h30; B = 8'h5D; #100;
A = 8'h30; B = 8'h5E; #100;
A = 8'h30; B = 8'h5F; #100;
A = 8'h30; B = 8'h60; #100;
A = 8'h30; B = 8'h61; #100;
A = 8'h30; B = 8'h62; #100;
A = 8'h30; B = 8'h63; #100;
A = 8'h30; B = 8'h64; #100;
A = 8'h30; B = 8'h65; #100;
A = 8'h30; B = 8'h66; #100;
A = 8'h30; B = 8'h67; #100;
A = 8'h30; B = 8'h68; #100;
A = 8'h30; B = 8'h69; #100;
A = 8'h30; B = 8'h6A; #100;
A = 8'h30; B = 8'h6B; #100;
A = 8'h30; B = 8'h6C; #100;
A = 8'h30; B = 8'h6D; #100;
A = 8'h30; B = 8'h6E; #100;
A = 8'h30; B = 8'h6F; #100;
A = 8'h30; B = 8'h70; #100;
A = 8'h30; B = 8'h71; #100;
A = 8'h30; B = 8'h72; #100;
A = 8'h30; B = 8'h73; #100;
A = 8'h30; B = 8'h74; #100;
A = 8'h30; B = 8'h75; #100;
A = 8'h30; B = 8'h76; #100;
A = 8'h30; B = 8'h77; #100;
A = 8'h30; B = 8'h78; #100;
A = 8'h30; B = 8'h79; #100;
A = 8'h30; B = 8'h7A; #100;
A = 8'h30; B = 8'h7B; #100;
A = 8'h30; B = 8'h7C; #100;
A = 8'h30; B = 8'h7D; #100;
A = 8'h30; B = 8'h7E; #100;
A = 8'h30; B = 8'h7F; #100;
A = 8'h30; B = 8'h80; #100;
A = 8'h30; B = 8'h81; #100;
A = 8'h30; B = 8'h82; #100;
A = 8'h30; B = 8'h83; #100;
A = 8'h30; B = 8'h84; #100;
A = 8'h30; B = 8'h85; #100;
A = 8'h30; B = 8'h86; #100;
A = 8'h30; B = 8'h87; #100;
A = 8'h30; B = 8'h88; #100;
A = 8'h30; B = 8'h89; #100;
A = 8'h30; B = 8'h8A; #100;
A = 8'h30; B = 8'h8B; #100;
A = 8'h30; B = 8'h8C; #100;
A = 8'h30; B = 8'h8D; #100;
A = 8'h30; B = 8'h8E; #100;
A = 8'h30; B = 8'h8F; #100;
A = 8'h30; B = 8'h90; #100;
A = 8'h30; B = 8'h91; #100;
A = 8'h30; B = 8'h92; #100;
A = 8'h30; B = 8'h93; #100;
A = 8'h30; B = 8'h94; #100;
A = 8'h30; B = 8'h95; #100;
A = 8'h30; B = 8'h96; #100;
A = 8'h30; B = 8'h97; #100;
A = 8'h30; B = 8'h98; #100;
A = 8'h30; B = 8'h99; #100;
A = 8'h30; B = 8'h9A; #100;
A = 8'h30; B = 8'h9B; #100;
A = 8'h30; B = 8'h9C; #100;
A = 8'h30; B = 8'h9D; #100;
A = 8'h30; B = 8'h9E; #100;
A = 8'h30; B = 8'h9F; #100;
A = 8'h30; B = 8'hA0; #100;
A = 8'h30; B = 8'hA1; #100;
A = 8'h30; B = 8'hA2; #100;
A = 8'h30; B = 8'hA3; #100;
A = 8'h30; B = 8'hA4; #100;
A = 8'h30; B = 8'hA5; #100;
A = 8'h30; B = 8'hA6; #100;
A = 8'h30; B = 8'hA7; #100;
A = 8'h30; B = 8'hA8; #100;
A = 8'h30; B = 8'hA9; #100;
A = 8'h30; B = 8'hAA; #100;
A = 8'h30; B = 8'hAB; #100;
A = 8'h30; B = 8'hAC; #100;
A = 8'h30; B = 8'hAD; #100;
A = 8'h30; B = 8'hAE; #100;
A = 8'h30; B = 8'hAF; #100;
A = 8'h30; B = 8'hB0; #100;
A = 8'h30; B = 8'hB1; #100;
A = 8'h30; B = 8'hB2; #100;
A = 8'h30; B = 8'hB3; #100;
A = 8'h30; B = 8'hB4; #100;
A = 8'h30; B = 8'hB5; #100;
A = 8'h30; B = 8'hB6; #100;
A = 8'h30; B = 8'hB7; #100;
A = 8'h30; B = 8'hB8; #100;
A = 8'h30; B = 8'hB9; #100;
A = 8'h30; B = 8'hBA; #100;
A = 8'h30; B = 8'hBB; #100;
A = 8'h30; B = 8'hBC; #100;
A = 8'h30; B = 8'hBD; #100;
A = 8'h30; B = 8'hBE; #100;
A = 8'h30; B = 8'hBF; #100;
A = 8'h30; B = 8'hC0; #100;
A = 8'h30; B = 8'hC1; #100;
A = 8'h30; B = 8'hC2; #100;
A = 8'h30; B = 8'hC3; #100;
A = 8'h30; B = 8'hC4; #100;
A = 8'h30; B = 8'hC5; #100;
A = 8'h30; B = 8'hC6; #100;
A = 8'h30; B = 8'hC7; #100;
A = 8'h30; B = 8'hC8; #100;
A = 8'h30; B = 8'hC9; #100;
A = 8'h30; B = 8'hCA; #100;
A = 8'h30; B = 8'hCB; #100;
A = 8'h30; B = 8'hCC; #100;
A = 8'h30; B = 8'hCD; #100;
A = 8'h30; B = 8'hCE; #100;
A = 8'h30; B = 8'hCF; #100;
A = 8'h30; B = 8'hD0; #100;
A = 8'h30; B = 8'hD1; #100;
A = 8'h30; B = 8'hD2; #100;
A = 8'h30; B = 8'hD3; #100;
A = 8'h30; B = 8'hD4; #100;
A = 8'h30; B = 8'hD5; #100;
A = 8'h30; B = 8'hD6; #100;
A = 8'h30; B = 8'hD7; #100;
A = 8'h30; B = 8'hD8; #100;
A = 8'h30; B = 8'hD9; #100;
A = 8'h30; B = 8'hDA; #100;
A = 8'h30; B = 8'hDB; #100;
A = 8'h30; B = 8'hDC; #100;
A = 8'h30; B = 8'hDD; #100;
A = 8'h30; B = 8'hDE; #100;
A = 8'h30; B = 8'hDF; #100;
A = 8'h30; B = 8'hE0; #100;
A = 8'h30; B = 8'hE1; #100;
A = 8'h30; B = 8'hE2; #100;
A = 8'h30; B = 8'hE3; #100;
A = 8'h30; B = 8'hE4; #100;
A = 8'h30; B = 8'hE5; #100;
A = 8'h30; B = 8'hE6; #100;
A = 8'h30; B = 8'hE7; #100;
A = 8'h30; B = 8'hE8; #100;
A = 8'h30; B = 8'hE9; #100;
A = 8'h30; B = 8'hEA; #100;
A = 8'h30; B = 8'hEB; #100;
A = 8'h30; B = 8'hEC; #100;
A = 8'h30; B = 8'hED; #100;
A = 8'h30; B = 8'hEE; #100;
A = 8'h30; B = 8'hEF; #100;
A = 8'h30; B = 8'hF0; #100;
A = 8'h30; B = 8'hF1; #100;
A = 8'h30; B = 8'hF2; #100;
A = 8'h30; B = 8'hF3; #100;
A = 8'h30; B = 8'hF4; #100;
A = 8'h30; B = 8'hF5; #100;
A = 8'h30; B = 8'hF6; #100;
A = 8'h30; B = 8'hF7; #100;
A = 8'h30; B = 8'hF8; #100;
A = 8'h30; B = 8'hF9; #100;
A = 8'h30; B = 8'hFA; #100;
A = 8'h30; B = 8'hFB; #100;
A = 8'h30; B = 8'hFC; #100;
A = 8'h30; B = 8'hFD; #100;
A = 8'h30; B = 8'hFE; #100;
A = 8'h30; B = 8'hFF; #100;
A = 8'h31; B = 8'h0; #100;
A = 8'h31; B = 8'h1; #100;
A = 8'h31; B = 8'h2; #100;
A = 8'h31; B = 8'h3; #100;
A = 8'h31; B = 8'h4; #100;
A = 8'h31; B = 8'h5; #100;
A = 8'h31; B = 8'h6; #100;
A = 8'h31; B = 8'h7; #100;
A = 8'h31; B = 8'h8; #100;
A = 8'h31; B = 8'h9; #100;
A = 8'h31; B = 8'hA; #100;
A = 8'h31; B = 8'hB; #100;
A = 8'h31; B = 8'hC; #100;
A = 8'h31; B = 8'hD; #100;
A = 8'h31; B = 8'hE; #100;
A = 8'h31; B = 8'hF; #100;
A = 8'h31; B = 8'h10; #100;
A = 8'h31; B = 8'h11; #100;
A = 8'h31; B = 8'h12; #100;
A = 8'h31; B = 8'h13; #100;
A = 8'h31; B = 8'h14; #100;
A = 8'h31; B = 8'h15; #100;
A = 8'h31; B = 8'h16; #100;
A = 8'h31; B = 8'h17; #100;
A = 8'h31; B = 8'h18; #100;
A = 8'h31; B = 8'h19; #100;
A = 8'h31; B = 8'h1A; #100;
A = 8'h31; B = 8'h1B; #100;
A = 8'h31; B = 8'h1C; #100;
A = 8'h31; B = 8'h1D; #100;
A = 8'h31; B = 8'h1E; #100;
A = 8'h31; B = 8'h1F; #100;
A = 8'h31; B = 8'h20; #100;
A = 8'h31; B = 8'h21; #100;
A = 8'h31; B = 8'h22; #100;
A = 8'h31; B = 8'h23; #100;
A = 8'h31; B = 8'h24; #100;
A = 8'h31; B = 8'h25; #100;
A = 8'h31; B = 8'h26; #100;
A = 8'h31; B = 8'h27; #100;
A = 8'h31; B = 8'h28; #100;
A = 8'h31; B = 8'h29; #100;
A = 8'h31; B = 8'h2A; #100;
A = 8'h31; B = 8'h2B; #100;
A = 8'h31; B = 8'h2C; #100;
A = 8'h31; B = 8'h2D; #100;
A = 8'h31; B = 8'h2E; #100;
A = 8'h31; B = 8'h2F; #100;
A = 8'h31; B = 8'h30; #100;
A = 8'h31; B = 8'h31; #100;
A = 8'h31; B = 8'h32; #100;
A = 8'h31; B = 8'h33; #100;
A = 8'h31; B = 8'h34; #100;
A = 8'h31; B = 8'h35; #100;
A = 8'h31; B = 8'h36; #100;
A = 8'h31; B = 8'h37; #100;
A = 8'h31; B = 8'h38; #100;
A = 8'h31; B = 8'h39; #100;
A = 8'h31; B = 8'h3A; #100;
A = 8'h31; B = 8'h3B; #100;
A = 8'h31; B = 8'h3C; #100;
A = 8'h31; B = 8'h3D; #100;
A = 8'h31; B = 8'h3E; #100;
A = 8'h31; B = 8'h3F; #100;
A = 8'h31; B = 8'h40; #100;
A = 8'h31; B = 8'h41; #100;
A = 8'h31; B = 8'h42; #100;
A = 8'h31; B = 8'h43; #100;
A = 8'h31; B = 8'h44; #100;
A = 8'h31; B = 8'h45; #100;
A = 8'h31; B = 8'h46; #100;
A = 8'h31; B = 8'h47; #100;
A = 8'h31; B = 8'h48; #100;
A = 8'h31; B = 8'h49; #100;
A = 8'h31; B = 8'h4A; #100;
A = 8'h31; B = 8'h4B; #100;
A = 8'h31; B = 8'h4C; #100;
A = 8'h31; B = 8'h4D; #100;
A = 8'h31; B = 8'h4E; #100;
A = 8'h31; B = 8'h4F; #100;
A = 8'h31; B = 8'h50; #100;
A = 8'h31; B = 8'h51; #100;
A = 8'h31; B = 8'h52; #100;
A = 8'h31; B = 8'h53; #100;
A = 8'h31; B = 8'h54; #100;
A = 8'h31; B = 8'h55; #100;
A = 8'h31; B = 8'h56; #100;
A = 8'h31; B = 8'h57; #100;
A = 8'h31; B = 8'h58; #100;
A = 8'h31; B = 8'h59; #100;
A = 8'h31; B = 8'h5A; #100;
A = 8'h31; B = 8'h5B; #100;
A = 8'h31; B = 8'h5C; #100;
A = 8'h31; B = 8'h5D; #100;
A = 8'h31; B = 8'h5E; #100;
A = 8'h31; B = 8'h5F; #100;
A = 8'h31; B = 8'h60; #100;
A = 8'h31; B = 8'h61; #100;
A = 8'h31; B = 8'h62; #100;
A = 8'h31; B = 8'h63; #100;
A = 8'h31; B = 8'h64; #100;
A = 8'h31; B = 8'h65; #100;
A = 8'h31; B = 8'h66; #100;
A = 8'h31; B = 8'h67; #100;
A = 8'h31; B = 8'h68; #100;
A = 8'h31; B = 8'h69; #100;
A = 8'h31; B = 8'h6A; #100;
A = 8'h31; B = 8'h6B; #100;
A = 8'h31; B = 8'h6C; #100;
A = 8'h31; B = 8'h6D; #100;
A = 8'h31; B = 8'h6E; #100;
A = 8'h31; B = 8'h6F; #100;
A = 8'h31; B = 8'h70; #100;
A = 8'h31; B = 8'h71; #100;
A = 8'h31; B = 8'h72; #100;
A = 8'h31; B = 8'h73; #100;
A = 8'h31; B = 8'h74; #100;
A = 8'h31; B = 8'h75; #100;
A = 8'h31; B = 8'h76; #100;
A = 8'h31; B = 8'h77; #100;
A = 8'h31; B = 8'h78; #100;
A = 8'h31; B = 8'h79; #100;
A = 8'h31; B = 8'h7A; #100;
A = 8'h31; B = 8'h7B; #100;
A = 8'h31; B = 8'h7C; #100;
A = 8'h31; B = 8'h7D; #100;
A = 8'h31; B = 8'h7E; #100;
A = 8'h31; B = 8'h7F; #100;
A = 8'h31; B = 8'h80; #100;
A = 8'h31; B = 8'h81; #100;
A = 8'h31; B = 8'h82; #100;
A = 8'h31; B = 8'h83; #100;
A = 8'h31; B = 8'h84; #100;
A = 8'h31; B = 8'h85; #100;
A = 8'h31; B = 8'h86; #100;
A = 8'h31; B = 8'h87; #100;
A = 8'h31; B = 8'h88; #100;
A = 8'h31; B = 8'h89; #100;
A = 8'h31; B = 8'h8A; #100;
A = 8'h31; B = 8'h8B; #100;
A = 8'h31; B = 8'h8C; #100;
A = 8'h31; B = 8'h8D; #100;
A = 8'h31; B = 8'h8E; #100;
A = 8'h31; B = 8'h8F; #100;
A = 8'h31; B = 8'h90; #100;
A = 8'h31; B = 8'h91; #100;
A = 8'h31; B = 8'h92; #100;
A = 8'h31; B = 8'h93; #100;
A = 8'h31; B = 8'h94; #100;
A = 8'h31; B = 8'h95; #100;
A = 8'h31; B = 8'h96; #100;
A = 8'h31; B = 8'h97; #100;
A = 8'h31; B = 8'h98; #100;
A = 8'h31; B = 8'h99; #100;
A = 8'h31; B = 8'h9A; #100;
A = 8'h31; B = 8'h9B; #100;
A = 8'h31; B = 8'h9C; #100;
A = 8'h31; B = 8'h9D; #100;
A = 8'h31; B = 8'h9E; #100;
A = 8'h31; B = 8'h9F; #100;
A = 8'h31; B = 8'hA0; #100;
A = 8'h31; B = 8'hA1; #100;
A = 8'h31; B = 8'hA2; #100;
A = 8'h31; B = 8'hA3; #100;
A = 8'h31; B = 8'hA4; #100;
A = 8'h31; B = 8'hA5; #100;
A = 8'h31; B = 8'hA6; #100;
A = 8'h31; B = 8'hA7; #100;
A = 8'h31; B = 8'hA8; #100;
A = 8'h31; B = 8'hA9; #100;
A = 8'h31; B = 8'hAA; #100;
A = 8'h31; B = 8'hAB; #100;
A = 8'h31; B = 8'hAC; #100;
A = 8'h31; B = 8'hAD; #100;
A = 8'h31; B = 8'hAE; #100;
A = 8'h31; B = 8'hAF; #100;
A = 8'h31; B = 8'hB0; #100;
A = 8'h31; B = 8'hB1; #100;
A = 8'h31; B = 8'hB2; #100;
A = 8'h31; B = 8'hB3; #100;
A = 8'h31; B = 8'hB4; #100;
A = 8'h31; B = 8'hB5; #100;
A = 8'h31; B = 8'hB6; #100;
A = 8'h31; B = 8'hB7; #100;
A = 8'h31; B = 8'hB8; #100;
A = 8'h31; B = 8'hB9; #100;
A = 8'h31; B = 8'hBA; #100;
A = 8'h31; B = 8'hBB; #100;
A = 8'h31; B = 8'hBC; #100;
A = 8'h31; B = 8'hBD; #100;
A = 8'h31; B = 8'hBE; #100;
A = 8'h31; B = 8'hBF; #100;
A = 8'h31; B = 8'hC0; #100;
A = 8'h31; B = 8'hC1; #100;
A = 8'h31; B = 8'hC2; #100;
A = 8'h31; B = 8'hC3; #100;
A = 8'h31; B = 8'hC4; #100;
A = 8'h31; B = 8'hC5; #100;
A = 8'h31; B = 8'hC6; #100;
A = 8'h31; B = 8'hC7; #100;
A = 8'h31; B = 8'hC8; #100;
A = 8'h31; B = 8'hC9; #100;
A = 8'h31; B = 8'hCA; #100;
A = 8'h31; B = 8'hCB; #100;
A = 8'h31; B = 8'hCC; #100;
A = 8'h31; B = 8'hCD; #100;
A = 8'h31; B = 8'hCE; #100;
A = 8'h31; B = 8'hCF; #100;
A = 8'h31; B = 8'hD0; #100;
A = 8'h31; B = 8'hD1; #100;
A = 8'h31; B = 8'hD2; #100;
A = 8'h31; B = 8'hD3; #100;
A = 8'h31; B = 8'hD4; #100;
A = 8'h31; B = 8'hD5; #100;
A = 8'h31; B = 8'hD6; #100;
A = 8'h31; B = 8'hD7; #100;
A = 8'h31; B = 8'hD8; #100;
A = 8'h31; B = 8'hD9; #100;
A = 8'h31; B = 8'hDA; #100;
A = 8'h31; B = 8'hDB; #100;
A = 8'h31; B = 8'hDC; #100;
A = 8'h31; B = 8'hDD; #100;
A = 8'h31; B = 8'hDE; #100;
A = 8'h31; B = 8'hDF; #100;
A = 8'h31; B = 8'hE0; #100;
A = 8'h31; B = 8'hE1; #100;
A = 8'h31; B = 8'hE2; #100;
A = 8'h31; B = 8'hE3; #100;
A = 8'h31; B = 8'hE4; #100;
A = 8'h31; B = 8'hE5; #100;
A = 8'h31; B = 8'hE6; #100;
A = 8'h31; B = 8'hE7; #100;
A = 8'h31; B = 8'hE8; #100;
A = 8'h31; B = 8'hE9; #100;
A = 8'h31; B = 8'hEA; #100;
A = 8'h31; B = 8'hEB; #100;
A = 8'h31; B = 8'hEC; #100;
A = 8'h31; B = 8'hED; #100;
A = 8'h31; B = 8'hEE; #100;
A = 8'h31; B = 8'hEF; #100;
A = 8'h31; B = 8'hF0; #100;
A = 8'h31; B = 8'hF1; #100;
A = 8'h31; B = 8'hF2; #100;
A = 8'h31; B = 8'hF3; #100;
A = 8'h31; B = 8'hF4; #100;
A = 8'h31; B = 8'hF5; #100;
A = 8'h31; B = 8'hF6; #100;
A = 8'h31; B = 8'hF7; #100;
A = 8'h31; B = 8'hF8; #100;
A = 8'h31; B = 8'hF9; #100;
A = 8'h31; B = 8'hFA; #100;
A = 8'h31; B = 8'hFB; #100;
A = 8'h31; B = 8'hFC; #100;
A = 8'h31; B = 8'hFD; #100;
A = 8'h31; B = 8'hFE; #100;
A = 8'h31; B = 8'hFF; #100;
A = 8'h32; B = 8'h0; #100;
A = 8'h32; B = 8'h1; #100;
A = 8'h32; B = 8'h2; #100;
A = 8'h32; B = 8'h3; #100;
A = 8'h32; B = 8'h4; #100;
A = 8'h32; B = 8'h5; #100;
A = 8'h32; B = 8'h6; #100;
A = 8'h32; B = 8'h7; #100;
A = 8'h32; B = 8'h8; #100;
A = 8'h32; B = 8'h9; #100;
A = 8'h32; B = 8'hA; #100;
A = 8'h32; B = 8'hB; #100;
A = 8'h32; B = 8'hC; #100;
A = 8'h32; B = 8'hD; #100;
A = 8'h32; B = 8'hE; #100;
A = 8'h32; B = 8'hF; #100;
A = 8'h32; B = 8'h10; #100;
A = 8'h32; B = 8'h11; #100;
A = 8'h32; B = 8'h12; #100;
A = 8'h32; B = 8'h13; #100;
A = 8'h32; B = 8'h14; #100;
A = 8'h32; B = 8'h15; #100;
A = 8'h32; B = 8'h16; #100;
A = 8'h32; B = 8'h17; #100;
A = 8'h32; B = 8'h18; #100;
A = 8'h32; B = 8'h19; #100;
A = 8'h32; B = 8'h1A; #100;
A = 8'h32; B = 8'h1B; #100;
A = 8'h32; B = 8'h1C; #100;
A = 8'h32; B = 8'h1D; #100;
A = 8'h32; B = 8'h1E; #100;
A = 8'h32; B = 8'h1F; #100;
A = 8'h32; B = 8'h20; #100;
A = 8'h32; B = 8'h21; #100;
A = 8'h32; B = 8'h22; #100;
A = 8'h32; B = 8'h23; #100;
A = 8'h32; B = 8'h24; #100;
A = 8'h32; B = 8'h25; #100;
A = 8'h32; B = 8'h26; #100;
A = 8'h32; B = 8'h27; #100;
A = 8'h32; B = 8'h28; #100;
A = 8'h32; B = 8'h29; #100;
A = 8'h32; B = 8'h2A; #100;
A = 8'h32; B = 8'h2B; #100;
A = 8'h32; B = 8'h2C; #100;
A = 8'h32; B = 8'h2D; #100;
A = 8'h32; B = 8'h2E; #100;
A = 8'h32; B = 8'h2F; #100;
A = 8'h32; B = 8'h30; #100;
A = 8'h32; B = 8'h31; #100;
A = 8'h32; B = 8'h32; #100;
A = 8'h32; B = 8'h33; #100;
A = 8'h32; B = 8'h34; #100;
A = 8'h32; B = 8'h35; #100;
A = 8'h32; B = 8'h36; #100;
A = 8'h32; B = 8'h37; #100;
A = 8'h32; B = 8'h38; #100;
A = 8'h32; B = 8'h39; #100;
A = 8'h32; B = 8'h3A; #100;
A = 8'h32; B = 8'h3B; #100;
A = 8'h32; B = 8'h3C; #100;
A = 8'h32; B = 8'h3D; #100;
A = 8'h32; B = 8'h3E; #100;
A = 8'h32; B = 8'h3F; #100;
A = 8'h32; B = 8'h40; #100;
A = 8'h32; B = 8'h41; #100;
A = 8'h32; B = 8'h42; #100;
A = 8'h32; B = 8'h43; #100;
A = 8'h32; B = 8'h44; #100;
A = 8'h32; B = 8'h45; #100;
A = 8'h32; B = 8'h46; #100;
A = 8'h32; B = 8'h47; #100;
A = 8'h32; B = 8'h48; #100;
A = 8'h32; B = 8'h49; #100;
A = 8'h32; B = 8'h4A; #100;
A = 8'h32; B = 8'h4B; #100;
A = 8'h32; B = 8'h4C; #100;
A = 8'h32; B = 8'h4D; #100;
A = 8'h32; B = 8'h4E; #100;
A = 8'h32; B = 8'h4F; #100;
A = 8'h32; B = 8'h50; #100;
A = 8'h32; B = 8'h51; #100;
A = 8'h32; B = 8'h52; #100;
A = 8'h32; B = 8'h53; #100;
A = 8'h32; B = 8'h54; #100;
A = 8'h32; B = 8'h55; #100;
A = 8'h32; B = 8'h56; #100;
A = 8'h32; B = 8'h57; #100;
A = 8'h32; B = 8'h58; #100;
A = 8'h32; B = 8'h59; #100;
A = 8'h32; B = 8'h5A; #100;
A = 8'h32; B = 8'h5B; #100;
A = 8'h32; B = 8'h5C; #100;
A = 8'h32; B = 8'h5D; #100;
A = 8'h32; B = 8'h5E; #100;
A = 8'h32; B = 8'h5F; #100;
A = 8'h32; B = 8'h60; #100;
A = 8'h32; B = 8'h61; #100;
A = 8'h32; B = 8'h62; #100;
A = 8'h32; B = 8'h63; #100;
A = 8'h32; B = 8'h64; #100;
A = 8'h32; B = 8'h65; #100;
A = 8'h32; B = 8'h66; #100;
A = 8'h32; B = 8'h67; #100;
A = 8'h32; B = 8'h68; #100;
A = 8'h32; B = 8'h69; #100;
A = 8'h32; B = 8'h6A; #100;
A = 8'h32; B = 8'h6B; #100;
A = 8'h32; B = 8'h6C; #100;
A = 8'h32; B = 8'h6D; #100;
A = 8'h32; B = 8'h6E; #100;
A = 8'h32; B = 8'h6F; #100;
A = 8'h32; B = 8'h70; #100;
A = 8'h32; B = 8'h71; #100;
A = 8'h32; B = 8'h72; #100;
A = 8'h32; B = 8'h73; #100;
A = 8'h32; B = 8'h74; #100;
A = 8'h32; B = 8'h75; #100;
A = 8'h32; B = 8'h76; #100;
A = 8'h32; B = 8'h77; #100;
A = 8'h32; B = 8'h78; #100;
A = 8'h32; B = 8'h79; #100;
A = 8'h32; B = 8'h7A; #100;
A = 8'h32; B = 8'h7B; #100;
A = 8'h32; B = 8'h7C; #100;
A = 8'h32; B = 8'h7D; #100;
A = 8'h32; B = 8'h7E; #100;
A = 8'h32; B = 8'h7F; #100;
A = 8'h32; B = 8'h80; #100;
A = 8'h32; B = 8'h81; #100;
A = 8'h32; B = 8'h82; #100;
A = 8'h32; B = 8'h83; #100;
A = 8'h32; B = 8'h84; #100;
A = 8'h32; B = 8'h85; #100;
A = 8'h32; B = 8'h86; #100;
A = 8'h32; B = 8'h87; #100;
A = 8'h32; B = 8'h88; #100;
A = 8'h32; B = 8'h89; #100;
A = 8'h32; B = 8'h8A; #100;
A = 8'h32; B = 8'h8B; #100;
A = 8'h32; B = 8'h8C; #100;
A = 8'h32; B = 8'h8D; #100;
A = 8'h32; B = 8'h8E; #100;
A = 8'h32; B = 8'h8F; #100;
A = 8'h32; B = 8'h90; #100;
A = 8'h32; B = 8'h91; #100;
A = 8'h32; B = 8'h92; #100;
A = 8'h32; B = 8'h93; #100;
A = 8'h32; B = 8'h94; #100;
A = 8'h32; B = 8'h95; #100;
A = 8'h32; B = 8'h96; #100;
A = 8'h32; B = 8'h97; #100;
A = 8'h32; B = 8'h98; #100;
A = 8'h32; B = 8'h99; #100;
A = 8'h32; B = 8'h9A; #100;
A = 8'h32; B = 8'h9B; #100;
A = 8'h32; B = 8'h9C; #100;
A = 8'h32; B = 8'h9D; #100;
A = 8'h32; B = 8'h9E; #100;
A = 8'h32; B = 8'h9F; #100;
A = 8'h32; B = 8'hA0; #100;
A = 8'h32; B = 8'hA1; #100;
A = 8'h32; B = 8'hA2; #100;
A = 8'h32; B = 8'hA3; #100;
A = 8'h32; B = 8'hA4; #100;
A = 8'h32; B = 8'hA5; #100;
A = 8'h32; B = 8'hA6; #100;
A = 8'h32; B = 8'hA7; #100;
A = 8'h32; B = 8'hA8; #100;
A = 8'h32; B = 8'hA9; #100;
A = 8'h32; B = 8'hAA; #100;
A = 8'h32; B = 8'hAB; #100;
A = 8'h32; B = 8'hAC; #100;
A = 8'h32; B = 8'hAD; #100;
A = 8'h32; B = 8'hAE; #100;
A = 8'h32; B = 8'hAF; #100;
A = 8'h32; B = 8'hB0; #100;
A = 8'h32; B = 8'hB1; #100;
A = 8'h32; B = 8'hB2; #100;
A = 8'h32; B = 8'hB3; #100;
A = 8'h32; B = 8'hB4; #100;
A = 8'h32; B = 8'hB5; #100;
A = 8'h32; B = 8'hB6; #100;
A = 8'h32; B = 8'hB7; #100;
A = 8'h32; B = 8'hB8; #100;
A = 8'h32; B = 8'hB9; #100;
A = 8'h32; B = 8'hBA; #100;
A = 8'h32; B = 8'hBB; #100;
A = 8'h32; B = 8'hBC; #100;
A = 8'h32; B = 8'hBD; #100;
A = 8'h32; B = 8'hBE; #100;
A = 8'h32; B = 8'hBF; #100;
A = 8'h32; B = 8'hC0; #100;
A = 8'h32; B = 8'hC1; #100;
A = 8'h32; B = 8'hC2; #100;
A = 8'h32; B = 8'hC3; #100;
A = 8'h32; B = 8'hC4; #100;
A = 8'h32; B = 8'hC5; #100;
A = 8'h32; B = 8'hC6; #100;
A = 8'h32; B = 8'hC7; #100;
A = 8'h32; B = 8'hC8; #100;
A = 8'h32; B = 8'hC9; #100;
A = 8'h32; B = 8'hCA; #100;
A = 8'h32; B = 8'hCB; #100;
A = 8'h32; B = 8'hCC; #100;
A = 8'h32; B = 8'hCD; #100;
A = 8'h32; B = 8'hCE; #100;
A = 8'h32; B = 8'hCF; #100;
A = 8'h32; B = 8'hD0; #100;
A = 8'h32; B = 8'hD1; #100;
A = 8'h32; B = 8'hD2; #100;
A = 8'h32; B = 8'hD3; #100;
A = 8'h32; B = 8'hD4; #100;
A = 8'h32; B = 8'hD5; #100;
A = 8'h32; B = 8'hD6; #100;
A = 8'h32; B = 8'hD7; #100;
A = 8'h32; B = 8'hD8; #100;
A = 8'h32; B = 8'hD9; #100;
A = 8'h32; B = 8'hDA; #100;
A = 8'h32; B = 8'hDB; #100;
A = 8'h32; B = 8'hDC; #100;
A = 8'h32; B = 8'hDD; #100;
A = 8'h32; B = 8'hDE; #100;
A = 8'h32; B = 8'hDF; #100;
A = 8'h32; B = 8'hE0; #100;
A = 8'h32; B = 8'hE1; #100;
A = 8'h32; B = 8'hE2; #100;
A = 8'h32; B = 8'hE3; #100;
A = 8'h32; B = 8'hE4; #100;
A = 8'h32; B = 8'hE5; #100;
A = 8'h32; B = 8'hE6; #100;
A = 8'h32; B = 8'hE7; #100;
A = 8'h32; B = 8'hE8; #100;
A = 8'h32; B = 8'hE9; #100;
A = 8'h32; B = 8'hEA; #100;
A = 8'h32; B = 8'hEB; #100;
A = 8'h32; B = 8'hEC; #100;
A = 8'h32; B = 8'hED; #100;
A = 8'h32; B = 8'hEE; #100;
A = 8'h32; B = 8'hEF; #100;
A = 8'h32; B = 8'hF0; #100;
A = 8'h32; B = 8'hF1; #100;
A = 8'h32; B = 8'hF2; #100;
A = 8'h32; B = 8'hF3; #100;
A = 8'h32; B = 8'hF4; #100;
A = 8'h32; B = 8'hF5; #100;
A = 8'h32; B = 8'hF6; #100;
A = 8'h32; B = 8'hF7; #100;
A = 8'h32; B = 8'hF8; #100;
A = 8'h32; B = 8'hF9; #100;
A = 8'h32; B = 8'hFA; #100;
A = 8'h32; B = 8'hFB; #100;
A = 8'h32; B = 8'hFC; #100;
A = 8'h32; B = 8'hFD; #100;
A = 8'h32; B = 8'hFE; #100;
A = 8'h32; B = 8'hFF; #100;
A = 8'h33; B = 8'h0; #100;
A = 8'h33; B = 8'h1; #100;
A = 8'h33; B = 8'h2; #100;
A = 8'h33; B = 8'h3; #100;
A = 8'h33; B = 8'h4; #100;
A = 8'h33; B = 8'h5; #100;
A = 8'h33; B = 8'h6; #100;
A = 8'h33; B = 8'h7; #100;
A = 8'h33; B = 8'h8; #100;
A = 8'h33; B = 8'h9; #100;
A = 8'h33; B = 8'hA; #100;
A = 8'h33; B = 8'hB; #100;
A = 8'h33; B = 8'hC; #100;
A = 8'h33; B = 8'hD; #100;
A = 8'h33; B = 8'hE; #100;
A = 8'h33; B = 8'hF; #100;
A = 8'h33; B = 8'h10; #100;
A = 8'h33; B = 8'h11; #100;
A = 8'h33; B = 8'h12; #100;
A = 8'h33; B = 8'h13; #100;
A = 8'h33; B = 8'h14; #100;
A = 8'h33; B = 8'h15; #100;
A = 8'h33; B = 8'h16; #100;
A = 8'h33; B = 8'h17; #100;
A = 8'h33; B = 8'h18; #100;
A = 8'h33; B = 8'h19; #100;
A = 8'h33; B = 8'h1A; #100;
A = 8'h33; B = 8'h1B; #100;
A = 8'h33; B = 8'h1C; #100;
A = 8'h33; B = 8'h1D; #100;
A = 8'h33; B = 8'h1E; #100;
A = 8'h33; B = 8'h1F; #100;
A = 8'h33; B = 8'h20; #100;
A = 8'h33; B = 8'h21; #100;
A = 8'h33; B = 8'h22; #100;
A = 8'h33; B = 8'h23; #100;
A = 8'h33; B = 8'h24; #100;
A = 8'h33; B = 8'h25; #100;
A = 8'h33; B = 8'h26; #100;
A = 8'h33; B = 8'h27; #100;
A = 8'h33; B = 8'h28; #100;
A = 8'h33; B = 8'h29; #100;
A = 8'h33; B = 8'h2A; #100;
A = 8'h33; B = 8'h2B; #100;
A = 8'h33; B = 8'h2C; #100;
A = 8'h33; B = 8'h2D; #100;
A = 8'h33; B = 8'h2E; #100;
A = 8'h33; B = 8'h2F; #100;
A = 8'h33; B = 8'h30; #100;
A = 8'h33; B = 8'h31; #100;
A = 8'h33; B = 8'h32; #100;
A = 8'h33; B = 8'h33; #100;
A = 8'h33; B = 8'h34; #100;
A = 8'h33; B = 8'h35; #100;
A = 8'h33; B = 8'h36; #100;
A = 8'h33; B = 8'h37; #100;
A = 8'h33; B = 8'h38; #100;
A = 8'h33; B = 8'h39; #100;
A = 8'h33; B = 8'h3A; #100;
A = 8'h33; B = 8'h3B; #100;
A = 8'h33; B = 8'h3C; #100;
A = 8'h33; B = 8'h3D; #100;
A = 8'h33; B = 8'h3E; #100;
A = 8'h33; B = 8'h3F; #100;
A = 8'h33; B = 8'h40; #100;
A = 8'h33; B = 8'h41; #100;
A = 8'h33; B = 8'h42; #100;
A = 8'h33; B = 8'h43; #100;
A = 8'h33; B = 8'h44; #100;
A = 8'h33; B = 8'h45; #100;
A = 8'h33; B = 8'h46; #100;
A = 8'h33; B = 8'h47; #100;
A = 8'h33; B = 8'h48; #100;
A = 8'h33; B = 8'h49; #100;
A = 8'h33; B = 8'h4A; #100;
A = 8'h33; B = 8'h4B; #100;
A = 8'h33; B = 8'h4C; #100;
A = 8'h33; B = 8'h4D; #100;
A = 8'h33; B = 8'h4E; #100;
A = 8'h33; B = 8'h4F; #100;
A = 8'h33; B = 8'h50; #100;
A = 8'h33; B = 8'h51; #100;
A = 8'h33; B = 8'h52; #100;
A = 8'h33; B = 8'h53; #100;
A = 8'h33; B = 8'h54; #100;
A = 8'h33; B = 8'h55; #100;
A = 8'h33; B = 8'h56; #100;
A = 8'h33; B = 8'h57; #100;
A = 8'h33; B = 8'h58; #100;
A = 8'h33; B = 8'h59; #100;
A = 8'h33; B = 8'h5A; #100;
A = 8'h33; B = 8'h5B; #100;
A = 8'h33; B = 8'h5C; #100;
A = 8'h33; B = 8'h5D; #100;
A = 8'h33; B = 8'h5E; #100;
A = 8'h33; B = 8'h5F; #100;
A = 8'h33; B = 8'h60; #100;
A = 8'h33; B = 8'h61; #100;
A = 8'h33; B = 8'h62; #100;
A = 8'h33; B = 8'h63; #100;
A = 8'h33; B = 8'h64; #100;
A = 8'h33; B = 8'h65; #100;
A = 8'h33; B = 8'h66; #100;
A = 8'h33; B = 8'h67; #100;
A = 8'h33; B = 8'h68; #100;
A = 8'h33; B = 8'h69; #100;
A = 8'h33; B = 8'h6A; #100;
A = 8'h33; B = 8'h6B; #100;
A = 8'h33; B = 8'h6C; #100;
A = 8'h33; B = 8'h6D; #100;
A = 8'h33; B = 8'h6E; #100;
A = 8'h33; B = 8'h6F; #100;
A = 8'h33; B = 8'h70; #100;
A = 8'h33; B = 8'h71; #100;
A = 8'h33; B = 8'h72; #100;
A = 8'h33; B = 8'h73; #100;
A = 8'h33; B = 8'h74; #100;
A = 8'h33; B = 8'h75; #100;
A = 8'h33; B = 8'h76; #100;
A = 8'h33; B = 8'h77; #100;
A = 8'h33; B = 8'h78; #100;
A = 8'h33; B = 8'h79; #100;
A = 8'h33; B = 8'h7A; #100;
A = 8'h33; B = 8'h7B; #100;
A = 8'h33; B = 8'h7C; #100;
A = 8'h33; B = 8'h7D; #100;
A = 8'h33; B = 8'h7E; #100;
A = 8'h33; B = 8'h7F; #100;
A = 8'h33; B = 8'h80; #100;
A = 8'h33; B = 8'h81; #100;
A = 8'h33; B = 8'h82; #100;
A = 8'h33; B = 8'h83; #100;
A = 8'h33; B = 8'h84; #100;
A = 8'h33; B = 8'h85; #100;
A = 8'h33; B = 8'h86; #100;
A = 8'h33; B = 8'h87; #100;
A = 8'h33; B = 8'h88; #100;
A = 8'h33; B = 8'h89; #100;
A = 8'h33; B = 8'h8A; #100;
A = 8'h33; B = 8'h8B; #100;
A = 8'h33; B = 8'h8C; #100;
A = 8'h33; B = 8'h8D; #100;
A = 8'h33; B = 8'h8E; #100;
A = 8'h33; B = 8'h8F; #100;
A = 8'h33; B = 8'h90; #100;
A = 8'h33; B = 8'h91; #100;
A = 8'h33; B = 8'h92; #100;
A = 8'h33; B = 8'h93; #100;
A = 8'h33; B = 8'h94; #100;
A = 8'h33; B = 8'h95; #100;
A = 8'h33; B = 8'h96; #100;
A = 8'h33; B = 8'h97; #100;
A = 8'h33; B = 8'h98; #100;
A = 8'h33; B = 8'h99; #100;
A = 8'h33; B = 8'h9A; #100;
A = 8'h33; B = 8'h9B; #100;
A = 8'h33; B = 8'h9C; #100;
A = 8'h33; B = 8'h9D; #100;
A = 8'h33; B = 8'h9E; #100;
A = 8'h33; B = 8'h9F; #100;
A = 8'h33; B = 8'hA0; #100;
A = 8'h33; B = 8'hA1; #100;
A = 8'h33; B = 8'hA2; #100;
A = 8'h33; B = 8'hA3; #100;
A = 8'h33; B = 8'hA4; #100;
A = 8'h33; B = 8'hA5; #100;
A = 8'h33; B = 8'hA6; #100;
A = 8'h33; B = 8'hA7; #100;
A = 8'h33; B = 8'hA8; #100;
A = 8'h33; B = 8'hA9; #100;
A = 8'h33; B = 8'hAA; #100;
A = 8'h33; B = 8'hAB; #100;
A = 8'h33; B = 8'hAC; #100;
A = 8'h33; B = 8'hAD; #100;
A = 8'h33; B = 8'hAE; #100;
A = 8'h33; B = 8'hAF; #100;
A = 8'h33; B = 8'hB0; #100;
A = 8'h33; B = 8'hB1; #100;
A = 8'h33; B = 8'hB2; #100;
A = 8'h33; B = 8'hB3; #100;
A = 8'h33; B = 8'hB4; #100;
A = 8'h33; B = 8'hB5; #100;
A = 8'h33; B = 8'hB6; #100;
A = 8'h33; B = 8'hB7; #100;
A = 8'h33; B = 8'hB8; #100;
A = 8'h33; B = 8'hB9; #100;
A = 8'h33; B = 8'hBA; #100;
A = 8'h33; B = 8'hBB; #100;
A = 8'h33; B = 8'hBC; #100;
A = 8'h33; B = 8'hBD; #100;
A = 8'h33; B = 8'hBE; #100;
A = 8'h33; B = 8'hBF; #100;
A = 8'h33; B = 8'hC0; #100;
A = 8'h33; B = 8'hC1; #100;
A = 8'h33; B = 8'hC2; #100;
A = 8'h33; B = 8'hC3; #100;
A = 8'h33; B = 8'hC4; #100;
A = 8'h33; B = 8'hC5; #100;
A = 8'h33; B = 8'hC6; #100;
A = 8'h33; B = 8'hC7; #100;
A = 8'h33; B = 8'hC8; #100;
A = 8'h33; B = 8'hC9; #100;
A = 8'h33; B = 8'hCA; #100;
A = 8'h33; B = 8'hCB; #100;
A = 8'h33; B = 8'hCC; #100;
A = 8'h33; B = 8'hCD; #100;
A = 8'h33; B = 8'hCE; #100;
A = 8'h33; B = 8'hCF; #100;
A = 8'h33; B = 8'hD0; #100;
A = 8'h33; B = 8'hD1; #100;
A = 8'h33; B = 8'hD2; #100;
A = 8'h33; B = 8'hD3; #100;
A = 8'h33; B = 8'hD4; #100;
A = 8'h33; B = 8'hD5; #100;
A = 8'h33; B = 8'hD6; #100;
A = 8'h33; B = 8'hD7; #100;
A = 8'h33; B = 8'hD8; #100;
A = 8'h33; B = 8'hD9; #100;
A = 8'h33; B = 8'hDA; #100;
A = 8'h33; B = 8'hDB; #100;
A = 8'h33; B = 8'hDC; #100;
A = 8'h33; B = 8'hDD; #100;
A = 8'h33; B = 8'hDE; #100;
A = 8'h33; B = 8'hDF; #100;
A = 8'h33; B = 8'hE0; #100;
A = 8'h33; B = 8'hE1; #100;
A = 8'h33; B = 8'hE2; #100;
A = 8'h33; B = 8'hE3; #100;
A = 8'h33; B = 8'hE4; #100;
A = 8'h33; B = 8'hE5; #100;
A = 8'h33; B = 8'hE6; #100;
A = 8'h33; B = 8'hE7; #100;
A = 8'h33; B = 8'hE8; #100;
A = 8'h33; B = 8'hE9; #100;
A = 8'h33; B = 8'hEA; #100;
A = 8'h33; B = 8'hEB; #100;
A = 8'h33; B = 8'hEC; #100;
A = 8'h33; B = 8'hED; #100;
A = 8'h33; B = 8'hEE; #100;
A = 8'h33; B = 8'hEF; #100;
A = 8'h33; B = 8'hF0; #100;
A = 8'h33; B = 8'hF1; #100;
A = 8'h33; B = 8'hF2; #100;
A = 8'h33; B = 8'hF3; #100;
A = 8'h33; B = 8'hF4; #100;
A = 8'h33; B = 8'hF5; #100;
A = 8'h33; B = 8'hF6; #100;
A = 8'h33; B = 8'hF7; #100;
A = 8'h33; B = 8'hF8; #100;
A = 8'h33; B = 8'hF9; #100;
A = 8'h33; B = 8'hFA; #100;
A = 8'h33; B = 8'hFB; #100;
A = 8'h33; B = 8'hFC; #100;
A = 8'h33; B = 8'hFD; #100;
A = 8'h33; B = 8'hFE; #100;
A = 8'h33; B = 8'hFF; #100;
A = 8'h34; B = 8'h0; #100;
A = 8'h34; B = 8'h1; #100;
A = 8'h34; B = 8'h2; #100;
A = 8'h34; B = 8'h3; #100;
A = 8'h34; B = 8'h4; #100;
A = 8'h34; B = 8'h5; #100;
A = 8'h34; B = 8'h6; #100;
A = 8'h34; B = 8'h7; #100;
A = 8'h34; B = 8'h8; #100;
A = 8'h34; B = 8'h9; #100;
A = 8'h34; B = 8'hA; #100;
A = 8'h34; B = 8'hB; #100;
A = 8'h34; B = 8'hC; #100;
A = 8'h34; B = 8'hD; #100;
A = 8'h34; B = 8'hE; #100;
A = 8'h34; B = 8'hF; #100;
A = 8'h34; B = 8'h10; #100;
A = 8'h34; B = 8'h11; #100;
A = 8'h34; B = 8'h12; #100;
A = 8'h34; B = 8'h13; #100;
A = 8'h34; B = 8'h14; #100;
A = 8'h34; B = 8'h15; #100;
A = 8'h34; B = 8'h16; #100;
A = 8'h34; B = 8'h17; #100;
A = 8'h34; B = 8'h18; #100;
A = 8'h34; B = 8'h19; #100;
A = 8'h34; B = 8'h1A; #100;
A = 8'h34; B = 8'h1B; #100;
A = 8'h34; B = 8'h1C; #100;
A = 8'h34; B = 8'h1D; #100;
A = 8'h34; B = 8'h1E; #100;
A = 8'h34; B = 8'h1F; #100;
A = 8'h34; B = 8'h20; #100;
A = 8'h34; B = 8'h21; #100;
A = 8'h34; B = 8'h22; #100;
A = 8'h34; B = 8'h23; #100;
A = 8'h34; B = 8'h24; #100;
A = 8'h34; B = 8'h25; #100;
A = 8'h34; B = 8'h26; #100;
A = 8'h34; B = 8'h27; #100;
A = 8'h34; B = 8'h28; #100;
A = 8'h34; B = 8'h29; #100;
A = 8'h34; B = 8'h2A; #100;
A = 8'h34; B = 8'h2B; #100;
A = 8'h34; B = 8'h2C; #100;
A = 8'h34; B = 8'h2D; #100;
A = 8'h34; B = 8'h2E; #100;
A = 8'h34; B = 8'h2F; #100;
A = 8'h34; B = 8'h30; #100;
A = 8'h34; B = 8'h31; #100;
A = 8'h34; B = 8'h32; #100;
A = 8'h34; B = 8'h33; #100;
A = 8'h34; B = 8'h34; #100;
A = 8'h34; B = 8'h35; #100;
A = 8'h34; B = 8'h36; #100;
A = 8'h34; B = 8'h37; #100;
A = 8'h34; B = 8'h38; #100;
A = 8'h34; B = 8'h39; #100;
A = 8'h34; B = 8'h3A; #100;
A = 8'h34; B = 8'h3B; #100;
A = 8'h34; B = 8'h3C; #100;
A = 8'h34; B = 8'h3D; #100;
A = 8'h34; B = 8'h3E; #100;
A = 8'h34; B = 8'h3F; #100;
A = 8'h34; B = 8'h40; #100;
A = 8'h34; B = 8'h41; #100;
A = 8'h34; B = 8'h42; #100;
A = 8'h34; B = 8'h43; #100;
A = 8'h34; B = 8'h44; #100;
A = 8'h34; B = 8'h45; #100;
A = 8'h34; B = 8'h46; #100;
A = 8'h34; B = 8'h47; #100;
A = 8'h34; B = 8'h48; #100;
A = 8'h34; B = 8'h49; #100;
A = 8'h34; B = 8'h4A; #100;
A = 8'h34; B = 8'h4B; #100;
A = 8'h34; B = 8'h4C; #100;
A = 8'h34; B = 8'h4D; #100;
A = 8'h34; B = 8'h4E; #100;
A = 8'h34; B = 8'h4F; #100;
A = 8'h34; B = 8'h50; #100;
A = 8'h34; B = 8'h51; #100;
A = 8'h34; B = 8'h52; #100;
A = 8'h34; B = 8'h53; #100;
A = 8'h34; B = 8'h54; #100;
A = 8'h34; B = 8'h55; #100;
A = 8'h34; B = 8'h56; #100;
A = 8'h34; B = 8'h57; #100;
A = 8'h34; B = 8'h58; #100;
A = 8'h34; B = 8'h59; #100;
A = 8'h34; B = 8'h5A; #100;
A = 8'h34; B = 8'h5B; #100;
A = 8'h34; B = 8'h5C; #100;
A = 8'h34; B = 8'h5D; #100;
A = 8'h34; B = 8'h5E; #100;
A = 8'h34; B = 8'h5F; #100;
A = 8'h34; B = 8'h60; #100;
A = 8'h34; B = 8'h61; #100;
A = 8'h34; B = 8'h62; #100;
A = 8'h34; B = 8'h63; #100;
A = 8'h34; B = 8'h64; #100;
A = 8'h34; B = 8'h65; #100;
A = 8'h34; B = 8'h66; #100;
A = 8'h34; B = 8'h67; #100;
A = 8'h34; B = 8'h68; #100;
A = 8'h34; B = 8'h69; #100;
A = 8'h34; B = 8'h6A; #100;
A = 8'h34; B = 8'h6B; #100;
A = 8'h34; B = 8'h6C; #100;
A = 8'h34; B = 8'h6D; #100;
A = 8'h34; B = 8'h6E; #100;
A = 8'h34; B = 8'h6F; #100;
A = 8'h34; B = 8'h70; #100;
A = 8'h34; B = 8'h71; #100;
A = 8'h34; B = 8'h72; #100;
A = 8'h34; B = 8'h73; #100;
A = 8'h34; B = 8'h74; #100;
A = 8'h34; B = 8'h75; #100;
A = 8'h34; B = 8'h76; #100;
A = 8'h34; B = 8'h77; #100;
A = 8'h34; B = 8'h78; #100;
A = 8'h34; B = 8'h79; #100;
A = 8'h34; B = 8'h7A; #100;
A = 8'h34; B = 8'h7B; #100;
A = 8'h34; B = 8'h7C; #100;
A = 8'h34; B = 8'h7D; #100;
A = 8'h34; B = 8'h7E; #100;
A = 8'h34; B = 8'h7F; #100;
A = 8'h34; B = 8'h80; #100;
A = 8'h34; B = 8'h81; #100;
A = 8'h34; B = 8'h82; #100;
A = 8'h34; B = 8'h83; #100;
A = 8'h34; B = 8'h84; #100;
A = 8'h34; B = 8'h85; #100;
A = 8'h34; B = 8'h86; #100;
A = 8'h34; B = 8'h87; #100;
A = 8'h34; B = 8'h88; #100;
A = 8'h34; B = 8'h89; #100;
A = 8'h34; B = 8'h8A; #100;
A = 8'h34; B = 8'h8B; #100;
A = 8'h34; B = 8'h8C; #100;
A = 8'h34; B = 8'h8D; #100;
A = 8'h34; B = 8'h8E; #100;
A = 8'h34; B = 8'h8F; #100;
A = 8'h34; B = 8'h90; #100;
A = 8'h34; B = 8'h91; #100;
A = 8'h34; B = 8'h92; #100;
A = 8'h34; B = 8'h93; #100;
A = 8'h34; B = 8'h94; #100;
A = 8'h34; B = 8'h95; #100;
A = 8'h34; B = 8'h96; #100;
A = 8'h34; B = 8'h97; #100;
A = 8'h34; B = 8'h98; #100;
A = 8'h34; B = 8'h99; #100;
A = 8'h34; B = 8'h9A; #100;
A = 8'h34; B = 8'h9B; #100;
A = 8'h34; B = 8'h9C; #100;
A = 8'h34; B = 8'h9D; #100;
A = 8'h34; B = 8'h9E; #100;
A = 8'h34; B = 8'h9F; #100;
A = 8'h34; B = 8'hA0; #100;
A = 8'h34; B = 8'hA1; #100;
A = 8'h34; B = 8'hA2; #100;
A = 8'h34; B = 8'hA3; #100;
A = 8'h34; B = 8'hA4; #100;
A = 8'h34; B = 8'hA5; #100;
A = 8'h34; B = 8'hA6; #100;
A = 8'h34; B = 8'hA7; #100;
A = 8'h34; B = 8'hA8; #100;
A = 8'h34; B = 8'hA9; #100;
A = 8'h34; B = 8'hAA; #100;
A = 8'h34; B = 8'hAB; #100;
A = 8'h34; B = 8'hAC; #100;
A = 8'h34; B = 8'hAD; #100;
A = 8'h34; B = 8'hAE; #100;
A = 8'h34; B = 8'hAF; #100;
A = 8'h34; B = 8'hB0; #100;
A = 8'h34; B = 8'hB1; #100;
A = 8'h34; B = 8'hB2; #100;
A = 8'h34; B = 8'hB3; #100;
A = 8'h34; B = 8'hB4; #100;
A = 8'h34; B = 8'hB5; #100;
A = 8'h34; B = 8'hB6; #100;
A = 8'h34; B = 8'hB7; #100;
A = 8'h34; B = 8'hB8; #100;
A = 8'h34; B = 8'hB9; #100;
A = 8'h34; B = 8'hBA; #100;
A = 8'h34; B = 8'hBB; #100;
A = 8'h34; B = 8'hBC; #100;
A = 8'h34; B = 8'hBD; #100;
A = 8'h34; B = 8'hBE; #100;
A = 8'h34; B = 8'hBF; #100;
A = 8'h34; B = 8'hC0; #100;
A = 8'h34; B = 8'hC1; #100;
A = 8'h34; B = 8'hC2; #100;
A = 8'h34; B = 8'hC3; #100;
A = 8'h34; B = 8'hC4; #100;
A = 8'h34; B = 8'hC5; #100;
A = 8'h34; B = 8'hC6; #100;
A = 8'h34; B = 8'hC7; #100;
A = 8'h34; B = 8'hC8; #100;
A = 8'h34; B = 8'hC9; #100;
A = 8'h34; B = 8'hCA; #100;
A = 8'h34; B = 8'hCB; #100;
A = 8'h34; B = 8'hCC; #100;
A = 8'h34; B = 8'hCD; #100;
A = 8'h34; B = 8'hCE; #100;
A = 8'h34; B = 8'hCF; #100;
A = 8'h34; B = 8'hD0; #100;
A = 8'h34; B = 8'hD1; #100;
A = 8'h34; B = 8'hD2; #100;
A = 8'h34; B = 8'hD3; #100;
A = 8'h34; B = 8'hD4; #100;
A = 8'h34; B = 8'hD5; #100;
A = 8'h34; B = 8'hD6; #100;
A = 8'h34; B = 8'hD7; #100;
A = 8'h34; B = 8'hD8; #100;
A = 8'h34; B = 8'hD9; #100;
A = 8'h34; B = 8'hDA; #100;
A = 8'h34; B = 8'hDB; #100;
A = 8'h34; B = 8'hDC; #100;
A = 8'h34; B = 8'hDD; #100;
A = 8'h34; B = 8'hDE; #100;
A = 8'h34; B = 8'hDF; #100;
A = 8'h34; B = 8'hE0; #100;
A = 8'h34; B = 8'hE1; #100;
A = 8'h34; B = 8'hE2; #100;
A = 8'h34; B = 8'hE3; #100;
A = 8'h34; B = 8'hE4; #100;
A = 8'h34; B = 8'hE5; #100;
A = 8'h34; B = 8'hE6; #100;
A = 8'h34; B = 8'hE7; #100;
A = 8'h34; B = 8'hE8; #100;
A = 8'h34; B = 8'hE9; #100;
A = 8'h34; B = 8'hEA; #100;
A = 8'h34; B = 8'hEB; #100;
A = 8'h34; B = 8'hEC; #100;
A = 8'h34; B = 8'hED; #100;
A = 8'h34; B = 8'hEE; #100;
A = 8'h34; B = 8'hEF; #100;
A = 8'h34; B = 8'hF0; #100;
A = 8'h34; B = 8'hF1; #100;
A = 8'h34; B = 8'hF2; #100;
A = 8'h34; B = 8'hF3; #100;
A = 8'h34; B = 8'hF4; #100;
A = 8'h34; B = 8'hF5; #100;
A = 8'h34; B = 8'hF6; #100;
A = 8'h34; B = 8'hF7; #100;
A = 8'h34; B = 8'hF8; #100;
A = 8'h34; B = 8'hF9; #100;
A = 8'h34; B = 8'hFA; #100;
A = 8'h34; B = 8'hFB; #100;
A = 8'h34; B = 8'hFC; #100;
A = 8'h34; B = 8'hFD; #100;
A = 8'h34; B = 8'hFE; #100;
A = 8'h34; B = 8'hFF; #100;
A = 8'h35; B = 8'h0; #100;
A = 8'h35; B = 8'h1; #100;
A = 8'h35; B = 8'h2; #100;
A = 8'h35; B = 8'h3; #100;
A = 8'h35; B = 8'h4; #100;
A = 8'h35; B = 8'h5; #100;
A = 8'h35; B = 8'h6; #100;
A = 8'h35; B = 8'h7; #100;
A = 8'h35; B = 8'h8; #100;
A = 8'h35; B = 8'h9; #100;
A = 8'h35; B = 8'hA; #100;
A = 8'h35; B = 8'hB; #100;
A = 8'h35; B = 8'hC; #100;
A = 8'h35; B = 8'hD; #100;
A = 8'h35; B = 8'hE; #100;
A = 8'h35; B = 8'hF; #100;
A = 8'h35; B = 8'h10; #100;
A = 8'h35; B = 8'h11; #100;
A = 8'h35; B = 8'h12; #100;
A = 8'h35; B = 8'h13; #100;
A = 8'h35; B = 8'h14; #100;
A = 8'h35; B = 8'h15; #100;
A = 8'h35; B = 8'h16; #100;
A = 8'h35; B = 8'h17; #100;
A = 8'h35; B = 8'h18; #100;
A = 8'h35; B = 8'h19; #100;
A = 8'h35; B = 8'h1A; #100;
A = 8'h35; B = 8'h1B; #100;
A = 8'h35; B = 8'h1C; #100;
A = 8'h35; B = 8'h1D; #100;
A = 8'h35; B = 8'h1E; #100;
A = 8'h35; B = 8'h1F; #100;
A = 8'h35; B = 8'h20; #100;
A = 8'h35; B = 8'h21; #100;
A = 8'h35; B = 8'h22; #100;
A = 8'h35; B = 8'h23; #100;
A = 8'h35; B = 8'h24; #100;
A = 8'h35; B = 8'h25; #100;
A = 8'h35; B = 8'h26; #100;
A = 8'h35; B = 8'h27; #100;
A = 8'h35; B = 8'h28; #100;
A = 8'h35; B = 8'h29; #100;
A = 8'h35; B = 8'h2A; #100;
A = 8'h35; B = 8'h2B; #100;
A = 8'h35; B = 8'h2C; #100;
A = 8'h35; B = 8'h2D; #100;
A = 8'h35; B = 8'h2E; #100;
A = 8'h35; B = 8'h2F; #100;
A = 8'h35; B = 8'h30; #100;
A = 8'h35; B = 8'h31; #100;
A = 8'h35; B = 8'h32; #100;
A = 8'h35; B = 8'h33; #100;
A = 8'h35; B = 8'h34; #100;
A = 8'h35; B = 8'h35; #100;
A = 8'h35; B = 8'h36; #100;
A = 8'h35; B = 8'h37; #100;
A = 8'h35; B = 8'h38; #100;
A = 8'h35; B = 8'h39; #100;
A = 8'h35; B = 8'h3A; #100;
A = 8'h35; B = 8'h3B; #100;
A = 8'h35; B = 8'h3C; #100;
A = 8'h35; B = 8'h3D; #100;
A = 8'h35; B = 8'h3E; #100;
A = 8'h35; B = 8'h3F; #100;
A = 8'h35; B = 8'h40; #100;
A = 8'h35; B = 8'h41; #100;
A = 8'h35; B = 8'h42; #100;
A = 8'h35; B = 8'h43; #100;
A = 8'h35; B = 8'h44; #100;
A = 8'h35; B = 8'h45; #100;
A = 8'h35; B = 8'h46; #100;
A = 8'h35; B = 8'h47; #100;
A = 8'h35; B = 8'h48; #100;
A = 8'h35; B = 8'h49; #100;
A = 8'h35; B = 8'h4A; #100;
A = 8'h35; B = 8'h4B; #100;
A = 8'h35; B = 8'h4C; #100;
A = 8'h35; B = 8'h4D; #100;
A = 8'h35; B = 8'h4E; #100;
A = 8'h35; B = 8'h4F; #100;
A = 8'h35; B = 8'h50; #100;
A = 8'h35; B = 8'h51; #100;
A = 8'h35; B = 8'h52; #100;
A = 8'h35; B = 8'h53; #100;
A = 8'h35; B = 8'h54; #100;
A = 8'h35; B = 8'h55; #100;
A = 8'h35; B = 8'h56; #100;
A = 8'h35; B = 8'h57; #100;
A = 8'h35; B = 8'h58; #100;
A = 8'h35; B = 8'h59; #100;
A = 8'h35; B = 8'h5A; #100;
A = 8'h35; B = 8'h5B; #100;
A = 8'h35; B = 8'h5C; #100;
A = 8'h35; B = 8'h5D; #100;
A = 8'h35; B = 8'h5E; #100;
A = 8'h35; B = 8'h5F; #100;
A = 8'h35; B = 8'h60; #100;
A = 8'h35; B = 8'h61; #100;
A = 8'h35; B = 8'h62; #100;
A = 8'h35; B = 8'h63; #100;
A = 8'h35; B = 8'h64; #100;
A = 8'h35; B = 8'h65; #100;
A = 8'h35; B = 8'h66; #100;
A = 8'h35; B = 8'h67; #100;
A = 8'h35; B = 8'h68; #100;
A = 8'h35; B = 8'h69; #100;
A = 8'h35; B = 8'h6A; #100;
A = 8'h35; B = 8'h6B; #100;
A = 8'h35; B = 8'h6C; #100;
A = 8'h35; B = 8'h6D; #100;
A = 8'h35; B = 8'h6E; #100;
A = 8'h35; B = 8'h6F; #100;
A = 8'h35; B = 8'h70; #100;
A = 8'h35; B = 8'h71; #100;
A = 8'h35; B = 8'h72; #100;
A = 8'h35; B = 8'h73; #100;
A = 8'h35; B = 8'h74; #100;
A = 8'h35; B = 8'h75; #100;
A = 8'h35; B = 8'h76; #100;
A = 8'h35; B = 8'h77; #100;
A = 8'h35; B = 8'h78; #100;
A = 8'h35; B = 8'h79; #100;
A = 8'h35; B = 8'h7A; #100;
A = 8'h35; B = 8'h7B; #100;
A = 8'h35; B = 8'h7C; #100;
A = 8'h35; B = 8'h7D; #100;
A = 8'h35; B = 8'h7E; #100;
A = 8'h35; B = 8'h7F; #100;
A = 8'h35; B = 8'h80; #100;
A = 8'h35; B = 8'h81; #100;
A = 8'h35; B = 8'h82; #100;
A = 8'h35; B = 8'h83; #100;
A = 8'h35; B = 8'h84; #100;
A = 8'h35; B = 8'h85; #100;
A = 8'h35; B = 8'h86; #100;
A = 8'h35; B = 8'h87; #100;
A = 8'h35; B = 8'h88; #100;
A = 8'h35; B = 8'h89; #100;
A = 8'h35; B = 8'h8A; #100;
A = 8'h35; B = 8'h8B; #100;
A = 8'h35; B = 8'h8C; #100;
A = 8'h35; B = 8'h8D; #100;
A = 8'h35; B = 8'h8E; #100;
A = 8'h35; B = 8'h8F; #100;
A = 8'h35; B = 8'h90; #100;
A = 8'h35; B = 8'h91; #100;
A = 8'h35; B = 8'h92; #100;
A = 8'h35; B = 8'h93; #100;
A = 8'h35; B = 8'h94; #100;
A = 8'h35; B = 8'h95; #100;
A = 8'h35; B = 8'h96; #100;
A = 8'h35; B = 8'h97; #100;
A = 8'h35; B = 8'h98; #100;
A = 8'h35; B = 8'h99; #100;
A = 8'h35; B = 8'h9A; #100;
A = 8'h35; B = 8'h9B; #100;
A = 8'h35; B = 8'h9C; #100;
A = 8'h35; B = 8'h9D; #100;
A = 8'h35; B = 8'h9E; #100;
A = 8'h35; B = 8'h9F; #100;
A = 8'h35; B = 8'hA0; #100;
A = 8'h35; B = 8'hA1; #100;
A = 8'h35; B = 8'hA2; #100;
A = 8'h35; B = 8'hA3; #100;
A = 8'h35; B = 8'hA4; #100;
A = 8'h35; B = 8'hA5; #100;
A = 8'h35; B = 8'hA6; #100;
A = 8'h35; B = 8'hA7; #100;
A = 8'h35; B = 8'hA8; #100;
A = 8'h35; B = 8'hA9; #100;
A = 8'h35; B = 8'hAA; #100;
A = 8'h35; B = 8'hAB; #100;
A = 8'h35; B = 8'hAC; #100;
A = 8'h35; B = 8'hAD; #100;
A = 8'h35; B = 8'hAE; #100;
A = 8'h35; B = 8'hAF; #100;
A = 8'h35; B = 8'hB0; #100;
A = 8'h35; B = 8'hB1; #100;
A = 8'h35; B = 8'hB2; #100;
A = 8'h35; B = 8'hB3; #100;
A = 8'h35; B = 8'hB4; #100;
A = 8'h35; B = 8'hB5; #100;
A = 8'h35; B = 8'hB6; #100;
A = 8'h35; B = 8'hB7; #100;
A = 8'h35; B = 8'hB8; #100;
A = 8'h35; B = 8'hB9; #100;
A = 8'h35; B = 8'hBA; #100;
A = 8'h35; B = 8'hBB; #100;
A = 8'h35; B = 8'hBC; #100;
A = 8'h35; B = 8'hBD; #100;
A = 8'h35; B = 8'hBE; #100;
A = 8'h35; B = 8'hBF; #100;
A = 8'h35; B = 8'hC0; #100;
A = 8'h35; B = 8'hC1; #100;
A = 8'h35; B = 8'hC2; #100;
A = 8'h35; B = 8'hC3; #100;
A = 8'h35; B = 8'hC4; #100;
A = 8'h35; B = 8'hC5; #100;
A = 8'h35; B = 8'hC6; #100;
A = 8'h35; B = 8'hC7; #100;
A = 8'h35; B = 8'hC8; #100;
A = 8'h35; B = 8'hC9; #100;
A = 8'h35; B = 8'hCA; #100;
A = 8'h35; B = 8'hCB; #100;
A = 8'h35; B = 8'hCC; #100;
A = 8'h35; B = 8'hCD; #100;
A = 8'h35; B = 8'hCE; #100;
A = 8'h35; B = 8'hCF; #100;
A = 8'h35; B = 8'hD0; #100;
A = 8'h35; B = 8'hD1; #100;
A = 8'h35; B = 8'hD2; #100;
A = 8'h35; B = 8'hD3; #100;
A = 8'h35; B = 8'hD4; #100;
A = 8'h35; B = 8'hD5; #100;
A = 8'h35; B = 8'hD6; #100;
A = 8'h35; B = 8'hD7; #100;
A = 8'h35; B = 8'hD8; #100;
A = 8'h35; B = 8'hD9; #100;
A = 8'h35; B = 8'hDA; #100;
A = 8'h35; B = 8'hDB; #100;
A = 8'h35; B = 8'hDC; #100;
A = 8'h35; B = 8'hDD; #100;
A = 8'h35; B = 8'hDE; #100;
A = 8'h35; B = 8'hDF; #100;
A = 8'h35; B = 8'hE0; #100;
A = 8'h35; B = 8'hE1; #100;
A = 8'h35; B = 8'hE2; #100;
A = 8'h35; B = 8'hE3; #100;
A = 8'h35; B = 8'hE4; #100;
A = 8'h35; B = 8'hE5; #100;
A = 8'h35; B = 8'hE6; #100;
A = 8'h35; B = 8'hE7; #100;
A = 8'h35; B = 8'hE8; #100;
A = 8'h35; B = 8'hE9; #100;
A = 8'h35; B = 8'hEA; #100;
A = 8'h35; B = 8'hEB; #100;
A = 8'h35; B = 8'hEC; #100;
A = 8'h35; B = 8'hED; #100;
A = 8'h35; B = 8'hEE; #100;
A = 8'h35; B = 8'hEF; #100;
A = 8'h35; B = 8'hF0; #100;
A = 8'h35; B = 8'hF1; #100;
A = 8'h35; B = 8'hF2; #100;
A = 8'h35; B = 8'hF3; #100;
A = 8'h35; B = 8'hF4; #100;
A = 8'h35; B = 8'hF5; #100;
A = 8'h35; B = 8'hF6; #100;
A = 8'h35; B = 8'hF7; #100;
A = 8'h35; B = 8'hF8; #100;
A = 8'h35; B = 8'hF9; #100;
A = 8'h35; B = 8'hFA; #100;
A = 8'h35; B = 8'hFB; #100;
A = 8'h35; B = 8'hFC; #100;
A = 8'h35; B = 8'hFD; #100;
A = 8'h35; B = 8'hFE; #100;
A = 8'h35; B = 8'hFF; #100;
A = 8'h36; B = 8'h0; #100;
A = 8'h36; B = 8'h1; #100;
A = 8'h36; B = 8'h2; #100;
A = 8'h36; B = 8'h3; #100;
A = 8'h36; B = 8'h4; #100;
A = 8'h36; B = 8'h5; #100;
A = 8'h36; B = 8'h6; #100;
A = 8'h36; B = 8'h7; #100;
A = 8'h36; B = 8'h8; #100;
A = 8'h36; B = 8'h9; #100;
A = 8'h36; B = 8'hA; #100;
A = 8'h36; B = 8'hB; #100;
A = 8'h36; B = 8'hC; #100;
A = 8'h36; B = 8'hD; #100;
A = 8'h36; B = 8'hE; #100;
A = 8'h36; B = 8'hF; #100;
A = 8'h36; B = 8'h10; #100;
A = 8'h36; B = 8'h11; #100;
A = 8'h36; B = 8'h12; #100;
A = 8'h36; B = 8'h13; #100;
A = 8'h36; B = 8'h14; #100;
A = 8'h36; B = 8'h15; #100;
A = 8'h36; B = 8'h16; #100;
A = 8'h36; B = 8'h17; #100;
A = 8'h36; B = 8'h18; #100;
A = 8'h36; B = 8'h19; #100;
A = 8'h36; B = 8'h1A; #100;
A = 8'h36; B = 8'h1B; #100;
A = 8'h36; B = 8'h1C; #100;
A = 8'h36; B = 8'h1D; #100;
A = 8'h36; B = 8'h1E; #100;
A = 8'h36; B = 8'h1F; #100;
A = 8'h36; B = 8'h20; #100;
A = 8'h36; B = 8'h21; #100;
A = 8'h36; B = 8'h22; #100;
A = 8'h36; B = 8'h23; #100;
A = 8'h36; B = 8'h24; #100;
A = 8'h36; B = 8'h25; #100;
A = 8'h36; B = 8'h26; #100;
A = 8'h36; B = 8'h27; #100;
A = 8'h36; B = 8'h28; #100;
A = 8'h36; B = 8'h29; #100;
A = 8'h36; B = 8'h2A; #100;
A = 8'h36; B = 8'h2B; #100;
A = 8'h36; B = 8'h2C; #100;
A = 8'h36; B = 8'h2D; #100;
A = 8'h36; B = 8'h2E; #100;
A = 8'h36; B = 8'h2F; #100;
A = 8'h36; B = 8'h30; #100;
A = 8'h36; B = 8'h31; #100;
A = 8'h36; B = 8'h32; #100;
A = 8'h36; B = 8'h33; #100;
A = 8'h36; B = 8'h34; #100;
A = 8'h36; B = 8'h35; #100;
A = 8'h36; B = 8'h36; #100;
A = 8'h36; B = 8'h37; #100;
A = 8'h36; B = 8'h38; #100;
A = 8'h36; B = 8'h39; #100;
A = 8'h36; B = 8'h3A; #100;
A = 8'h36; B = 8'h3B; #100;
A = 8'h36; B = 8'h3C; #100;
A = 8'h36; B = 8'h3D; #100;
A = 8'h36; B = 8'h3E; #100;
A = 8'h36; B = 8'h3F; #100;
A = 8'h36; B = 8'h40; #100;
A = 8'h36; B = 8'h41; #100;
A = 8'h36; B = 8'h42; #100;
A = 8'h36; B = 8'h43; #100;
A = 8'h36; B = 8'h44; #100;
A = 8'h36; B = 8'h45; #100;
A = 8'h36; B = 8'h46; #100;
A = 8'h36; B = 8'h47; #100;
A = 8'h36; B = 8'h48; #100;
A = 8'h36; B = 8'h49; #100;
A = 8'h36; B = 8'h4A; #100;
A = 8'h36; B = 8'h4B; #100;
A = 8'h36; B = 8'h4C; #100;
A = 8'h36; B = 8'h4D; #100;
A = 8'h36; B = 8'h4E; #100;
A = 8'h36; B = 8'h4F; #100;
A = 8'h36; B = 8'h50; #100;
A = 8'h36; B = 8'h51; #100;
A = 8'h36; B = 8'h52; #100;
A = 8'h36; B = 8'h53; #100;
A = 8'h36; B = 8'h54; #100;
A = 8'h36; B = 8'h55; #100;
A = 8'h36; B = 8'h56; #100;
A = 8'h36; B = 8'h57; #100;
A = 8'h36; B = 8'h58; #100;
A = 8'h36; B = 8'h59; #100;
A = 8'h36; B = 8'h5A; #100;
A = 8'h36; B = 8'h5B; #100;
A = 8'h36; B = 8'h5C; #100;
A = 8'h36; B = 8'h5D; #100;
A = 8'h36; B = 8'h5E; #100;
A = 8'h36; B = 8'h5F; #100;
A = 8'h36; B = 8'h60; #100;
A = 8'h36; B = 8'h61; #100;
A = 8'h36; B = 8'h62; #100;
A = 8'h36; B = 8'h63; #100;
A = 8'h36; B = 8'h64; #100;
A = 8'h36; B = 8'h65; #100;
A = 8'h36; B = 8'h66; #100;
A = 8'h36; B = 8'h67; #100;
A = 8'h36; B = 8'h68; #100;
A = 8'h36; B = 8'h69; #100;
A = 8'h36; B = 8'h6A; #100;
A = 8'h36; B = 8'h6B; #100;
A = 8'h36; B = 8'h6C; #100;
A = 8'h36; B = 8'h6D; #100;
A = 8'h36; B = 8'h6E; #100;
A = 8'h36; B = 8'h6F; #100;
A = 8'h36; B = 8'h70; #100;
A = 8'h36; B = 8'h71; #100;
A = 8'h36; B = 8'h72; #100;
A = 8'h36; B = 8'h73; #100;
A = 8'h36; B = 8'h74; #100;
A = 8'h36; B = 8'h75; #100;
A = 8'h36; B = 8'h76; #100;
A = 8'h36; B = 8'h77; #100;
A = 8'h36; B = 8'h78; #100;
A = 8'h36; B = 8'h79; #100;
A = 8'h36; B = 8'h7A; #100;
A = 8'h36; B = 8'h7B; #100;
A = 8'h36; B = 8'h7C; #100;
A = 8'h36; B = 8'h7D; #100;
A = 8'h36; B = 8'h7E; #100;
A = 8'h36; B = 8'h7F; #100;
A = 8'h36; B = 8'h80; #100;
A = 8'h36; B = 8'h81; #100;
A = 8'h36; B = 8'h82; #100;
A = 8'h36; B = 8'h83; #100;
A = 8'h36; B = 8'h84; #100;
A = 8'h36; B = 8'h85; #100;
A = 8'h36; B = 8'h86; #100;
A = 8'h36; B = 8'h87; #100;
A = 8'h36; B = 8'h88; #100;
A = 8'h36; B = 8'h89; #100;
A = 8'h36; B = 8'h8A; #100;
A = 8'h36; B = 8'h8B; #100;
A = 8'h36; B = 8'h8C; #100;
A = 8'h36; B = 8'h8D; #100;
A = 8'h36; B = 8'h8E; #100;
A = 8'h36; B = 8'h8F; #100;
A = 8'h36; B = 8'h90; #100;
A = 8'h36; B = 8'h91; #100;
A = 8'h36; B = 8'h92; #100;
A = 8'h36; B = 8'h93; #100;
A = 8'h36; B = 8'h94; #100;
A = 8'h36; B = 8'h95; #100;
A = 8'h36; B = 8'h96; #100;
A = 8'h36; B = 8'h97; #100;
A = 8'h36; B = 8'h98; #100;
A = 8'h36; B = 8'h99; #100;
A = 8'h36; B = 8'h9A; #100;
A = 8'h36; B = 8'h9B; #100;
A = 8'h36; B = 8'h9C; #100;
A = 8'h36; B = 8'h9D; #100;
A = 8'h36; B = 8'h9E; #100;
A = 8'h36; B = 8'h9F; #100;
A = 8'h36; B = 8'hA0; #100;
A = 8'h36; B = 8'hA1; #100;
A = 8'h36; B = 8'hA2; #100;
A = 8'h36; B = 8'hA3; #100;
A = 8'h36; B = 8'hA4; #100;
A = 8'h36; B = 8'hA5; #100;
A = 8'h36; B = 8'hA6; #100;
A = 8'h36; B = 8'hA7; #100;
A = 8'h36; B = 8'hA8; #100;
A = 8'h36; B = 8'hA9; #100;
A = 8'h36; B = 8'hAA; #100;
A = 8'h36; B = 8'hAB; #100;
A = 8'h36; B = 8'hAC; #100;
A = 8'h36; B = 8'hAD; #100;
A = 8'h36; B = 8'hAE; #100;
A = 8'h36; B = 8'hAF; #100;
A = 8'h36; B = 8'hB0; #100;
A = 8'h36; B = 8'hB1; #100;
A = 8'h36; B = 8'hB2; #100;
A = 8'h36; B = 8'hB3; #100;
A = 8'h36; B = 8'hB4; #100;
A = 8'h36; B = 8'hB5; #100;
A = 8'h36; B = 8'hB6; #100;
A = 8'h36; B = 8'hB7; #100;
A = 8'h36; B = 8'hB8; #100;
A = 8'h36; B = 8'hB9; #100;
A = 8'h36; B = 8'hBA; #100;
A = 8'h36; B = 8'hBB; #100;
A = 8'h36; B = 8'hBC; #100;
A = 8'h36; B = 8'hBD; #100;
A = 8'h36; B = 8'hBE; #100;
A = 8'h36; B = 8'hBF; #100;
A = 8'h36; B = 8'hC0; #100;
A = 8'h36; B = 8'hC1; #100;
A = 8'h36; B = 8'hC2; #100;
A = 8'h36; B = 8'hC3; #100;
A = 8'h36; B = 8'hC4; #100;
A = 8'h36; B = 8'hC5; #100;
A = 8'h36; B = 8'hC6; #100;
A = 8'h36; B = 8'hC7; #100;
A = 8'h36; B = 8'hC8; #100;
A = 8'h36; B = 8'hC9; #100;
A = 8'h36; B = 8'hCA; #100;
A = 8'h36; B = 8'hCB; #100;
A = 8'h36; B = 8'hCC; #100;
A = 8'h36; B = 8'hCD; #100;
A = 8'h36; B = 8'hCE; #100;
A = 8'h36; B = 8'hCF; #100;
A = 8'h36; B = 8'hD0; #100;
A = 8'h36; B = 8'hD1; #100;
A = 8'h36; B = 8'hD2; #100;
A = 8'h36; B = 8'hD3; #100;
A = 8'h36; B = 8'hD4; #100;
A = 8'h36; B = 8'hD5; #100;
A = 8'h36; B = 8'hD6; #100;
A = 8'h36; B = 8'hD7; #100;
A = 8'h36; B = 8'hD8; #100;
A = 8'h36; B = 8'hD9; #100;
A = 8'h36; B = 8'hDA; #100;
A = 8'h36; B = 8'hDB; #100;
A = 8'h36; B = 8'hDC; #100;
A = 8'h36; B = 8'hDD; #100;
A = 8'h36; B = 8'hDE; #100;
A = 8'h36; B = 8'hDF; #100;
A = 8'h36; B = 8'hE0; #100;
A = 8'h36; B = 8'hE1; #100;
A = 8'h36; B = 8'hE2; #100;
A = 8'h36; B = 8'hE3; #100;
A = 8'h36; B = 8'hE4; #100;
A = 8'h36; B = 8'hE5; #100;
A = 8'h36; B = 8'hE6; #100;
A = 8'h36; B = 8'hE7; #100;
A = 8'h36; B = 8'hE8; #100;
A = 8'h36; B = 8'hE9; #100;
A = 8'h36; B = 8'hEA; #100;
A = 8'h36; B = 8'hEB; #100;
A = 8'h36; B = 8'hEC; #100;
A = 8'h36; B = 8'hED; #100;
A = 8'h36; B = 8'hEE; #100;
A = 8'h36; B = 8'hEF; #100;
A = 8'h36; B = 8'hF0; #100;
A = 8'h36; B = 8'hF1; #100;
A = 8'h36; B = 8'hF2; #100;
A = 8'h36; B = 8'hF3; #100;
A = 8'h36; B = 8'hF4; #100;
A = 8'h36; B = 8'hF5; #100;
A = 8'h36; B = 8'hF6; #100;
A = 8'h36; B = 8'hF7; #100;
A = 8'h36; B = 8'hF8; #100;
A = 8'h36; B = 8'hF9; #100;
A = 8'h36; B = 8'hFA; #100;
A = 8'h36; B = 8'hFB; #100;
A = 8'h36; B = 8'hFC; #100;
A = 8'h36; B = 8'hFD; #100;
A = 8'h36; B = 8'hFE; #100;
A = 8'h36; B = 8'hFF; #100;
A = 8'h37; B = 8'h0; #100;
A = 8'h37; B = 8'h1; #100;
A = 8'h37; B = 8'h2; #100;
A = 8'h37; B = 8'h3; #100;
A = 8'h37; B = 8'h4; #100;
A = 8'h37; B = 8'h5; #100;
A = 8'h37; B = 8'h6; #100;
A = 8'h37; B = 8'h7; #100;
A = 8'h37; B = 8'h8; #100;
A = 8'h37; B = 8'h9; #100;
A = 8'h37; B = 8'hA; #100;
A = 8'h37; B = 8'hB; #100;
A = 8'h37; B = 8'hC; #100;
A = 8'h37; B = 8'hD; #100;
A = 8'h37; B = 8'hE; #100;
A = 8'h37; B = 8'hF; #100;
A = 8'h37; B = 8'h10; #100;
A = 8'h37; B = 8'h11; #100;
A = 8'h37; B = 8'h12; #100;
A = 8'h37; B = 8'h13; #100;
A = 8'h37; B = 8'h14; #100;
A = 8'h37; B = 8'h15; #100;
A = 8'h37; B = 8'h16; #100;
A = 8'h37; B = 8'h17; #100;
A = 8'h37; B = 8'h18; #100;
A = 8'h37; B = 8'h19; #100;
A = 8'h37; B = 8'h1A; #100;
A = 8'h37; B = 8'h1B; #100;
A = 8'h37; B = 8'h1C; #100;
A = 8'h37; B = 8'h1D; #100;
A = 8'h37; B = 8'h1E; #100;
A = 8'h37; B = 8'h1F; #100;
A = 8'h37; B = 8'h20; #100;
A = 8'h37; B = 8'h21; #100;
A = 8'h37; B = 8'h22; #100;
A = 8'h37; B = 8'h23; #100;
A = 8'h37; B = 8'h24; #100;
A = 8'h37; B = 8'h25; #100;
A = 8'h37; B = 8'h26; #100;
A = 8'h37; B = 8'h27; #100;
A = 8'h37; B = 8'h28; #100;
A = 8'h37; B = 8'h29; #100;
A = 8'h37; B = 8'h2A; #100;
A = 8'h37; B = 8'h2B; #100;
A = 8'h37; B = 8'h2C; #100;
A = 8'h37; B = 8'h2D; #100;
A = 8'h37; B = 8'h2E; #100;
A = 8'h37; B = 8'h2F; #100;
A = 8'h37; B = 8'h30; #100;
A = 8'h37; B = 8'h31; #100;
A = 8'h37; B = 8'h32; #100;
A = 8'h37; B = 8'h33; #100;
A = 8'h37; B = 8'h34; #100;
A = 8'h37; B = 8'h35; #100;
A = 8'h37; B = 8'h36; #100;
A = 8'h37; B = 8'h37; #100;
A = 8'h37; B = 8'h38; #100;
A = 8'h37; B = 8'h39; #100;
A = 8'h37; B = 8'h3A; #100;
A = 8'h37; B = 8'h3B; #100;
A = 8'h37; B = 8'h3C; #100;
A = 8'h37; B = 8'h3D; #100;
A = 8'h37; B = 8'h3E; #100;
A = 8'h37; B = 8'h3F; #100;
A = 8'h37; B = 8'h40; #100;
A = 8'h37; B = 8'h41; #100;
A = 8'h37; B = 8'h42; #100;
A = 8'h37; B = 8'h43; #100;
A = 8'h37; B = 8'h44; #100;
A = 8'h37; B = 8'h45; #100;
A = 8'h37; B = 8'h46; #100;
A = 8'h37; B = 8'h47; #100;
A = 8'h37; B = 8'h48; #100;
A = 8'h37; B = 8'h49; #100;
A = 8'h37; B = 8'h4A; #100;
A = 8'h37; B = 8'h4B; #100;
A = 8'h37; B = 8'h4C; #100;
A = 8'h37; B = 8'h4D; #100;
A = 8'h37; B = 8'h4E; #100;
A = 8'h37; B = 8'h4F; #100;
A = 8'h37; B = 8'h50; #100;
A = 8'h37; B = 8'h51; #100;
A = 8'h37; B = 8'h52; #100;
A = 8'h37; B = 8'h53; #100;
A = 8'h37; B = 8'h54; #100;
A = 8'h37; B = 8'h55; #100;
A = 8'h37; B = 8'h56; #100;
A = 8'h37; B = 8'h57; #100;
A = 8'h37; B = 8'h58; #100;
A = 8'h37; B = 8'h59; #100;
A = 8'h37; B = 8'h5A; #100;
A = 8'h37; B = 8'h5B; #100;
A = 8'h37; B = 8'h5C; #100;
A = 8'h37; B = 8'h5D; #100;
A = 8'h37; B = 8'h5E; #100;
A = 8'h37; B = 8'h5F; #100;
A = 8'h37; B = 8'h60; #100;
A = 8'h37; B = 8'h61; #100;
A = 8'h37; B = 8'h62; #100;
A = 8'h37; B = 8'h63; #100;
A = 8'h37; B = 8'h64; #100;
A = 8'h37; B = 8'h65; #100;
A = 8'h37; B = 8'h66; #100;
A = 8'h37; B = 8'h67; #100;
A = 8'h37; B = 8'h68; #100;
A = 8'h37; B = 8'h69; #100;
A = 8'h37; B = 8'h6A; #100;
A = 8'h37; B = 8'h6B; #100;
A = 8'h37; B = 8'h6C; #100;
A = 8'h37; B = 8'h6D; #100;
A = 8'h37; B = 8'h6E; #100;
A = 8'h37; B = 8'h6F; #100;
A = 8'h37; B = 8'h70; #100;
A = 8'h37; B = 8'h71; #100;
A = 8'h37; B = 8'h72; #100;
A = 8'h37; B = 8'h73; #100;
A = 8'h37; B = 8'h74; #100;
A = 8'h37; B = 8'h75; #100;
A = 8'h37; B = 8'h76; #100;
A = 8'h37; B = 8'h77; #100;
A = 8'h37; B = 8'h78; #100;
A = 8'h37; B = 8'h79; #100;
A = 8'h37; B = 8'h7A; #100;
A = 8'h37; B = 8'h7B; #100;
A = 8'h37; B = 8'h7C; #100;
A = 8'h37; B = 8'h7D; #100;
A = 8'h37; B = 8'h7E; #100;
A = 8'h37; B = 8'h7F; #100;
A = 8'h37; B = 8'h80; #100;
A = 8'h37; B = 8'h81; #100;
A = 8'h37; B = 8'h82; #100;
A = 8'h37; B = 8'h83; #100;
A = 8'h37; B = 8'h84; #100;
A = 8'h37; B = 8'h85; #100;
A = 8'h37; B = 8'h86; #100;
A = 8'h37; B = 8'h87; #100;
A = 8'h37; B = 8'h88; #100;
A = 8'h37; B = 8'h89; #100;
A = 8'h37; B = 8'h8A; #100;
A = 8'h37; B = 8'h8B; #100;
A = 8'h37; B = 8'h8C; #100;
A = 8'h37; B = 8'h8D; #100;
A = 8'h37; B = 8'h8E; #100;
A = 8'h37; B = 8'h8F; #100;
A = 8'h37; B = 8'h90; #100;
A = 8'h37; B = 8'h91; #100;
A = 8'h37; B = 8'h92; #100;
A = 8'h37; B = 8'h93; #100;
A = 8'h37; B = 8'h94; #100;
A = 8'h37; B = 8'h95; #100;
A = 8'h37; B = 8'h96; #100;
A = 8'h37; B = 8'h97; #100;
A = 8'h37; B = 8'h98; #100;
A = 8'h37; B = 8'h99; #100;
A = 8'h37; B = 8'h9A; #100;
A = 8'h37; B = 8'h9B; #100;
A = 8'h37; B = 8'h9C; #100;
A = 8'h37; B = 8'h9D; #100;
A = 8'h37; B = 8'h9E; #100;
A = 8'h37; B = 8'h9F; #100;
A = 8'h37; B = 8'hA0; #100;
A = 8'h37; B = 8'hA1; #100;
A = 8'h37; B = 8'hA2; #100;
A = 8'h37; B = 8'hA3; #100;
A = 8'h37; B = 8'hA4; #100;
A = 8'h37; B = 8'hA5; #100;
A = 8'h37; B = 8'hA6; #100;
A = 8'h37; B = 8'hA7; #100;
A = 8'h37; B = 8'hA8; #100;
A = 8'h37; B = 8'hA9; #100;
A = 8'h37; B = 8'hAA; #100;
A = 8'h37; B = 8'hAB; #100;
A = 8'h37; B = 8'hAC; #100;
A = 8'h37; B = 8'hAD; #100;
A = 8'h37; B = 8'hAE; #100;
A = 8'h37; B = 8'hAF; #100;
A = 8'h37; B = 8'hB0; #100;
A = 8'h37; B = 8'hB1; #100;
A = 8'h37; B = 8'hB2; #100;
A = 8'h37; B = 8'hB3; #100;
A = 8'h37; B = 8'hB4; #100;
A = 8'h37; B = 8'hB5; #100;
A = 8'h37; B = 8'hB6; #100;
A = 8'h37; B = 8'hB7; #100;
A = 8'h37; B = 8'hB8; #100;
A = 8'h37; B = 8'hB9; #100;
A = 8'h37; B = 8'hBA; #100;
A = 8'h37; B = 8'hBB; #100;
A = 8'h37; B = 8'hBC; #100;
A = 8'h37; B = 8'hBD; #100;
A = 8'h37; B = 8'hBE; #100;
A = 8'h37; B = 8'hBF; #100;
A = 8'h37; B = 8'hC0; #100;
A = 8'h37; B = 8'hC1; #100;
A = 8'h37; B = 8'hC2; #100;
A = 8'h37; B = 8'hC3; #100;
A = 8'h37; B = 8'hC4; #100;
A = 8'h37; B = 8'hC5; #100;
A = 8'h37; B = 8'hC6; #100;
A = 8'h37; B = 8'hC7; #100;
A = 8'h37; B = 8'hC8; #100;
A = 8'h37; B = 8'hC9; #100;
A = 8'h37; B = 8'hCA; #100;
A = 8'h37; B = 8'hCB; #100;
A = 8'h37; B = 8'hCC; #100;
A = 8'h37; B = 8'hCD; #100;
A = 8'h37; B = 8'hCE; #100;
A = 8'h37; B = 8'hCF; #100;
A = 8'h37; B = 8'hD0; #100;
A = 8'h37; B = 8'hD1; #100;
A = 8'h37; B = 8'hD2; #100;
A = 8'h37; B = 8'hD3; #100;
A = 8'h37; B = 8'hD4; #100;
A = 8'h37; B = 8'hD5; #100;
A = 8'h37; B = 8'hD6; #100;
A = 8'h37; B = 8'hD7; #100;
A = 8'h37; B = 8'hD8; #100;
A = 8'h37; B = 8'hD9; #100;
A = 8'h37; B = 8'hDA; #100;
A = 8'h37; B = 8'hDB; #100;
A = 8'h37; B = 8'hDC; #100;
A = 8'h37; B = 8'hDD; #100;
A = 8'h37; B = 8'hDE; #100;
A = 8'h37; B = 8'hDF; #100;
A = 8'h37; B = 8'hE0; #100;
A = 8'h37; B = 8'hE1; #100;
A = 8'h37; B = 8'hE2; #100;
A = 8'h37; B = 8'hE3; #100;
A = 8'h37; B = 8'hE4; #100;
A = 8'h37; B = 8'hE5; #100;
A = 8'h37; B = 8'hE6; #100;
A = 8'h37; B = 8'hE7; #100;
A = 8'h37; B = 8'hE8; #100;
A = 8'h37; B = 8'hE9; #100;
A = 8'h37; B = 8'hEA; #100;
A = 8'h37; B = 8'hEB; #100;
A = 8'h37; B = 8'hEC; #100;
A = 8'h37; B = 8'hED; #100;
A = 8'h37; B = 8'hEE; #100;
A = 8'h37; B = 8'hEF; #100;
A = 8'h37; B = 8'hF0; #100;
A = 8'h37; B = 8'hF1; #100;
A = 8'h37; B = 8'hF2; #100;
A = 8'h37; B = 8'hF3; #100;
A = 8'h37; B = 8'hF4; #100;
A = 8'h37; B = 8'hF5; #100;
A = 8'h37; B = 8'hF6; #100;
A = 8'h37; B = 8'hF7; #100;
A = 8'h37; B = 8'hF8; #100;
A = 8'h37; B = 8'hF9; #100;
A = 8'h37; B = 8'hFA; #100;
A = 8'h37; B = 8'hFB; #100;
A = 8'h37; B = 8'hFC; #100;
A = 8'h37; B = 8'hFD; #100;
A = 8'h37; B = 8'hFE; #100;
A = 8'h37; B = 8'hFF; #100;
A = 8'h38; B = 8'h0; #100;
A = 8'h38; B = 8'h1; #100;
A = 8'h38; B = 8'h2; #100;
A = 8'h38; B = 8'h3; #100;
A = 8'h38; B = 8'h4; #100;
A = 8'h38; B = 8'h5; #100;
A = 8'h38; B = 8'h6; #100;
A = 8'h38; B = 8'h7; #100;
A = 8'h38; B = 8'h8; #100;
A = 8'h38; B = 8'h9; #100;
A = 8'h38; B = 8'hA; #100;
A = 8'h38; B = 8'hB; #100;
A = 8'h38; B = 8'hC; #100;
A = 8'h38; B = 8'hD; #100;
A = 8'h38; B = 8'hE; #100;
A = 8'h38; B = 8'hF; #100;
A = 8'h38; B = 8'h10; #100;
A = 8'h38; B = 8'h11; #100;
A = 8'h38; B = 8'h12; #100;
A = 8'h38; B = 8'h13; #100;
A = 8'h38; B = 8'h14; #100;
A = 8'h38; B = 8'h15; #100;
A = 8'h38; B = 8'h16; #100;
A = 8'h38; B = 8'h17; #100;
A = 8'h38; B = 8'h18; #100;
A = 8'h38; B = 8'h19; #100;
A = 8'h38; B = 8'h1A; #100;
A = 8'h38; B = 8'h1B; #100;
A = 8'h38; B = 8'h1C; #100;
A = 8'h38; B = 8'h1D; #100;
A = 8'h38; B = 8'h1E; #100;
A = 8'h38; B = 8'h1F; #100;
A = 8'h38; B = 8'h20; #100;
A = 8'h38; B = 8'h21; #100;
A = 8'h38; B = 8'h22; #100;
A = 8'h38; B = 8'h23; #100;
A = 8'h38; B = 8'h24; #100;
A = 8'h38; B = 8'h25; #100;
A = 8'h38; B = 8'h26; #100;
A = 8'h38; B = 8'h27; #100;
A = 8'h38; B = 8'h28; #100;
A = 8'h38; B = 8'h29; #100;
A = 8'h38; B = 8'h2A; #100;
A = 8'h38; B = 8'h2B; #100;
A = 8'h38; B = 8'h2C; #100;
A = 8'h38; B = 8'h2D; #100;
A = 8'h38; B = 8'h2E; #100;
A = 8'h38; B = 8'h2F; #100;
A = 8'h38; B = 8'h30; #100;
A = 8'h38; B = 8'h31; #100;
A = 8'h38; B = 8'h32; #100;
A = 8'h38; B = 8'h33; #100;
A = 8'h38; B = 8'h34; #100;
A = 8'h38; B = 8'h35; #100;
A = 8'h38; B = 8'h36; #100;
A = 8'h38; B = 8'h37; #100;
A = 8'h38; B = 8'h38; #100;
A = 8'h38; B = 8'h39; #100;
A = 8'h38; B = 8'h3A; #100;
A = 8'h38; B = 8'h3B; #100;
A = 8'h38; B = 8'h3C; #100;
A = 8'h38; B = 8'h3D; #100;
A = 8'h38; B = 8'h3E; #100;
A = 8'h38; B = 8'h3F; #100;
A = 8'h38; B = 8'h40; #100;
A = 8'h38; B = 8'h41; #100;
A = 8'h38; B = 8'h42; #100;
A = 8'h38; B = 8'h43; #100;
A = 8'h38; B = 8'h44; #100;
A = 8'h38; B = 8'h45; #100;
A = 8'h38; B = 8'h46; #100;
A = 8'h38; B = 8'h47; #100;
A = 8'h38; B = 8'h48; #100;
A = 8'h38; B = 8'h49; #100;
A = 8'h38; B = 8'h4A; #100;
A = 8'h38; B = 8'h4B; #100;
A = 8'h38; B = 8'h4C; #100;
A = 8'h38; B = 8'h4D; #100;
A = 8'h38; B = 8'h4E; #100;
A = 8'h38; B = 8'h4F; #100;
A = 8'h38; B = 8'h50; #100;
A = 8'h38; B = 8'h51; #100;
A = 8'h38; B = 8'h52; #100;
A = 8'h38; B = 8'h53; #100;
A = 8'h38; B = 8'h54; #100;
A = 8'h38; B = 8'h55; #100;
A = 8'h38; B = 8'h56; #100;
A = 8'h38; B = 8'h57; #100;
A = 8'h38; B = 8'h58; #100;
A = 8'h38; B = 8'h59; #100;
A = 8'h38; B = 8'h5A; #100;
A = 8'h38; B = 8'h5B; #100;
A = 8'h38; B = 8'h5C; #100;
A = 8'h38; B = 8'h5D; #100;
A = 8'h38; B = 8'h5E; #100;
A = 8'h38; B = 8'h5F; #100;
A = 8'h38; B = 8'h60; #100;
A = 8'h38; B = 8'h61; #100;
A = 8'h38; B = 8'h62; #100;
A = 8'h38; B = 8'h63; #100;
A = 8'h38; B = 8'h64; #100;
A = 8'h38; B = 8'h65; #100;
A = 8'h38; B = 8'h66; #100;
A = 8'h38; B = 8'h67; #100;
A = 8'h38; B = 8'h68; #100;
A = 8'h38; B = 8'h69; #100;
A = 8'h38; B = 8'h6A; #100;
A = 8'h38; B = 8'h6B; #100;
A = 8'h38; B = 8'h6C; #100;
A = 8'h38; B = 8'h6D; #100;
A = 8'h38; B = 8'h6E; #100;
A = 8'h38; B = 8'h6F; #100;
A = 8'h38; B = 8'h70; #100;
A = 8'h38; B = 8'h71; #100;
A = 8'h38; B = 8'h72; #100;
A = 8'h38; B = 8'h73; #100;
A = 8'h38; B = 8'h74; #100;
A = 8'h38; B = 8'h75; #100;
A = 8'h38; B = 8'h76; #100;
A = 8'h38; B = 8'h77; #100;
A = 8'h38; B = 8'h78; #100;
A = 8'h38; B = 8'h79; #100;
A = 8'h38; B = 8'h7A; #100;
A = 8'h38; B = 8'h7B; #100;
A = 8'h38; B = 8'h7C; #100;
A = 8'h38; B = 8'h7D; #100;
A = 8'h38; B = 8'h7E; #100;
A = 8'h38; B = 8'h7F; #100;
A = 8'h38; B = 8'h80; #100;
A = 8'h38; B = 8'h81; #100;
A = 8'h38; B = 8'h82; #100;
A = 8'h38; B = 8'h83; #100;
A = 8'h38; B = 8'h84; #100;
A = 8'h38; B = 8'h85; #100;
A = 8'h38; B = 8'h86; #100;
A = 8'h38; B = 8'h87; #100;
A = 8'h38; B = 8'h88; #100;
A = 8'h38; B = 8'h89; #100;
A = 8'h38; B = 8'h8A; #100;
A = 8'h38; B = 8'h8B; #100;
A = 8'h38; B = 8'h8C; #100;
A = 8'h38; B = 8'h8D; #100;
A = 8'h38; B = 8'h8E; #100;
A = 8'h38; B = 8'h8F; #100;
A = 8'h38; B = 8'h90; #100;
A = 8'h38; B = 8'h91; #100;
A = 8'h38; B = 8'h92; #100;
A = 8'h38; B = 8'h93; #100;
A = 8'h38; B = 8'h94; #100;
A = 8'h38; B = 8'h95; #100;
A = 8'h38; B = 8'h96; #100;
A = 8'h38; B = 8'h97; #100;
A = 8'h38; B = 8'h98; #100;
A = 8'h38; B = 8'h99; #100;
A = 8'h38; B = 8'h9A; #100;
A = 8'h38; B = 8'h9B; #100;
A = 8'h38; B = 8'h9C; #100;
A = 8'h38; B = 8'h9D; #100;
A = 8'h38; B = 8'h9E; #100;
A = 8'h38; B = 8'h9F; #100;
A = 8'h38; B = 8'hA0; #100;
A = 8'h38; B = 8'hA1; #100;
A = 8'h38; B = 8'hA2; #100;
A = 8'h38; B = 8'hA3; #100;
A = 8'h38; B = 8'hA4; #100;
A = 8'h38; B = 8'hA5; #100;
A = 8'h38; B = 8'hA6; #100;
A = 8'h38; B = 8'hA7; #100;
A = 8'h38; B = 8'hA8; #100;
A = 8'h38; B = 8'hA9; #100;
A = 8'h38; B = 8'hAA; #100;
A = 8'h38; B = 8'hAB; #100;
A = 8'h38; B = 8'hAC; #100;
A = 8'h38; B = 8'hAD; #100;
A = 8'h38; B = 8'hAE; #100;
A = 8'h38; B = 8'hAF; #100;
A = 8'h38; B = 8'hB0; #100;
A = 8'h38; B = 8'hB1; #100;
A = 8'h38; B = 8'hB2; #100;
A = 8'h38; B = 8'hB3; #100;
A = 8'h38; B = 8'hB4; #100;
A = 8'h38; B = 8'hB5; #100;
A = 8'h38; B = 8'hB6; #100;
A = 8'h38; B = 8'hB7; #100;
A = 8'h38; B = 8'hB8; #100;
A = 8'h38; B = 8'hB9; #100;
A = 8'h38; B = 8'hBA; #100;
A = 8'h38; B = 8'hBB; #100;
A = 8'h38; B = 8'hBC; #100;
A = 8'h38; B = 8'hBD; #100;
A = 8'h38; B = 8'hBE; #100;
A = 8'h38; B = 8'hBF; #100;
A = 8'h38; B = 8'hC0; #100;
A = 8'h38; B = 8'hC1; #100;
A = 8'h38; B = 8'hC2; #100;
A = 8'h38; B = 8'hC3; #100;
A = 8'h38; B = 8'hC4; #100;
A = 8'h38; B = 8'hC5; #100;
A = 8'h38; B = 8'hC6; #100;
A = 8'h38; B = 8'hC7; #100;
A = 8'h38; B = 8'hC8; #100;
A = 8'h38; B = 8'hC9; #100;
A = 8'h38; B = 8'hCA; #100;
A = 8'h38; B = 8'hCB; #100;
A = 8'h38; B = 8'hCC; #100;
A = 8'h38; B = 8'hCD; #100;
A = 8'h38; B = 8'hCE; #100;
A = 8'h38; B = 8'hCF; #100;
A = 8'h38; B = 8'hD0; #100;
A = 8'h38; B = 8'hD1; #100;
A = 8'h38; B = 8'hD2; #100;
A = 8'h38; B = 8'hD3; #100;
A = 8'h38; B = 8'hD4; #100;
A = 8'h38; B = 8'hD5; #100;
A = 8'h38; B = 8'hD6; #100;
A = 8'h38; B = 8'hD7; #100;
A = 8'h38; B = 8'hD8; #100;
A = 8'h38; B = 8'hD9; #100;
A = 8'h38; B = 8'hDA; #100;
A = 8'h38; B = 8'hDB; #100;
A = 8'h38; B = 8'hDC; #100;
A = 8'h38; B = 8'hDD; #100;
A = 8'h38; B = 8'hDE; #100;
A = 8'h38; B = 8'hDF; #100;
A = 8'h38; B = 8'hE0; #100;
A = 8'h38; B = 8'hE1; #100;
A = 8'h38; B = 8'hE2; #100;
A = 8'h38; B = 8'hE3; #100;
A = 8'h38; B = 8'hE4; #100;
A = 8'h38; B = 8'hE5; #100;
A = 8'h38; B = 8'hE6; #100;
A = 8'h38; B = 8'hE7; #100;
A = 8'h38; B = 8'hE8; #100;
A = 8'h38; B = 8'hE9; #100;
A = 8'h38; B = 8'hEA; #100;
A = 8'h38; B = 8'hEB; #100;
A = 8'h38; B = 8'hEC; #100;
A = 8'h38; B = 8'hED; #100;
A = 8'h38; B = 8'hEE; #100;
A = 8'h38; B = 8'hEF; #100;
A = 8'h38; B = 8'hF0; #100;
A = 8'h38; B = 8'hF1; #100;
A = 8'h38; B = 8'hF2; #100;
A = 8'h38; B = 8'hF3; #100;
A = 8'h38; B = 8'hF4; #100;
A = 8'h38; B = 8'hF5; #100;
A = 8'h38; B = 8'hF6; #100;
A = 8'h38; B = 8'hF7; #100;
A = 8'h38; B = 8'hF8; #100;
A = 8'h38; B = 8'hF9; #100;
A = 8'h38; B = 8'hFA; #100;
A = 8'h38; B = 8'hFB; #100;
A = 8'h38; B = 8'hFC; #100;
A = 8'h38; B = 8'hFD; #100;
A = 8'h38; B = 8'hFE; #100;
A = 8'h38; B = 8'hFF; #100;
A = 8'h39; B = 8'h0; #100;
A = 8'h39; B = 8'h1; #100;
A = 8'h39; B = 8'h2; #100;
A = 8'h39; B = 8'h3; #100;
A = 8'h39; B = 8'h4; #100;
A = 8'h39; B = 8'h5; #100;
A = 8'h39; B = 8'h6; #100;
A = 8'h39; B = 8'h7; #100;
A = 8'h39; B = 8'h8; #100;
A = 8'h39; B = 8'h9; #100;
A = 8'h39; B = 8'hA; #100;
A = 8'h39; B = 8'hB; #100;
A = 8'h39; B = 8'hC; #100;
A = 8'h39; B = 8'hD; #100;
A = 8'h39; B = 8'hE; #100;
A = 8'h39; B = 8'hF; #100;
A = 8'h39; B = 8'h10; #100;
A = 8'h39; B = 8'h11; #100;
A = 8'h39; B = 8'h12; #100;
A = 8'h39; B = 8'h13; #100;
A = 8'h39; B = 8'h14; #100;
A = 8'h39; B = 8'h15; #100;
A = 8'h39; B = 8'h16; #100;
A = 8'h39; B = 8'h17; #100;
A = 8'h39; B = 8'h18; #100;
A = 8'h39; B = 8'h19; #100;
A = 8'h39; B = 8'h1A; #100;
A = 8'h39; B = 8'h1B; #100;
A = 8'h39; B = 8'h1C; #100;
A = 8'h39; B = 8'h1D; #100;
A = 8'h39; B = 8'h1E; #100;
A = 8'h39; B = 8'h1F; #100;
A = 8'h39; B = 8'h20; #100;
A = 8'h39; B = 8'h21; #100;
A = 8'h39; B = 8'h22; #100;
A = 8'h39; B = 8'h23; #100;
A = 8'h39; B = 8'h24; #100;
A = 8'h39; B = 8'h25; #100;
A = 8'h39; B = 8'h26; #100;
A = 8'h39; B = 8'h27; #100;
A = 8'h39; B = 8'h28; #100;
A = 8'h39; B = 8'h29; #100;
A = 8'h39; B = 8'h2A; #100;
A = 8'h39; B = 8'h2B; #100;
A = 8'h39; B = 8'h2C; #100;
A = 8'h39; B = 8'h2D; #100;
A = 8'h39; B = 8'h2E; #100;
A = 8'h39; B = 8'h2F; #100;
A = 8'h39; B = 8'h30; #100;
A = 8'h39; B = 8'h31; #100;
A = 8'h39; B = 8'h32; #100;
A = 8'h39; B = 8'h33; #100;
A = 8'h39; B = 8'h34; #100;
A = 8'h39; B = 8'h35; #100;
A = 8'h39; B = 8'h36; #100;
A = 8'h39; B = 8'h37; #100;
A = 8'h39; B = 8'h38; #100;
A = 8'h39; B = 8'h39; #100;
A = 8'h39; B = 8'h3A; #100;
A = 8'h39; B = 8'h3B; #100;
A = 8'h39; B = 8'h3C; #100;
A = 8'h39; B = 8'h3D; #100;
A = 8'h39; B = 8'h3E; #100;
A = 8'h39; B = 8'h3F; #100;
A = 8'h39; B = 8'h40; #100;
A = 8'h39; B = 8'h41; #100;
A = 8'h39; B = 8'h42; #100;
A = 8'h39; B = 8'h43; #100;
A = 8'h39; B = 8'h44; #100;
A = 8'h39; B = 8'h45; #100;
A = 8'h39; B = 8'h46; #100;
A = 8'h39; B = 8'h47; #100;
A = 8'h39; B = 8'h48; #100;
A = 8'h39; B = 8'h49; #100;
A = 8'h39; B = 8'h4A; #100;
A = 8'h39; B = 8'h4B; #100;
A = 8'h39; B = 8'h4C; #100;
A = 8'h39; B = 8'h4D; #100;
A = 8'h39; B = 8'h4E; #100;
A = 8'h39; B = 8'h4F; #100;
A = 8'h39; B = 8'h50; #100;
A = 8'h39; B = 8'h51; #100;
A = 8'h39; B = 8'h52; #100;
A = 8'h39; B = 8'h53; #100;
A = 8'h39; B = 8'h54; #100;
A = 8'h39; B = 8'h55; #100;
A = 8'h39; B = 8'h56; #100;
A = 8'h39; B = 8'h57; #100;
A = 8'h39; B = 8'h58; #100;
A = 8'h39; B = 8'h59; #100;
A = 8'h39; B = 8'h5A; #100;
A = 8'h39; B = 8'h5B; #100;
A = 8'h39; B = 8'h5C; #100;
A = 8'h39; B = 8'h5D; #100;
A = 8'h39; B = 8'h5E; #100;
A = 8'h39; B = 8'h5F; #100;
A = 8'h39; B = 8'h60; #100;
A = 8'h39; B = 8'h61; #100;
A = 8'h39; B = 8'h62; #100;
A = 8'h39; B = 8'h63; #100;
A = 8'h39; B = 8'h64; #100;
A = 8'h39; B = 8'h65; #100;
A = 8'h39; B = 8'h66; #100;
A = 8'h39; B = 8'h67; #100;
A = 8'h39; B = 8'h68; #100;
A = 8'h39; B = 8'h69; #100;
A = 8'h39; B = 8'h6A; #100;
A = 8'h39; B = 8'h6B; #100;
A = 8'h39; B = 8'h6C; #100;
A = 8'h39; B = 8'h6D; #100;
A = 8'h39; B = 8'h6E; #100;
A = 8'h39; B = 8'h6F; #100;
A = 8'h39; B = 8'h70; #100;
A = 8'h39; B = 8'h71; #100;
A = 8'h39; B = 8'h72; #100;
A = 8'h39; B = 8'h73; #100;
A = 8'h39; B = 8'h74; #100;
A = 8'h39; B = 8'h75; #100;
A = 8'h39; B = 8'h76; #100;
A = 8'h39; B = 8'h77; #100;
A = 8'h39; B = 8'h78; #100;
A = 8'h39; B = 8'h79; #100;
A = 8'h39; B = 8'h7A; #100;
A = 8'h39; B = 8'h7B; #100;
A = 8'h39; B = 8'h7C; #100;
A = 8'h39; B = 8'h7D; #100;
A = 8'h39; B = 8'h7E; #100;
A = 8'h39; B = 8'h7F; #100;
A = 8'h39; B = 8'h80; #100;
A = 8'h39; B = 8'h81; #100;
A = 8'h39; B = 8'h82; #100;
A = 8'h39; B = 8'h83; #100;
A = 8'h39; B = 8'h84; #100;
A = 8'h39; B = 8'h85; #100;
A = 8'h39; B = 8'h86; #100;
A = 8'h39; B = 8'h87; #100;
A = 8'h39; B = 8'h88; #100;
A = 8'h39; B = 8'h89; #100;
A = 8'h39; B = 8'h8A; #100;
A = 8'h39; B = 8'h8B; #100;
A = 8'h39; B = 8'h8C; #100;
A = 8'h39; B = 8'h8D; #100;
A = 8'h39; B = 8'h8E; #100;
A = 8'h39; B = 8'h8F; #100;
A = 8'h39; B = 8'h90; #100;
A = 8'h39; B = 8'h91; #100;
A = 8'h39; B = 8'h92; #100;
A = 8'h39; B = 8'h93; #100;
A = 8'h39; B = 8'h94; #100;
A = 8'h39; B = 8'h95; #100;
A = 8'h39; B = 8'h96; #100;
A = 8'h39; B = 8'h97; #100;
A = 8'h39; B = 8'h98; #100;
A = 8'h39; B = 8'h99; #100;
A = 8'h39; B = 8'h9A; #100;
A = 8'h39; B = 8'h9B; #100;
A = 8'h39; B = 8'h9C; #100;
A = 8'h39; B = 8'h9D; #100;
A = 8'h39; B = 8'h9E; #100;
A = 8'h39; B = 8'h9F; #100;
A = 8'h39; B = 8'hA0; #100;
A = 8'h39; B = 8'hA1; #100;
A = 8'h39; B = 8'hA2; #100;
A = 8'h39; B = 8'hA3; #100;
A = 8'h39; B = 8'hA4; #100;
A = 8'h39; B = 8'hA5; #100;
A = 8'h39; B = 8'hA6; #100;
A = 8'h39; B = 8'hA7; #100;
A = 8'h39; B = 8'hA8; #100;
A = 8'h39; B = 8'hA9; #100;
A = 8'h39; B = 8'hAA; #100;
A = 8'h39; B = 8'hAB; #100;
A = 8'h39; B = 8'hAC; #100;
A = 8'h39; B = 8'hAD; #100;
A = 8'h39; B = 8'hAE; #100;
A = 8'h39; B = 8'hAF; #100;
A = 8'h39; B = 8'hB0; #100;
A = 8'h39; B = 8'hB1; #100;
A = 8'h39; B = 8'hB2; #100;
A = 8'h39; B = 8'hB3; #100;
A = 8'h39; B = 8'hB4; #100;
A = 8'h39; B = 8'hB5; #100;
A = 8'h39; B = 8'hB6; #100;
A = 8'h39; B = 8'hB7; #100;
A = 8'h39; B = 8'hB8; #100;
A = 8'h39; B = 8'hB9; #100;
A = 8'h39; B = 8'hBA; #100;
A = 8'h39; B = 8'hBB; #100;
A = 8'h39; B = 8'hBC; #100;
A = 8'h39; B = 8'hBD; #100;
A = 8'h39; B = 8'hBE; #100;
A = 8'h39; B = 8'hBF; #100;
A = 8'h39; B = 8'hC0; #100;
A = 8'h39; B = 8'hC1; #100;
A = 8'h39; B = 8'hC2; #100;
A = 8'h39; B = 8'hC3; #100;
A = 8'h39; B = 8'hC4; #100;
A = 8'h39; B = 8'hC5; #100;
A = 8'h39; B = 8'hC6; #100;
A = 8'h39; B = 8'hC7; #100;
A = 8'h39; B = 8'hC8; #100;
A = 8'h39; B = 8'hC9; #100;
A = 8'h39; B = 8'hCA; #100;
A = 8'h39; B = 8'hCB; #100;
A = 8'h39; B = 8'hCC; #100;
A = 8'h39; B = 8'hCD; #100;
A = 8'h39; B = 8'hCE; #100;
A = 8'h39; B = 8'hCF; #100;
A = 8'h39; B = 8'hD0; #100;
A = 8'h39; B = 8'hD1; #100;
A = 8'h39; B = 8'hD2; #100;
A = 8'h39; B = 8'hD3; #100;
A = 8'h39; B = 8'hD4; #100;
A = 8'h39; B = 8'hD5; #100;
A = 8'h39; B = 8'hD6; #100;
A = 8'h39; B = 8'hD7; #100;
A = 8'h39; B = 8'hD8; #100;
A = 8'h39; B = 8'hD9; #100;
A = 8'h39; B = 8'hDA; #100;
A = 8'h39; B = 8'hDB; #100;
A = 8'h39; B = 8'hDC; #100;
A = 8'h39; B = 8'hDD; #100;
A = 8'h39; B = 8'hDE; #100;
A = 8'h39; B = 8'hDF; #100;
A = 8'h39; B = 8'hE0; #100;
A = 8'h39; B = 8'hE1; #100;
A = 8'h39; B = 8'hE2; #100;
A = 8'h39; B = 8'hE3; #100;
A = 8'h39; B = 8'hE4; #100;
A = 8'h39; B = 8'hE5; #100;
A = 8'h39; B = 8'hE6; #100;
A = 8'h39; B = 8'hE7; #100;
A = 8'h39; B = 8'hE8; #100;
A = 8'h39; B = 8'hE9; #100;
A = 8'h39; B = 8'hEA; #100;
A = 8'h39; B = 8'hEB; #100;
A = 8'h39; B = 8'hEC; #100;
A = 8'h39; B = 8'hED; #100;
A = 8'h39; B = 8'hEE; #100;
A = 8'h39; B = 8'hEF; #100;
A = 8'h39; B = 8'hF0; #100;
A = 8'h39; B = 8'hF1; #100;
A = 8'h39; B = 8'hF2; #100;
A = 8'h39; B = 8'hF3; #100;
A = 8'h39; B = 8'hF4; #100;
A = 8'h39; B = 8'hF5; #100;
A = 8'h39; B = 8'hF6; #100;
A = 8'h39; B = 8'hF7; #100;
A = 8'h39; B = 8'hF8; #100;
A = 8'h39; B = 8'hF9; #100;
A = 8'h39; B = 8'hFA; #100;
A = 8'h39; B = 8'hFB; #100;
A = 8'h39; B = 8'hFC; #100;
A = 8'h39; B = 8'hFD; #100;
A = 8'h39; B = 8'hFE; #100;
A = 8'h39; B = 8'hFF; #100;
A = 8'h3A; B = 8'h0; #100;
A = 8'h3A; B = 8'h1; #100;
A = 8'h3A; B = 8'h2; #100;
A = 8'h3A; B = 8'h3; #100;
A = 8'h3A; B = 8'h4; #100;
A = 8'h3A; B = 8'h5; #100;
A = 8'h3A; B = 8'h6; #100;
A = 8'h3A; B = 8'h7; #100;
A = 8'h3A; B = 8'h8; #100;
A = 8'h3A; B = 8'h9; #100;
A = 8'h3A; B = 8'hA; #100;
A = 8'h3A; B = 8'hB; #100;
A = 8'h3A; B = 8'hC; #100;
A = 8'h3A; B = 8'hD; #100;
A = 8'h3A; B = 8'hE; #100;
A = 8'h3A; B = 8'hF; #100;
A = 8'h3A; B = 8'h10; #100;
A = 8'h3A; B = 8'h11; #100;
A = 8'h3A; B = 8'h12; #100;
A = 8'h3A; B = 8'h13; #100;
A = 8'h3A; B = 8'h14; #100;
A = 8'h3A; B = 8'h15; #100;
A = 8'h3A; B = 8'h16; #100;
A = 8'h3A; B = 8'h17; #100;
A = 8'h3A; B = 8'h18; #100;
A = 8'h3A; B = 8'h19; #100;
A = 8'h3A; B = 8'h1A; #100;
A = 8'h3A; B = 8'h1B; #100;
A = 8'h3A; B = 8'h1C; #100;
A = 8'h3A; B = 8'h1D; #100;
A = 8'h3A; B = 8'h1E; #100;
A = 8'h3A; B = 8'h1F; #100;
A = 8'h3A; B = 8'h20; #100;
A = 8'h3A; B = 8'h21; #100;
A = 8'h3A; B = 8'h22; #100;
A = 8'h3A; B = 8'h23; #100;
A = 8'h3A; B = 8'h24; #100;
A = 8'h3A; B = 8'h25; #100;
A = 8'h3A; B = 8'h26; #100;
A = 8'h3A; B = 8'h27; #100;
A = 8'h3A; B = 8'h28; #100;
A = 8'h3A; B = 8'h29; #100;
A = 8'h3A; B = 8'h2A; #100;
A = 8'h3A; B = 8'h2B; #100;
A = 8'h3A; B = 8'h2C; #100;
A = 8'h3A; B = 8'h2D; #100;
A = 8'h3A; B = 8'h2E; #100;
A = 8'h3A; B = 8'h2F; #100;
A = 8'h3A; B = 8'h30; #100;
A = 8'h3A; B = 8'h31; #100;
A = 8'h3A; B = 8'h32; #100;
A = 8'h3A; B = 8'h33; #100;
A = 8'h3A; B = 8'h34; #100;
A = 8'h3A; B = 8'h35; #100;
A = 8'h3A; B = 8'h36; #100;
A = 8'h3A; B = 8'h37; #100;
A = 8'h3A; B = 8'h38; #100;
A = 8'h3A; B = 8'h39; #100;
A = 8'h3A; B = 8'h3A; #100;
A = 8'h3A; B = 8'h3B; #100;
A = 8'h3A; B = 8'h3C; #100;
A = 8'h3A; B = 8'h3D; #100;
A = 8'h3A; B = 8'h3E; #100;
A = 8'h3A; B = 8'h3F; #100;
A = 8'h3A; B = 8'h40; #100;
A = 8'h3A; B = 8'h41; #100;
A = 8'h3A; B = 8'h42; #100;
A = 8'h3A; B = 8'h43; #100;
A = 8'h3A; B = 8'h44; #100;
A = 8'h3A; B = 8'h45; #100;
A = 8'h3A; B = 8'h46; #100;
A = 8'h3A; B = 8'h47; #100;
A = 8'h3A; B = 8'h48; #100;
A = 8'h3A; B = 8'h49; #100;
A = 8'h3A; B = 8'h4A; #100;
A = 8'h3A; B = 8'h4B; #100;
A = 8'h3A; B = 8'h4C; #100;
A = 8'h3A; B = 8'h4D; #100;
A = 8'h3A; B = 8'h4E; #100;
A = 8'h3A; B = 8'h4F; #100;
A = 8'h3A; B = 8'h50; #100;
A = 8'h3A; B = 8'h51; #100;
A = 8'h3A; B = 8'h52; #100;
A = 8'h3A; B = 8'h53; #100;
A = 8'h3A; B = 8'h54; #100;
A = 8'h3A; B = 8'h55; #100;
A = 8'h3A; B = 8'h56; #100;
A = 8'h3A; B = 8'h57; #100;
A = 8'h3A; B = 8'h58; #100;
A = 8'h3A; B = 8'h59; #100;
A = 8'h3A; B = 8'h5A; #100;
A = 8'h3A; B = 8'h5B; #100;
A = 8'h3A; B = 8'h5C; #100;
A = 8'h3A; B = 8'h5D; #100;
A = 8'h3A; B = 8'h5E; #100;
A = 8'h3A; B = 8'h5F; #100;
A = 8'h3A; B = 8'h60; #100;
A = 8'h3A; B = 8'h61; #100;
A = 8'h3A; B = 8'h62; #100;
A = 8'h3A; B = 8'h63; #100;
A = 8'h3A; B = 8'h64; #100;
A = 8'h3A; B = 8'h65; #100;
A = 8'h3A; B = 8'h66; #100;
A = 8'h3A; B = 8'h67; #100;
A = 8'h3A; B = 8'h68; #100;
A = 8'h3A; B = 8'h69; #100;
A = 8'h3A; B = 8'h6A; #100;
A = 8'h3A; B = 8'h6B; #100;
A = 8'h3A; B = 8'h6C; #100;
A = 8'h3A; B = 8'h6D; #100;
A = 8'h3A; B = 8'h6E; #100;
A = 8'h3A; B = 8'h6F; #100;
A = 8'h3A; B = 8'h70; #100;
A = 8'h3A; B = 8'h71; #100;
A = 8'h3A; B = 8'h72; #100;
A = 8'h3A; B = 8'h73; #100;
A = 8'h3A; B = 8'h74; #100;
A = 8'h3A; B = 8'h75; #100;
A = 8'h3A; B = 8'h76; #100;
A = 8'h3A; B = 8'h77; #100;
A = 8'h3A; B = 8'h78; #100;
A = 8'h3A; B = 8'h79; #100;
A = 8'h3A; B = 8'h7A; #100;
A = 8'h3A; B = 8'h7B; #100;
A = 8'h3A; B = 8'h7C; #100;
A = 8'h3A; B = 8'h7D; #100;
A = 8'h3A; B = 8'h7E; #100;
A = 8'h3A; B = 8'h7F; #100;
A = 8'h3A; B = 8'h80; #100;
A = 8'h3A; B = 8'h81; #100;
A = 8'h3A; B = 8'h82; #100;
A = 8'h3A; B = 8'h83; #100;
A = 8'h3A; B = 8'h84; #100;
A = 8'h3A; B = 8'h85; #100;
A = 8'h3A; B = 8'h86; #100;
A = 8'h3A; B = 8'h87; #100;
A = 8'h3A; B = 8'h88; #100;
A = 8'h3A; B = 8'h89; #100;
A = 8'h3A; B = 8'h8A; #100;
A = 8'h3A; B = 8'h8B; #100;
A = 8'h3A; B = 8'h8C; #100;
A = 8'h3A; B = 8'h8D; #100;
A = 8'h3A; B = 8'h8E; #100;
A = 8'h3A; B = 8'h8F; #100;
A = 8'h3A; B = 8'h90; #100;
A = 8'h3A; B = 8'h91; #100;
A = 8'h3A; B = 8'h92; #100;
A = 8'h3A; B = 8'h93; #100;
A = 8'h3A; B = 8'h94; #100;
A = 8'h3A; B = 8'h95; #100;
A = 8'h3A; B = 8'h96; #100;
A = 8'h3A; B = 8'h97; #100;
A = 8'h3A; B = 8'h98; #100;
A = 8'h3A; B = 8'h99; #100;
A = 8'h3A; B = 8'h9A; #100;
A = 8'h3A; B = 8'h9B; #100;
A = 8'h3A; B = 8'h9C; #100;
A = 8'h3A; B = 8'h9D; #100;
A = 8'h3A; B = 8'h9E; #100;
A = 8'h3A; B = 8'h9F; #100;
A = 8'h3A; B = 8'hA0; #100;
A = 8'h3A; B = 8'hA1; #100;
A = 8'h3A; B = 8'hA2; #100;
A = 8'h3A; B = 8'hA3; #100;
A = 8'h3A; B = 8'hA4; #100;
A = 8'h3A; B = 8'hA5; #100;
A = 8'h3A; B = 8'hA6; #100;
A = 8'h3A; B = 8'hA7; #100;
A = 8'h3A; B = 8'hA8; #100;
A = 8'h3A; B = 8'hA9; #100;
A = 8'h3A; B = 8'hAA; #100;
A = 8'h3A; B = 8'hAB; #100;
A = 8'h3A; B = 8'hAC; #100;
A = 8'h3A; B = 8'hAD; #100;
A = 8'h3A; B = 8'hAE; #100;
A = 8'h3A; B = 8'hAF; #100;
A = 8'h3A; B = 8'hB0; #100;
A = 8'h3A; B = 8'hB1; #100;
A = 8'h3A; B = 8'hB2; #100;
A = 8'h3A; B = 8'hB3; #100;
A = 8'h3A; B = 8'hB4; #100;
A = 8'h3A; B = 8'hB5; #100;
A = 8'h3A; B = 8'hB6; #100;
A = 8'h3A; B = 8'hB7; #100;
A = 8'h3A; B = 8'hB8; #100;
A = 8'h3A; B = 8'hB9; #100;
A = 8'h3A; B = 8'hBA; #100;
A = 8'h3A; B = 8'hBB; #100;
A = 8'h3A; B = 8'hBC; #100;
A = 8'h3A; B = 8'hBD; #100;
A = 8'h3A; B = 8'hBE; #100;
A = 8'h3A; B = 8'hBF; #100;
A = 8'h3A; B = 8'hC0; #100;
A = 8'h3A; B = 8'hC1; #100;
A = 8'h3A; B = 8'hC2; #100;
A = 8'h3A; B = 8'hC3; #100;
A = 8'h3A; B = 8'hC4; #100;
A = 8'h3A; B = 8'hC5; #100;
A = 8'h3A; B = 8'hC6; #100;
A = 8'h3A; B = 8'hC7; #100;
A = 8'h3A; B = 8'hC8; #100;
A = 8'h3A; B = 8'hC9; #100;
A = 8'h3A; B = 8'hCA; #100;
A = 8'h3A; B = 8'hCB; #100;
A = 8'h3A; B = 8'hCC; #100;
A = 8'h3A; B = 8'hCD; #100;
A = 8'h3A; B = 8'hCE; #100;
A = 8'h3A; B = 8'hCF; #100;
A = 8'h3A; B = 8'hD0; #100;
A = 8'h3A; B = 8'hD1; #100;
A = 8'h3A; B = 8'hD2; #100;
A = 8'h3A; B = 8'hD3; #100;
A = 8'h3A; B = 8'hD4; #100;
A = 8'h3A; B = 8'hD5; #100;
A = 8'h3A; B = 8'hD6; #100;
A = 8'h3A; B = 8'hD7; #100;
A = 8'h3A; B = 8'hD8; #100;
A = 8'h3A; B = 8'hD9; #100;
A = 8'h3A; B = 8'hDA; #100;
A = 8'h3A; B = 8'hDB; #100;
A = 8'h3A; B = 8'hDC; #100;
A = 8'h3A; B = 8'hDD; #100;
A = 8'h3A; B = 8'hDE; #100;
A = 8'h3A; B = 8'hDF; #100;
A = 8'h3A; B = 8'hE0; #100;
A = 8'h3A; B = 8'hE1; #100;
A = 8'h3A; B = 8'hE2; #100;
A = 8'h3A; B = 8'hE3; #100;
A = 8'h3A; B = 8'hE4; #100;
A = 8'h3A; B = 8'hE5; #100;
A = 8'h3A; B = 8'hE6; #100;
A = 8'h3A; B = 8'hE7; #100;
A = 8'h3A; B = 8'hE8; #100;
A = 8'h3A; B = 8'hE9; #100;
A = 8'h3A; B = 8'hEA; #100;
A = 8'h3A; B = 8'hEB; #100;
A = 8'h3A; B = 8'hEC; #100;
A = 8'h3A; B = 8'hED; #100;
A = 8'h3A; B = 8'hEE; #100;
A = 8'h3A; B = 8'hEF; #100;
A = 8'h3A; B = 8'hF0; #100;
A = 8'h3A; B = 8'hF1; #100;
A = 8'h3A; B = 8'hF2; #100;
A = 8'h3A; B = 8'hF3; #100;
A = 8'h3A; B = 8'hF4; #100;
A = 8'h3A; B = 8'hF5; #100;
A = 8'h3A; B = 8'hF6; #100;
A = 8'h3A; B = 8'hF7; #100;
A = 8'h3A; B = 8'hF8; #100;
A = 8'h3A; B = 8'hF9; #100;
A = 8'h3A; B = 8'hFA; #100;
A = 8'h3A; B = 8'hFB; #100;
A = 8'h3A; B = 8'hFC; #100;
A = 8'h3A; B = 8'hFD; #100;
A = 8'h3A; B = 8'hFE; #100;
A = 8'h3A; B = 8'hFF; #100;
A = 8'h3B; B = 8'h0; #100;
A = 8'h3B; B = 8'h1; #100;
A = 8'h3B; B = 8'h2; #100;
A = 8'h3B; B = 8'h3; #100;
A = 8'h3B; B = 8'h4; #100;
A = 8'h3B; B = 8'h5; #100;
A = 8'h3B; B = 8'h6; #100;
A = 8'h3B; B = 8'h7; #100;
A = 8'h3B; B = 8'h8; #100;
A = 8'h3B; B = 8'h9; #100;
A = 8'h3B; B = 8'hA; #100;
A = 8'h3B; B = 8'hB; #100;
A = 8'h3B; B = 8'hC; #100;
A = 8'h3B; B = 8'hD; #100;
A = 8'h3B; B = 8'hE; #100;
A = 8'h3B; B = 8'hF; #100;
A = 8'h3B; B = 8'h10; #100;
A = 8'h3B; B = 8'h11; #100;
A = 8'h3B; B = 8'h12; #100;
A = 8'h3B; B = 8'h13; #100;
A = 8'h3B; B = 8'h14; #100;
A = 8'h3B; B = 8'h15; #100;
A = 8'h3B; B = 8'h16; #100;
A = 8'h3B; B = 8'h17; #100;
A = 8'h3B; B = 8'h18; #100;
A = 8'h3B; B = 8'h19; #100;
A = 8'h3B; B = 8'h1A; #100;
A = 8'h3B; B = 8'h1B; #100;
A = 8'h3B; B = 8'h1C; #100;
A = 8'h3B; B = 8'h1D; #100;
A = 8'h3B; B = 8'h1E; #100;
A = 8'h3B; B = 8'h1F; #100;
A = 8'h3B; B = 8'h20; #100;
A = 8'h3B; B = 8'h21; #100;
A = 8'h3B; B = 8'h22; #100;
A = 8'h3B; B = 8'h23; #100;
A = 8'h3B; B = 8'h24; #100;
A = 8'h3B; B = 8'h25; #100;
A = 8'h3B; B = 8'h26; #100;
A = 8'h3B; B = 8'h27; #100;
A = 8'h3B; B = 8'h28; #100;
A = 8'h3B; B = 8'h29; #100;
A = 8'h3B; B = 8'h2A; #100;
A = 8'h3B; B = 8'h2B; #100;
A = 8'h3B; B = 8'h2C; #100;
A = 8'h3B; B = 8'h2D; #100;
A = 8'h3B; B = 8'h2E; #100;
A = 8'h3B; B = 8'h2F; #100;
A = 8'h3B; B = 8'h30; #100;
A = 8'h3B; B = 8'h31; #100;
A = 8'h3B; B = 8'h32; #100;
A = 8'h3B; B = 8'h33; #100;
A = 8'h3B; B = 8'h34; #100;
A = 8'h3B; B = 8'h35; #100;
A = 8'h3B; B = 8'h36; #100;
A = 8'h3B; B = 8'h37; #100;
A = 8'h3B; B = 8'h38; #100;
A = 8'h3B; B = 8'h39; #100;
A = 8'h3B; B = 8'h3A; #100;
A = 8'h3B; B = 8'h3B; #100;
A = 8'h3B; B = 8'h3C; #100;
A = 8'h3B; B = 8'h3D; #100;
A = 8'h3B; B = 8'h3E; #100;
A = 8'h3B; B = 8'h3F; #100;
A = 8'h3B; B = 8'h40; #100;
A = 8'h3B; B = 8'h41; #100;
A = 8'h3B; B = 8'h42; #100;
A = 8'h3B; B = 8'h43; #100;
A = 8'h3B; B = 8'h44; #100;
A = 8'h3B; B = 8'h45; #100;
A = 8'h3B; B = 8'h46; #100;
A = 8'h3B; B = 8'h47; #100;
A = 8'h3B; B = 8'h48; #100;
A = 8'h3B; B = 8'h49; #100;
A = 8'h3B; B = 8'h4A; #100;
A = 8'h3B; B = 8'h4B; #100;
A = 8'h3B; B = 8'h4C; #100;
A = 8'h3B; B = 8'h4D; #100;
A = 8'h3B; B = 8'h4E; #100;
A = 8'h3B; B = 8'h4F; #100;
A = 8'h3B; B = 8'h50; #100;
A = 8'h3B; B = 8'h51; #100;
A = 8'h3B; B = 8'h52; #100;
A = 8'h3B; B = 8'h53; #100;
A = 8'h3B; B = 8'h54; #100;
A = 8'h3B; B = 8'h55; #100;
A = 8'h3B; B = 8'h56; #100;
A = 8'h3B; B = 8'h57; #100;
A = 8'h3B; B = 8'h58; #100;
A = 8'h3B; B = 8'h59; #100;
A = 8'h3B; B = 8'h5A; #100;
A = 8'h3B; B = 8'h5B; #100;
A = 8'h3B; B = 8'h5C; #100;
A = 8'h3B; B = 8'h5D; #100;
A = 8'h3B; B = 8'h5E; #100;
A = 8'h3B; B = 8'h5F; #100;
A = 8'h3B; B = 8'h60; #100;
A = 8'h3B; B = 8'h61; #100;
A = 8'h3B; B = 8'h62; #100;
A = 8'h3B; B = 8'h63; #100;
A = 8'h3B; B = 8'h64; #100;
A = 8'h3B; B = 8'h65; #100;
A = 8'h3B; B = 8'h66; #100;
A = 8'h3B; B = 8'h67; #100;
A = 8'h3B; B = 8'h68; #100;
A = 8'h3B; B = 8'h69; #100;
A = 8'h3B; B = 8'h6A; #100;
A = 8'h3B; B = 8'h6B; #100;
A = 8'h3B; B = 8'h6C; #100;
A = 8'h3B; B = 8'h6D; #100;
A = 8'h3B; B = 8'h6E; #100;
A = 8'h3B; B = 8'h6F; #100;
A = 8'h3B; B = 8'h70; #100;
A = 8'h3B; B = 8'h71; #100;
A = 8'h3B; B = 8'h72; #100;
A = 8'h3B; B = 8'h73; #100;
A = 8'h3B; B = 8'h74; #100;
A = 8'h3B; B = 8'h75; #100;
A = 8'h3B; B = 8'h76; #100;
A = 8'h3B; B = 8'h77; #100;
A = 8'h3B; B = 8'h78; #100;
A = 8'h3B; B = 8'h79; #100;
A = 8'h3B; B = 8'h7A; #100;
A = 8'h3B; B = 8'h7B; #100;
A = 8'h3B; B = 8'h7C; #100;
A = 8'h3B; B = 8'h7D; #100;
A = 8'h3B; B = 8'h7E; #100;
A = 8'h3B; B = 8'h7F; #100;
A = 8'h3B; B = 8'h80; #100;
A = 8'h3B; B = 8'h81; #100;
A = 8'h3B; B = 8'h82; #100;
A = 8'h3B; B = 8'h83; #100;
A = 8'h3B; B = 8'h84; #100;
A = 8'h3B; B = 8'h85; #100;
A = 8'h3B; B = 8'h86; #100;
A = 8'h3B; B = 8'h87; #100;
A = 8'h3B; B = 8'h88; #100;
A = 8'h3B; B = 8'h89; #100;
A = 8'h3B; B = 8'h8A; #100;
A = 8'h3B; B = 8'h8B; #100;
A = 8'h3B; B = 8'h8C; #100;
A = 8'h3B; B = 8'h8D; #100;
A = 8'h3B; B = 8'h8E; #100;
A = 8'h3B; B = 8'h8F; #100;
A = 8'h3B; B = 8'h90; #100;
A = 8'h3B; B = 8'h91; #100;
A = 8'h3B; B = 8'h92; #100;
A = 8'h3B; B = 8'h93; #100;
A = 8'h3B; B = 8'h94; #100;
A = 8'h3B; B = 8'h95; #100;
A = 8'h3B; B = 8'h96; #100;
A = 8'h3B; B = 8'h97; #100;
A = 8'h3B; B = 8'h98; #100;
A = 8'h3B; B = 8'h99; #100;
A = 8'h3B; B = 8'h9A; #100;
A = 8'h3B; B = 8'h9B; #100;
A = 8'h3B; B = 8'h9C; #100;
A = 8'h3B; B = 8'h9D; #100;
A = 8'h3B; B = 8'h9E; #100;
A = 8'h3B; B = 8'h9F; #100;
A = 8'h3B; B = 8'hA0; #100;
A = 8'h3B; B = 8'hA1; #100;
A = 8'h3B; B = 8'hA2; #100;
A = 8'h3B; B = 8'hA3; #100;
A = 8'h3B; B = 8'hA4; #100;
A = 8'h3B; B = 8'hA5; #100;
A = 8'h3B; B = 8'hA6; #100;
A = 8'h3B; B = 8'hA7; #100;
A = 8'h3B; B = 8'hA8; #100;
A = 8'h3B; B = 8'hA9; #100;
A = 8'h3B; B = 8'hAA; #100;
A = 8'h3B; B = 8'hAB; #100;
A = 8'h3B; B = 8'hAC; #100;
A = 8'h3B; B = 8'hAD; #100;
A = 8'h3B; B = 8'hAE; #100;
A = 8'h3B; B = 8'hAF; #100;
A = 8'h3B; B = 8'hB0; #100;
A = 8'h3B; B = 8'hB1; #100;
A = 8'h3B; B = 8'hB2; #100;
A = 8'h3B; B = 8'hB3; #100;
A = 8'h3B; B = 8'hB4; #100;
A = 8'h3B; B = 8'hB5; #100;
A = 8'h3B; B = 8'hB6; #100;
A = 8'h3B; B = 8'hB7; #100;
A = 8'h3B; B = 8'hB8; #100;
A = 8'h3B; B = 8'hB9; #100;
A = 8'h3B; B = 8'hBA; #100;
A = 8'h3B; B = 8'hBB; #100;
A = 8'h3B; B = 8'hBC; #100;
A = 8'h3B; B = 8'hBD; #100;
A = 8'h3B; B = 8'hBE; #100;
A = 8'h3B; B = 8'hBF; #100;
A = 8'h3B; B = 8'hC0; #100;
A = 8'h3B; B = 8'hC1; #100;
A = 8'h3B; B = 8'hC2; #100;
A = 8'h3B; B = 8'hC3; #100;
A = 8'h3B; B = 8'hC4; #100;
A = 8'h3B; B = 8'hC5; #100;
A = 8'h3B; B = 8'hC6; #100;
A = 8'h3B; B = 8'hC7; #100;
A = 8'h3B; B = 8'hC8; #100;
A = 8'h3B; B = 8'hC9; #100;
A = 8'h3B; B = 8'hCA; #100;
A = 8'h3B; B = 8'hCB; #100;
A = 8'h3B; B = 8'hCC; #100;
A = 8'h3B; B = 8'hCD; #100;
A = 8'h3B; B = 8'hCE; #100;
A = 8'h3B; B = 8'hCF; #100;
A = 8'h3B; B = 8'hD0; #100;
A = 8'h3B; B = 8'hD1; #100;
A = 8'h3B; B = 8'hD2; #100;
A = 8'h3B; B = 8'hD3; #100;
A = 8'h3B; B = 8'hD4; #100;
A = 8'h3B; B = 8'hD5; #100;
A = 8'h3B; B = 8'hD6; #100;
A = 8'h3B; B = 8'hD7; #100;
A = 8'h3B; B = 8'hD8; #100;
A = 8'h3B; B = 8'hD9; #100;
A = 8'h3B; B = 8'hDA; #100;
A = 8'h3B; B = 8'hDB; #100;
A = 8'h3B; B = 8'hDC; #100;
A = 8'h3B; B = 8'hDD; #100;
A = 8'h3B; B = 8'hDE; #100;
A = 8'h3B; B = 8'hDF; #100;
A = 8'h3B; B = 8'hE0; #100;
A = 8'h3B; B = 8'hE1; #100;
A = 8'h3B; B = 8'hE2; #100;
A = 8'h3B; B = 8'hE3; #100;
A = 8'h3B; B = 8'hE4; #100;
A = 8'h3B; B = 8'hE5; #100;
A = 8'h3B; B = 8'hE6; #100;
A = 8'h3B; B = 8'hE7; #100;
A = 8'h3B; B = 8'hE8; #100;
A = 8'h3B; B = 8'hE9; #100;
A = 8'h3B; B = 8'hEA; #100;
A = 8'h3B; B = 8'hEB; #100;
A = 8'h3B; B = 8'hEC; #100;
A = 8'h3B; B = 8'hED; #100;
A = 8'h3B; B = 8'hEE; #100;
A = 8'h3B; B = 8'hEF; #100;
A = 8'h3B; B = 8'hF0; #100;
A = 8'h3B; B = 8'hF1; #100;
A = 8'h3B; B = 8'hF2; #100;
A = 8'h3B; B = 8'hF3; #100;
A = 8'h3B; B = 8'hF4; #100;
A = 8'h3B; B = 8'hF5; #100;
A = 8'h3B; B = 8'hF6; #100;
A = 8'h3B; B = 8'hF7; #100;
A = 8'h3B; B = 8'hF8; #100;
A = 8'h3B; B = 8'hF9; #100;
A = 8'h3B; B = 8'hFA; #100;
A = 8'h3B; B = 8'hFB; #100;
A = 8'h3B; B = 8'hFC; #100;
A = 8'h3B; B = 8'hFD; #100;
A = 8'h3B; B = 8'hFE; #100;
A = 8'h3B; B = 8'hFF; #100;
A = 8'h3C; B = 8'h0; #100;
A = 8'h3C; B = 8'h1; #100;
A = 8'h3C; B = 8'h2; #100;
A = 8'h3C; B = 8'h3; #100;
A = 8'h3C; B = 8'h4; #100;
A = 8'h3C; B = 8'h5; #100;
A = 8'h3C; B = 8'h6; #100;
A = 8'h3C; B = 8'h7; #100;
A = 8'h3C; B = 8'h8; #100;
A = 8'h3C; B = 8'h9; #100;
A = 8'h3C; B = 8'hA; #100;
A = 8'h3C; B = 8'hB; #100;
A = 8'h3C; B = 8'hC; #100;
A = 8'h3C; B = 8'hD; #100;
A = 8'h3C; B = 8'hE; #100;
A = 8'h3C; B = 8'hF; #100;
A = 8'h3C; B = 8'h10; #100;
A = 8'h3C; B = 8'h11; #100;
A = 8'h3C; B = 8'h12; #100;
A = 8'h3C; B = 8'h13; #100;
A = 8'h3C; B = 8'h14; #100;
A = 8'h3C; B = 8'h15; #100;
A = 8'h3C; B = 8'h16; #100;
A = 8'h3C; B = 8'h17; #100;
A = 8'h3C; B = 8'h18; #100;
A = 8'h3C; B = 8'h19; #100;
A = 8'h3C; B = 8'h1A; #100;
A = 8'h3C; B = 8'h1B; #100;
A = 8'h3C; B = 8'h1C; #100;
A = 8'h3C; B = 8'h1D; #100;
A = 8'h3C; B = 8'h1E; #100;
A = 8'h3C; B = 8'h1F; #100;
A = 8'h3C; B = 8'h20; #100;
A = 8'h3C; B = 8'h21; #100;
A = 8'h3C; B = 8'h22; #100;
A = 8'h3C; B = 8'h23; #100;
A = 8'h3C; B = 8'h24; #100;
A = 8'h3C; B = 8'h25; #100;
A = 8'h3C; B = 8'h26; #100;
A = 8'h3C; B = 8'h27; #100;
A = 8'h3C; B = 8'h28; #100;
A = 8'h3C; B = 8'h29; #100;
A = 8'h3C; B = 8'h2A; #100;
A = 8'h3C; B = 8'h2B; #100;
A = 8'h3C; B = 8'h2C; #100;
A = 8'h3C; B = 8'h2D; #100;
A = 8'h3C; B = 8'h2E; #100;
A = 8'h3C; B = 8'h2F; #100;
A = 8'h3C; B = 8'h30; #100;
A = 8'h3C; B = 8'h31; #100;
A = 8'h3C; B = 8'h32; #100;
A = 8'h3C; B = 8'h33; #100;
A = 8'h3C; B = 8'h34; #100;
A = 8'h3C; B = 8'h35; #100;
A = 8'h3C; B = 8'h36; #100;
A = 8'h3C; B = 8'h37; #100;
A = 8'h3C; B = 8'h38; #100;
A = 8'h3C; B = 8'h39; #100;
A = 8'h3C; B = 8'h3A; #100;
A = 8'h3C; B = 8'h3B; #100;
A = 8'h3C; B = 8'h3C; #100;
A = 8'h3C; B = 8'h3D; #100;
A = 8'h3C; B = 8'h3E; #100;
A = 8'h3C; B = 8'h3F; #100;
A = 8'h3C; B = 8'h40; #100;
A = 8'h3C; B = 8'h41; #100;
A = 8'h3C; B = 8'h42; #100;
A = 8'h3C; B = 8'h43; #100;
A = 8'h3C; B = 8'h44; #100;
A = 8'h3C; B = 8'h45; #100;
A = 8'h3C; B = 8'h46; #100;
A = 8'h3C; B = 8'h47; #100;
A = 8'h3C; B = 8'h48; #100;
A = 8'h3C; B = 8'h49; #100;
A = 8'h3C; B = 8'h4A; #100;
A = 8'h3C; B = 8'h4B; #100;
A = 8'h3C; B = 8'h4C; #100;
A = 8'h3C; B = 8'h4D; #100;
A = 8'h3C; B = 8'h4E; #100;
A = 8'h3C; B = 8'h4F; #100;
A = 8'h3C; B = 8'h50; #100;
A = 8'h3C; B = 8'h51; #100;
A = 8'h3C; B = 8'h52; #100;
A = 8'h3C; B = 8'h53; #100;
A = 8'h3C; B = 8'h54; #100;
A = 8'h3C; B = 8'h55; #100;
A = 8'h3C; B = 8'h56; #100;
A = 8'h3C; B = 8'h57; #100;
A = 8'h3C; B = 8'h58; #100;
A = 8'h3C; B = 8'h59; #100;
A = 8'h3C; B = 8'h5A; #100;
A = 8'h3C; B = 8'h5B; #100;
A = 8'h3C; B = 8'h5C; #100;
A = 8'h3C; B = 8'h5D; #100;
A = 8'h3C; B = 8'h5E; #100;
A = 8'h3C; B = 8'h5F; #100;
A = 8'h3C; B = 8'h60; #100;
A = 8'h3C; B = 8'h61; #100;
A = 8'h3C; B = 8'h62; #100;
A = 8'h3C; B = 8'h63; #100;
A = 8'h3C; B = 8'h64; #100;
A = 8'h3C; B = 8'h65; #100;
A = 8'h3C; B = 8'h66; #100;
A = 8'h3C; B = 8'h67; #100;
A = 8'h3C; B = 8'h68; #100;
A = 8'h3C; B = 8'h69; #100;
A = 8'h3C; B = 8'h6A; #100;
A = 8'h3C; B = 8'h6B; #100;
A = 8'h3C; B = 8'h6C; #100;
A = 8'h3C; B = 8'h6D; #100;
A = 8'h3C; B = 8'h6E; #100;
A = 8'h3C; B = 8'h6F; #100;
A = 8'h3C; B = 8'h70; #100;
A = 8'h3C; B = 8'h71; #100;
A = 8'h3C; B = 8'h72; #100;
A = 8'h3C; B = 8'h73; #100;
A = 8'h3C; B = 8'h74; #100;
A = 8'h3C; B = 8'h75; #100;
A = 8'h3C; B = 8'h76; #100;
A = 8'h3C; B = 8'h77; #100;
A = 8'h3C; B = 8'h78; #100;
A = 8'h3C; B = 8'h79; #100;
A = 8'h3C; B = 8'h7A; #100;
A = 8'h3C; B = 8'h7B; #100;
A = 8'h3C; B = 8'h7C; #100;
A = 8'h3C; B = 8'h7D; #100;
A = 8'h3C; B = 8'h7E; #100;
A = 8'h3C; B = 8'h7F; #100;
A = 8'h3C; B = 8'h80; #100;
A = 8'h3C; B = 8'h81; #100;
A = 8'h3C; B = 8'h82; #100;
A = 8'h3C; B = 8'h83; #100;
A = 8'h3C; B = 8'h84; #100;
A = 8'h3C; B = 8'h85; #100;
A = 8'h3C; B = 8'h86; #100;
A = 8'h3C; B = 8'h87; #100;
A = 8'h3C; B = 8'h88; #100;
A = 8'h3C; B = 8'h89; #100;
A = 8'h3C; B = 8'h8A; #100;
A = 8'h3C; B = 8'h8B; #100;
A = 8'h3C; B = 8'h8C; #100;
A = 8'h3C; B = 8'h8D; #100;
A = 8'h3C; B = 8'h8E; #100;
A = 8'h3C; B = 8'h8F; #100;
A = 8'h3C; B = 8'h90; #100;
A = 8'h3C; B = 8'h91; #100;
A = 8'h3C; B = 8'h92; #100;
A = 8'h3C; B = 8'h93; #100;
A = 8'h3C; B = 8'h94; #100;
A = 8'h3C; B = 8'h95; #100;
A = 8'h3C; B = 8'h96; #100;
A = 8'h3C; B = 8'h97; #100;
A = 8'h3C; B = 8'h98; #100;
A = 8'h3C; B = 8'h99; #100;
A = 8'h3C; B = 8'h9A; #100;
A = 8'h3C; B = 8'h9B; #100;
A = 8'h3C; B = 8'h9C; #100;
A = 8'h3C; B = 8'h9D; #100;
A = 8'h3C; B = 8'h9E; #100;
A = 8'h3C; B = 8'h9F; #100;
A = 8'h3C; B = 8'hA0; #100;
A = 8'h3C; B = 8'hA1; #100;
A = 8'h3C; B = 8'hA2; #100;
A = 8'h3C; B = 8'hA3; #100;
A = 8'h3C; B = 8'hA4; #100;
A = 8'h3C; B = 8'hA5; #100;
A = 8'h3C; B = 8'hA6; #100;
A = 8'h3C; B = 8'hA7; #100;
A = 8'h3C; B = 8'hA8; #100;
A = 8'h3C; B = 8'hA9; #100;
A = 8'h3C; B = 8'hAA; #100;
A = 8'h3C; B = 8'hAB; #100;
A = 8'h3C; B = 8'hAC; #100;
A = 8'h3C; B = 8'hAD; #100;
A = 8'h3C; B = 8'hAE; #100;
A = 8'h3C; B = 8'hAF; #100;
A = 8'h3C; B = 8'hB0; #100;
A = 8'h3C; B = 8'hB1; #100;
A = 8'h3C; B = 8'hB2; #100;
A = 8'h3C; B = 8'hB3; #100;
A = 8'h3C; B = 8'hB4; #100;
A = 8'h3C; B = 8'hB5; #100;
A = 8'h3C; B = 8'hB6; #100;
A = 8'h3C; B = 8'hB7; #100;
A = 8'h3C; B = 8'hB8; #100;
A = 8'h3C; B = 8'hB9; #100;
A = 8'h3C; B = 8'hBA; #100;
A = 8'h3C; B = 8'hBB; #100;
A = 8'h3C; B = 8'hBC; #100;
A = 8'h3C; B = 8'hBD; #100;
A = 8'h3C; B = 8'hBE; #100;
A = 8'h3C; B = 8'hBF; #100;
A = 8'h3C; B = 8'hC0; #100;
A = 8'h3C; B = 8'hC1; #100;
A = 8'h3C; B = 8'hC2; #100;
A = 8'h3C; B = 8'hC3; #100;
A = 8'h3C; B = 8'hC4; #100;
A = 8'h3C; B = 8'hC5; #100;
A = 8'h3C; B = 8'hC6; #100;
A = 8'h3C; B = 8'hC7; #100;
A = 8'h3C; B = 8'hC8; #100;
A = 8'h3C; B = 8'hC9; #100;
A = 8'h3C; B = 8'hCA; #100;
A = 8'h3C; B = 8'hCB; #100;
A = 8'h3C; B = 8'hCC; #100;
A = 8'h3C; B = 8'hCD; #100;
A = 8'h3C; B = 8'hCE; #100;
A = 8'h3C; B = 8'hCF; #100;
A = 8'h3C; B = 8'hD0; #100;
A = 8'h3C; B = 8'hD1; #100;
A = 8'h3C; B = 8'hD2; #100;
A = 8'h3C; B = 8'hD3; #100;
A = 8'h3C; B = 8'hD4; #100;
A = 8'h3C; B = 8'hD5; #100;
A = 8'h3C; B = 8'hD6; #100;
A = 8'h3C; B = 8'hD7; #100;
A = 8'h3C; B = 8'hD8; #100;
A = 8'h3C; B = 8'hD9; #100;
A = 8'h3C; B = 8'hDA; #100;
A = 8'h3C; B = 8'hDB; #100;
A = 8'h3C; B = 8'hDC; #100;
A = 8'h3C; B = 8'hDD; #100;
A = 8'h3C; B = 8'hDE; #100;
A = 8'h3C; B = 8'hDF; #100;
A = 8'h3C; B = 8'hE0; #100;
A = 8'h3C; B = 8'hE1; #100;
A = 8'h3C; B = 8'hE2; #100;
A = 8'h3C; B = 8'hE3; #100;
A = 8'h3C; B = 8'hE4; #100;
A = 8'h3C; B = 8'hE5; #100;
A = 8'h3C; B = 8'hE6; #100;
A = 8'h3C; B = 8'hE7; #100;
A = 8'h3C; B = 8'hE8; #100;
A = 8'h3C; B = 8'hE9; #100;
A = 8'h3C; B = 8'hEA; #100;
A = 8'h3C; B = 8'hEB; #100;
A = 8'h3C; B = 8'hEC; #100;
A = 8'h3C; B = 8'hED; #100;
A = 8'h3C; B = 8'hEE; #100;
A = 8'h3C; B = 8'hEF; #100;
A = 8'h3C; B = 8'hF0; #100;
A = 8'h3C; B = 8'hF1; #100;
A = 8'h3C; B = 8'hF2; #100;
A = 8'h3C; B = 8'hF3; #100;
A = 8'h3C; B = 8'hF4; #100;
A = 8'h3C; B = 8'hF5; #100;
A = 8'h3C; B = 8'hF6; #100;
A = 8'h3C; B = 8'hF7; #100;
A = 8'h3C; B = 8'hF8; #100;
A = 8'h3C; B = 8'hF9; #100;
A = 8'h3C; B = 8'hFA; #100;
A = 8'h3C; B = 8'hFB; #100;
A = 8'h3C; B = 8'hFC; #100;
A = 8'h3C; B = 8'hFD; #100;
A = 8'h3C; B = 8'hFE; #100;
A = 8'h3C; B = 8'hFF; #100;
A = 8'h3D; B = 8'h0; #100;
A = 8'h3D; B = 8'h1; #100;
A = 8'h3D; B = 8'h2; #100;
A = 8'h3D; B = 8'h3; #100;
A = 8'h3D; B = 8'h4; #100;
A = 8'h3D; B = 8'h5; #100;
A = 8'h3D; B = 8'h6; #100;
A = 8'h3D; B = 8'h7; #100;
A = 8'h3D; B = 8'h8; #100;
A = 8'h3D; B = 8'h9; #100;
A = 8'h3D; B = 8'hA; #100;
A = 8'h3D; B = 8'hB; #100;
A = 8'h3D; B = 8'hC; #100;
A = 8'h3D; B = 8'hD; #100;
A = 8'h3D; B = 8'hE; #100;
A = 8'h3D; B = 8'hF; #100;
A = 8'h3D; B = 8'h10; #100;
A = 8'h3D; B = 8'h11; #100;
A = 8'h3D; B = 8'h12; #100;
A = 8'h3D; B = 8'h13; #100;
A = 8'h3D; B = 8'h14; #100;
A = 8'h3D; B = 8'h15; #100;
A = 8'h3D; B = 8'h16; #100;
A = 8'h3D; B = 8'h17; #100;
A = 8'h3D; B = 8'h18; #100;
A = 8'h3D; B = 8'h19; #100;
A = 8'h3D; B = 8'h1A; #100;
A = 8'h3D; B = 8'h1B; #100;
A = 8'h3D; B = 8'h1C; #100;
A = 8'h3D; B = 8'h1D; #100;
A = 8'h3D; B = 8'h1E; #100;
A = 8'h3D; B = 8'h1F; #100;
A = 8'h3D; B = 8'h20; #100;
A = 8'h3D; B = 8'h21; #100;
A = 8'h3D; B = 8'h22; #100;
A = 8'h3D; B = 8'h23; #100;
A = 8'h3D; B = 8'h24; #100;
A = 8'h3D; B = 8'h25; #100;
A = 8'h3D; B = 8'h26; #100;
A = 8'h3D; B = 8'h27; #100;
A = 8'h3D; B = 8'h28; #100;
A = 8'h3D; B = 8'h29; #100;
A = 8'h3D; B = 8'h2A; #100;
A = 8'h3D; B = 8'h2B; #100;
A = 8'h3D; B = 8'h2C; #100;
A = 8'h3D; B = 8'h2D; #100;
A = 8'h3D; B = 8'h2E; #100;
A = 8'h3D; B = 8'h2F; #100;
A = 8'h3D; B = 8'h30; #100;
A = 8'h3D; B = 8'h31; #100;
A = 8'h3D; B = 8'h32; #100;
A = 8'h3D; B = 8'h33; #100;
A = 8'h3D; B = 8'h34; #100;
A = 8'h3D; B = 8'h35; #100;
A = 8'h3D; B = 8'h36; #100;
A = 8'h3D; B = 8'h37; #100;
A = 8'h3D; B = 8'h38; #100;
A = 8'h3D; B = 8'h39; #100;
A = 8'h3D; B = 8'h3A; #100;
A = 8'h3D; B = 8'h3B; #100;
A = 8'h3D; B = 8'h3C; #100;
A = 8'h3D; B = 8'h3D; #100;
A = 8'h3D; B = 8'h3E; #100;
A = 8'h3D; B = 8'h3F; #100;
A = 8'h3D; B = 8'h40; #100;
A = 8'h3D; B = 8'h41; #100;
A = 8'h3D; B = 8'h42; #100;
A = 8'h3D; B = 8'h43; #100;
A = 8'h3D; B = 8'h44; #100;
A = 8'h3D; B = 8'h45; #100;
A = 8'h3D; B = 8'h46; #100;
A = 8'h3D; B = 8'h47; #100;
A = 8'h3D; B = 8'h48; #100;
A = 8'h3D; B = 8'h49; #100;
A = 8'h3D; B = 8'h4A; #100;
A = 8'h3D; B = 8'h4B; #100;
A = 8'h3D; B = 8'h4C; #100;
A = 8'h3D; B = 8'h4D; #100;
A = 8'h3D; B = 8'h4E; #100;
A = 8'h3D; B = 8'h4F; #100;
A = 8'h3D; B = 8'h50; #100;
A = 8'h3D; B = 8'h51; #100;
A = 8'h3D; B = 8'h52; #100;
A = 8'h3D; B = 8'h53; #100;
A = 8'h3D; B = 8'h54; #100;
A = 8'h3D; B = 8'h55; #100;
A = 8'h3D; B = 8'h56; #100;
A = 8'h3D; B = 8'h57; #100;
A = 8'h3D; B = 8'h58; #100;
A = 8'h3D; B = 8'h59; #100;
A = 8'h3D; B = 8'h5A; #100;
A = 8'h3D; B = 8'h5B; #100;
A = 8'h3D; B = 8'h5C; #100;
A = 8'h3D; B = 8'h5D; #100;
A = 8'h3D; B = 8'h5E; #100;
A = 8'h3D; B = 8'h5F; #100;
A = 8'h3D; B = 8'h60; #100;
A = 8'h3D; B = 8'h61; #100;
A = 8'h3D; B = 8'h62; #100;
A = 8'h3D; B = 8'h63; #100;
A = 8'h3D; B = 8'h64; #100;
A = 8'h3D; B = 8'h65; #100;
A = 8'h3D; B = 8'h66; #100;
A = 8'h3D; B = 8'h67; #100;
A = 8'h3D; B = 8'h68; #100;
A = 8'h3D; B = 8'h69; #100;
A = 8'h3D; B = 8'h6A; #100;
A = 8'h3D; B = 8'h6B; #100;
A = 8'h3D; B = 8'h6C; #100;
A = 8'h3D; B = 8'h6D; #100;
A = 8'h3D; B = 8'h6E; #100;
A = 8'h3D; B = 8'h6F; #100;
A = 8'h3D; B = 8'h70; #100;
A = 8'h3D; B = 8'h71; #100;
A = 8'h3D; B = 8'h72; #100;
A = 8'h3D; B = 8'h73; #100;
A = 8'h3D; B = 8'h74; #100;
A = 8'h3D; B = 8'h75; #100;
A = 8'h3D; B = 8'h76; #100;
A = 8'h3D; B = 8'h77; #100;
A = 8'h3D; B = 8'h78; #100;
A = 8'h3D; B = 8'h79; #100;
A = 8'h3D; B = 8'h7A; #100;
A = 8'h3D; B = 8'h7B; #100;
A = 8'h3D; B = 8'h7C; #100;
A = 8'h3D; B = 8'h7D; #100;
A = 8'h3D; B = 8'h7E; #100;
A = 8'h3D; B = 8'h7F; #100;
A = 8'h3D; B = 8'h80; #100;
A = 8'h3D; B = 8'h81; #100;
A = 8'h3D; B = 8'h82; #100;
A = 8'h3D; B = 8'h83; #100;
A = 8'h3D; B = 8'h84; #100;
A = 8'h3D; B = 8'h85; #100;
A = 8'h3D; B = 8'h86; #100;
A = 8'h3D; B = 8'h87; #100;
A = 8'h3D; B = 8'h88; #100;
A = 8'h3D; B = 8'h89; #100;
A = 8'h3D; B = 8'h8A; #100;
A = 8'h3D; B = 8'h8B; #100;
A = 8'h3D; B = 8'h8C; #100;
A = 8'h3D; B = 8'h8D; #100;
A = 8'h3D; B = 8'h8E; #100;
A = 8'h3D; B = 8'h8F; #100;
A = 8'h3D; B = 8'h90; #100;
A = 8'h3D; B = 8'h91; #100;
A = 8'h3D; B = 8'h92; #100;
A = 8'h3D; B = 8'h93; #100;
A = 8'h3D; B = 8'h94; #100;
A = 8'h3D; B = 8'h95; #100;
A = 8'h3D; B = 8'h96; #100;
A = 8'h3D; B = 8'h97; #100;
A = 8'h3D; B = 8'h98; #100;
A = 8'h3D; B = 8'h99; #100;
A = 8'h3D; B = 8'h9A; #100;
A = 8'h3D; B = 8'h9B; #100;
A = 8'h3D; B = 8'h9C; #100;
A = 8'h3D; B = 8'h9D; #100;
A = 8'h3D; B = 8'h9E; #100;
A = 8'h3D; B = 8'h9F; #100;
A = 8'h3D; B = 8'hA0; #100;
A = 8'h3D; B = 8'hA1; #100;
A = 8'h3D; B = 8'hA2; #100;
A = 8'h3D; B = 8'hA3; #100;
A = 8'h3D; B = 8'hA4; #100;
A = 8'h3D; B = 8'hA5; #100;
A = 8'h3D; B = 8'hA6; #100;
A = 8'h3D; B = 8'hA7; #100;
A = 8'h3D; B = 8'hA8; #100;
A = 8'h3D; B = 8'hA9; #100;
A = 8'h3D; B = 8'hAA; #100;
A = 8'h3D; B = 8'hAB; #100;
A = 8'h3D; B = 8'hAC; #100;
A = 8'h3D; B = 8'hAD; #100;
A = 8'h3D; B = 8'hAE; #100;
A = 8'h3D; B = 8'hAF; #100;
A = 8'h3D; B = 8'hB0; #100;
A = 8'h3D; B = 8'hB1; #100;
A = 8'h3D; B = 8'hB2; #100;
A = 8'h3D; B = 8'hB3; #100;
A = 8'h3D; B = 8'hB4; #100;
A = 8'h3D; B = 8'hB5; #100;
A = 8'h3D; B = 8'hB6; #100;
A = 8'h3D; B = 8'hB7; #100;
A = 8'h3D; B = 8'hB8; #100;
A = 8'h3D; B = 8'hB9; #100;
A = 8'h3D; B = 8'hBA; #100;
A = 8'h3D; B = 8'hBB; #100;
A = 8'h3D; B = 8'hBC; #100;
A = 8'h3D; B = 8'hBD; #100;
A = 8'h3D; B = 8'hBE; #100;
A = 8'h3D; B = 8'hBF; #100;
A = 8'h3D; B = 8'hC0; #100;
A = 8'h3D; B = 8'hC1; #100;
A = 8'h3D; B = 8'hC2; #100;
A = 8'h3D; B = 8'hC3; #100;
A = 8'h3D; B = 8'hC4; #100;
A = 8'h3D; B = 8'hC5; #100;
A = 8'h3D; B = 8'hC6; #100;
A = 8'h3D; B = 8'hC7; #100;
A = 8'h3D; B = 8'hC8; #100;
A = 8'h3D; B = 8'hC9; #100;
A = 8'h3D; B = 8'hCA; #100;
A = 8'h3D; B = 8'hCB; #100;
A = 8'h3D; B = 8'hCC; #100;
A = 8'h3D; B = 8'hCD; #100;
A = 8'h3D; B = 8'hCE; #100;
A = 8'h3D; B = 8'hCF; #100;
A = 8'h3D; B = 8'hD0; #100;
A = 8'h3D; B = 8'hD1; #100;
A = 8'h3D; B = 8'hD2; #100;
A = 8'h3D; B = 8'hD3; #100;
A = 8'h3D; B = 8'hD4; #100;
A = 8'h3D; B = 8'hD5; #100;
A = 8'h3D; B = 8'hD6; #100;
A = 8'h3D; B = 8'hD7; #100;
A = 8'h3D; B = 8'hD8; #100;
A = 8'h3D; B = 8'hD9; #100;
A = 8'h3D; B = 8'hDA; #100;
A = 8'h3D; B = 8'hDB; #100;
A = 8'h3D; B = 8'hDC; #100;
A = 8'h3D; B = 8'hDD; #100;
A = 8'h3D; B = 8'hDE; #100;
A = 8'h3D; B = 8'hDF; #100;
A = 8'h3D; B = 8'hE0; #100;
A = 8'h3D; B = 8'hE1; #100;
A = 8'h3D; B = 8'hE2; #100;
A = 8'h3D; B = 8'hE3; #100;
A = 8'h3D; B = 8'hE4; #100;
A = 8'h3D; B = 8'hE5; #100;
A = 8'h3D; B = 8'hE6; #100;
A = 8'h3D; B = 8'hE7; #100;
A = 8'h3D; B = 8'hE8; #100;
A = 8'h3D; B = 8'hE9; #100;
A = 8'h3D; B = 8'hEA; #100;
A = 8'h3D; B = 8'hEB; #100;
A = 8'h3D; B = 8'hEC; #100;
A = 8'h3D; B = 8'hED; #100;
A = 8'h3D; B = 8'hEE; #100;
A = 8'h3D; B = 8'hEF; #100;
A = 8'h3D; B = 8'hF0; #100;
A = 8'h3D; B = 8'hF1; #100;
A = 8'h3D; B = 8'hF2; #100;
A = 8'h3D; B = 8'hF3; #100;
A = 8'h3D; B = 8'hF4; #100;
A = 8'h3D; B = 8'hF5; #100;
A = 8'h3D; B = 8'hF6; #100;
A = 8'h3D; B = 8'hF7; #100;
A = 8'h3D; B = 8'hF8; #100;
A = 8'h3D; B = 8'hF9; #100;
A = 8'h3D; B = 8'hFA; #100;
A = 8'h3D; B = 8'hFB; #100;
A = 8'h3D; B = 8'hFC; #100;
A = 8'h3D; B = 8'hFD; #100;
A = 8'h3D; B = 8'hFE; #100;
A = 8'h3D; B = 8'hFF; #100;
A = 8'h3E; B = 8'h0; #100;
A = 8'h3E; B = 8'h1; #100;
A = 8'h3E; B = 8'h2; #100;
A = 8'h3E; B = 8'h3; #100;
A = 8'h3E; B = 8'h4; #100;
A = 8'h3E; B = 8'h5; #100;
A = 8'h3E; B = 8'h6; #100;
A = 8'h3E; B = 8'h7; #100;
A = 8'h3E; B = 8'h8; #100;
A = 8'h3E; B = 8'h9; #100;
A = 8'h3E; B = 8'hA; #100;
A = 8'h3E; B = 8'hB; #100;
A = 8'h3E; B = 8'hC; #100;
A = 8'h3E; B = 8'hD; #100;
A = 8'h3E; B = 8'hE; #100;
A = 8'h3E; B = 8'hF; #100;
A = 8'h3E; B = 8'h10; #100;
A = 8'h3E; B = 8'h11; #100;
A = 8'h3E; B = 8'h12; #100;
A = 8'h3E; B = 8'h13; #100;
A = 8'h3E; B = 8'h14; #100;
A = 8'h3E; B = 8'h15; #100;
A = 8'h3E; B = 8'h16; #100;
A = 8'h3E; B = 8'h17; #100;
A = 8'h3E; B = 8'h18; #100;
A = 8'h3E; B = 8'h19; #100;
A = 8'h3E; B = 8'h1A; #100;
A = 8'h3E; B = 8'h1B; #100;
A = 8'h3E; B = 8'h1C; #100;
A = 8'h3E; B = 8'h1D; #100;
A = 8'h3E; B = 8'h1E; #100;
A = 8'h3E; B = 8'h1F; #100;
A = 8'h3E; B = 8'h20; #100;
A = 8'h3E; B = 8'h21; #100;
A = 8'h3E; B = 8'h22; #100;
A = 8'h3E; B = 8'h23; #100;
A = 8'h3E; B = 8'h24; #100;
A = 8'h3E; B = 8'h25; #100;
A = 8'h3E; B = 8'h26; #100;
A = 8'h3E; B = 8'h27; #100;
A = 8'h3E; B = 8'h28; #100;
A = 8'h3E; B = 8'h29; #100;
A = 8'h3E; B = 8'h2A; #100;
A = 8'h3E; B = 8'h2B; #100;
A = 8'h3E; B = 8'h2C; #100;
A = 8'h3E; B = 8'h2D; #100;
A = 8'h3E; B = 8'h2E; #100;
A = 8'h3E; B = 8'h2F; #100;
A = 8'h3E; B = 8'h30; #100;
A = 8'h3E; B = 8'h31; #100;
A = 8'h3E; B = 8'h32; #100;
A = 8'h3E; B = 8'h33; #100;
A = 8'h3E; B = 8'h34; #100;
A = 8'h3E; B = 8'h35; #100;
A = 8'h3E; B = 8'h36; #100;
A = 8'h3E; B = 8'h37; #100;
A = 8'h3E; B = 8'h38; #100;
A = 8'h3E; B = 8'h39; #100;
A = 8'h3E; B = 8'h3A; #100;
A = 8'h3E; B = 8'h3B; #100;
A = 8'h3E; B = 8'h3C; #100;
A = 8'h3E; B = 8'h3D; #100;
A = 8'h3E; B = 8'h3E; #100;
A = 8'h3E; B = 8'h3F; #100;
A = 8'h3E; B = 8'h40; #100;
A = 8'h3E; B = 8'h41; #100;
A = 8'h3E; B = 8'h42; #100;
A = 8'h3E; B = 8'h43; #100;
A = 8'h3E; B = 8'h44; #100;
A = 8'h3E; B = 8'h45; #100;
A = 8'h3E; B = 8'h46; #100;
A = 8'h3E; B = 8'h47; #100;
A = 8'h3E; B = 8'h48; #100;
A = 8'h3E; B = 8'h49; #100;
A = 8'h3E; B = 8'h4A; #100;
A = 8'h3E; B = 8'h4B; #100;
A = 8'h3E; B = 8'h4C; #100;
A = 8'h3E; B = 8'h4D; #100;
A = 8'h3E; B = 8'h4E; #100;
A = 8'h3E; B = 8'h4F; #100;
A = 8'h3E; B = 8'h50; #100;
A = 8'h3E; B = 8'h51; #100;
A = 8'h3E; B = 8'h52; #100;
A = 8'h3E; B = 8'h53; #100;
A = 8'h3E; B = 8'h54; #100;
A = 8'h3E; B = 8'h55; #100;
A = 8'h3E; B = 8'h56; #100;
A = 8'h3E; B = 8'h57; #100;
A = 8'h3E; B = 8'h58; #100;
A = 8'h3E; B = 8'h59; #100;
A = 8'h3E; B = 8'h5A; #100;
A = 8'h3E; B = 8'h5B; #100;
A = 8'h3E; B = 8'h5C; #100;
A = 8'h3E; B = 8'h5D; #100;
A = 8'h3E; B = 8'h5E; #100;
A = 8'h3E; B = 8'h5F; #100;
A = 8'h3E; B = 8'h60; #100;
A = 8'h3E; B = 8'h61; #100;
A = 8'h3E; B = 8'h62; #100;
A = 8'h3E; B = 8'h63; #100;
A = 8'h3E; B = 8'h64; #100;
A = 8'h3E; B = 8'h65; #100;
A = 8'h3E; B = 8'h66; #100;
A = 8'h3E; B = 8'h67; #100;
A = 8'h3E; B = 8'h68; #100;
A = 8'h3E; B = 8'h69; #100;
A = 8'h3E; B = 8'h6A; #100;
A = 8'h3E; B = 8'h6B; #100;
A = 8'h3E; B = 8'h6C; #100;
A = 8'h3E; B = 8'h6D; #100;
A = 8'h3E; B = 8'h6E; #100;
A = 8'h3E; B = 8'h6F; #100;
A = 8'h3E; B = 8'h70; #100;
A = 8'h3E; B = 8'h71; #100;
A = 8'h3E; B = 8'h72; #100;
A = 8'h3E; B = 8'h73; #100;
A = 8'h3E; B = 8'h74; #100;
A = 8'h3E; B = 8'h75; #100;
A = 8'h3E; B = 8'h76; #100;
A = 8'h3E; B = 8'h77; #100;
A = 8'h3E; B = 8'h78; #100;
A = 8'h3E; B = 8'h79; #100;
A = 8'h3E; B = 8'h7A; #100;
A = 8'h3E; B = 8'h7B; #100;
A = 8'h3E; B = 8'h7C; #100;
A = 8'h3E; B = 8'h7D; #100;
A = 8'h3E; B = 8'h7E; #100;
A = 8'h3E; B = 8'h7F; #100;
A = 8'h3E; B = 8'h80; #100;
A = 8'h3E; B = 8'h81; #100;
A = 8'h3E; B = 8'h82; #100;
A = 8'h3E; B = 8'h83; #100;
A = 8'h3E; B = 8'h84; #100;
A = 8'h3E; B = 8'h85; #100;
A = 8'h3E; B = 8'h86; #100;
A = 8'h3E; B = 8'h87; #100;
A = 8'h3E; B = 8'h88; #100;
A = 8'h3E; B = 8'h89; #100;
A = 8'h3E; B = 8'h8A; #100;
A = 8'h3E; B = 8'h8B; #100;
A = 8'h3E; B = 8'h8C; #100;
A = 8'h3E; B = 8'h8D; #100;
A = 8'h3E; B = 8'h8E; #100;
A = 8'h3E; B = 8'h8F; #100;
A = 8'h3E; B = 8'h90; #100;
A = 8'h3E; B = 8'h91; #100;
A = 8'h3E; B = 8'h92; #100;
A = 8'h3E; B = 8'h93; #100;
A = 8'h3E; B = 8'h94; #100;
A = 8'h3E; B = 8'h95; #100;
A = 8'h3E; B = 8'h96; #100;
A = 8'h3E; B = 8'h97; #100;
A = 8'h3E; B = 8'h98; #100;
A = 8'h3E; B = 8'h99; #100;
A = 8'h3E; B = 8'h9A; #100;
A = 8'h3E; B = 8'h9B; #100;
A = 8'h3E; B = 8'h9C; #100;
A = 8'h3E; B = 8'h9D; #100;
A = 8'h3E; B = 8'h9E; #100;
A = 8'h3E; B = 8'h9F; #100;
A = 8'h3E; B = 8'hA0; #100;
A = 8'h3E; B = 8'hA1; #100;
A = 8'h3E; B = 8'hA2; #100;
A = 8'h3E; B = 8'hA3; #100;
A = 8'h3E; B = 8'hA4; #100;
A = 8'h3E; B = 8'hA5; #100;
A = 8'h3E; B = 8'hA6; #100;
A = 8'h3E; B = 8'hA7; #100;
A = 8'h3E; B = 8'hA8; #100;
A = 8'h3E; B = 8'hA9; #100;
A = 8'h3E; B = 8'hAA; #100;
A = 8'h3E; B = 8'hAB; #100;
A = 8'h3E; B = 8'hAC; #100;
A = 8'h3E; B = 8'hAD; #100;
A = 8'h3E; B = 8'hAE; #100;
A = 8'h3E; B = 8'hAF; #100;
A = 8'h3E; B = 8'hB0; #100;
A = 8'h3E; B = 8'hB1; #100;
A = 8'h3E; B = 8'hB2; #100;
A = 8'h3E; B = 8'hB3; #100;
A = 8'h3E; B = 8'hB4; #100;
A = 8'h3E; B = 8'hB5; #100;
A = 8'h3E; B = 8'hB6; #100;
A = 8'h3E; B = 8'hB7; #100;
A = 8'h3E; B = 8'hB8; #100;
A = 8'h3E; B = 8'hB9; #100;
A = 8'h3E; B = 8'hBA; #100;
A = 8'h3E; B = 8'hBB; #100;
A = 8'h3E; B = 8'hBC; #100;
A = 8'h3E; B = 8'hBD; #100;
A = 8'h3E; B = 8'hBE; #100;
A = 8'h3E; B = 8'hBF; #100;
A = 8'h3E; B = 8'hC0; #100;
A = 8'h3E; B = 8'hC1; #100;
A = 8'h3E; B = 8'hC2; #100;
A = 8'h3E; B = 8'hC3; #100;
A = 8'h3E; B = 8'hC4; #100;
A = 8'h3E; B = 8'hC5; #100;
A = 8'h3E; B = 8'hC6; #100;
A = 8'h3E; B = 8'hC7; #100;
A = 8'h3E; B = 8'hC8; #100;
A = 8'h3E; B = 8'hC9; #100;
A = 8'h3E; B = 8'hCA; #100;
A = 8'h3E; B = 8'hCB; #100;
A = 8'h3E; B = 8'hCC; #100;
A = 8'h3E; B = 8'hCD; #100;
A = 8'h3E; B = 8'hCE; #100;
A = 8'h3E; B = 8'hCF; #100;
A = 8'h3E; B = 8'hD0; #100;
A = 8'h3E; B = 8'hD1; #100;
A = 8'h3E; B = 8'hD2; #100;
A = 8'h3E; B = 8'hD3; #100;
A = 8'h3E; B = 8'hD4; #100;
A = 8'h3E; B = 8'hD5; #100;
A = 8'h3E; B = 8'hD6; #100;
A = 8'h3E; B = 8'hD7; #100;
A = 8'h3E; B = 8'hD8; #100;
A = 8'h3E; B = 8'hD9; #100;
A = 8'h3E; B = 8'hDA; #100;
A = 8'h3E; B = 8'hDB; #100;
A = 8'h3E; B = 8'hDC; #100;
A = 8'h3E; B = 8'hDD; #100;
A = 8'h3E; B = 8'hDE; #100;
A = 8'h3E; B = 8'hDF; #100;
A = 8'h3E; B = 8'hE0; #100;
A = 8'h3E; B = 8'hE1; #100;
A = 8'h3E; B = 8'hE2; #100;
A = 8'h3E; B = 8'hE3; #100;
A = 8'h3E; B = 8'hE4; #100;
A = 8'h3E; B = 8'hE5; #100;
A = 8'h3E; B = 8'hE6; #100;
A = 8'h3E; B = 8'hE7; #100;
A = 8'h3E; B = 8'hE8; #100;
A = 8'h3E; B = 8'hE9; #100;
A = 8'h3E; B = 8'hEA; #100;
A = 8'h3E; B = 8'hEB; #100;
A = 8'h3E; B = 8'hEC; #100;
A = 8'h3E; B = 8'hED; #100;
A = 8'h3E; B = 8'hEE; #100;
A = 8'h3E; B = 8'hEF; #100;
A = 8'h3E; B = 8'hF0; #100;
A = 8'h3E; B = 8'hF1; #100;
A = 8'h3E; B = 8'hF2; #100;
A = 8'h3E; B = 8'hF3; #100;
A = 8'h3E; B = 8'hF4; #100;
A = 8'h3E; B = 8'hF5; #100;
A = 8'h3E; B = 8'hF6; #100;
A = 8'h3E; B = 8'hF7; #100;
A = 8'h3E; B = 8'hF8; #100;
A = 8'h3E; B = 8'hF9; #100;
A = 8'h3E; B = 8'hFA; #100;
A = 8'h3E; B = 8'hFB; #100;
A = 8'h3E; B = 8'hFC; #100;
A = 8'h3E; B = 8'hFD; #100;
A = 8'h3E; B = 8'hFE; #100;
A = 8'h3E; B = 8'hFF; #100;
A = 8'h3F; B = 8'h0; #100;
A = 8'h3F; B = 8'h1; #100;
A = 8'h3F; B = 8'h2; #100;
A = 8'h3F; B = 8'h3; #100;
A = 8'h3F; B = 8'h4; #100;
A = 8'h3F; B = 8'h5; #100;
A = 8'h3F; B = 8'h6; #100;
A = 8'h3F; B = 8'h7; #100;
A = 8'h3F; B = 8'h8; #100;
A = 8'h3F; B = 8'h9; #100;
A = 8'h3F; B = 8'hA; #100;
A = 8'h3F; B = 8'hB; #100;
A = 8'h3F; B = 8'hC; #100;
A = 8'h3F; B = 8'hD; #100;
A = 8'h3F; B = 8'hE; #100;
A = 8'h3F; B = 8'hF; #100;
A = 8'h3F; B = 8'h10; #100;
A = 8'h3F; B = 8'h11; #100;
A = 8'h3F; B = 8'h12; #100;
A = 8'h3F; B = 8'h13; #100;
A = 8'h3F; B = 8'h14; #100;
A = 8'h3F; B = 8'h15; #100;
A = 8'h3F; B = 8'h16; #100;
A = 8'h3F; B = 8'h17; #100;
A = 8'h3F; B = 8'h18; #100;
A = 8'h3F; B = 8'h19; #100;
A = 8'h3F; B = 8'h1A; #100;
A = 8'h3F; B = 8'h1B; #100;
A = 8'h3F; B = 8'h1C; #100;
A = 8'h3F; B = 8'h1D; #100;
A = 8'h3F; B = 8'h1E; #100;
A = 8'h3F; B = 8'h1F; #100;
A = 8'h3F; B = 8'h20; #100;
A = 8'h3F; B = 8'h21; #100;
A = 8'h3F; B = 8'h22; #100;
A = 8'h3F; B = 8'h23; #100;
A = 8'h3F; B = 8'h24; #100;
A = 8'h3F; B = 8'h25; #100;
A = 8'h3F; B = 8'h26; #100;
A = 8'h3F; B = 8'h27; #100;
A = 8'h3F; B = 8'h28; #100;
A = 8'h3F; B = 8'h29; #100;
A = 8'h3F; B = 8'h2A; #100;
A = 8'h3F; B = 8'h2B; #100;
A = 8'h3F; B = 8'h2C; #100;
A = 8'h3F; B = 8'h2D; #100;
A = 8'h3F; B = 8'h2E; #100;
A = 8'h3F; B = 8'h2F; #100;
A = 8'h3F; B = 8'h30; #100;
A = 8'h3F; B = 8'h31; #100;
A = 8'h3F; B = 8'h32; #100;
A = 8'h3F; B = 8'h33; #100;
A = 8'h3F; B = 8'h34; #100;
A = 8'h3F; B = 8'h35; #100;
A = 8'h3F; B = 8'h36; #100;
A = 8'h3F; B = 8'h37; #100;
A = 8'h3F; B = 8'h38; #100;
A = 8'h3F; B = 8'h39; #100;
A = 8'h3F; B = 8'h3A; #100;
A = 8'h3F; B = 8'h3B; #100;
A = 8'h3F; B = 8'h3C; #100;
A = 8'h3F; B = 8'h3D; #100;
A = 8'h3F; B = 8'h3E; #100;
A = 8'h3F; B = 8'h3F; #100;
A = 8'h3F; B = 8'h40; #100;
A = 8'h3F; B = 8'h41; #100;
A = 8'h3F; B = 8'h42; #100;
A = 8'h3F; B = 8'h43; #100;
A = 8'h3F; B = 8'h44; #100;
A = 8'h3F; B = 8'h45; #100;
A = 8'h3F; B = 8'h46; #100;
A = 8'h3F; B = 8'h47; #100;
A = 8'h3F; B = 8'h48; #100;
A = 8'h3F; B = 8'h49; #100;
A = 8'h3F; B = 8'h4A; #100;
A = 8'h3F; B = 8'h4B; #100;
A = 8'h3F; B = 8'h4C; #100;
A = 8'h3F; B = 8'h4D; #100;
A = 8'h3F; B = 8'h4E; #100;
A = 8'h3F; B = 8'h4F; #100;
A = 8'h3F; B = 8'h50; #100;
A = 8'h3F; B = 8'h51; #100;
A = 8'h3F; B = 8'h52; #100;
A = 8'h3F; B = 8'h53; #100;
A = 8'h3F; B = 8'h54; #100;
A = 8'h3F; B = 8'h55; #100;
A = 8'h3F; B = 8'h56; #100;
A = 8'h3F; B = 8'h57; #100;
A = 8'h3F; B = 8'h58; #100;
A = 8'h3F; B = 8'h59; #100;
A = 8'h3F; B = 8'h5A; #100;
A = 8'h3F; B = 8'h5B; #100;
A = 8'h3F; B = 8'h5C; #100;
A = 8'h3F; B = 8'h5D; #100;
A = 8'h3F; B = 8'h5E; #100;
A = 8'h3F; B = 8'h5F; #100;
A = 8'h3F; B = 8'h60; #100;
A = 8'h3F; B = 8'h61; #100;
A = 8'h3F; B = 8'h62; #100;
A = 8'h3F; B = 8'h63; #100;
A = 8'h3F; B = 8'h64; #100;
A = 8'h3F; B = 8'h65; #100;
A = 8'h3F; B = 8'h66; #100;
A = 8'h3F; B = 8'h67; #100;
A = 8'h3F; B = 8'h68; #100;
A = 8'h3F; B = 8'h69; #100;
A = 8'h3F; B = 8'h6A; #100;
A = 8'h3F; B = 8'h6B; #100;
A = 8'h3F; B = 8'h6C; #100;
A = 8'h3F; B = 8'h6D; #100;
A = 8'h3F; B = 8'h6E; #100;
A = 8'h3F; B = 8'h6F; #100;
A = 8'h3F; B = 8'h70; #100;
A = 8'h3F; B = 8'h71; #100;
A = 8'h3F; B = 8'h72; #100;
A = 8'h3F; B = 8'h73; #100;
A = 8'h3F; B = 8'h74; #100;
A = 8'h3F; B = 8'h75; #100;
A = 8'h3F; B = 8'h76; #100;
A = 8'h3F; B = 8'h77; #100;
A = 8'h3F; B = 8'h78; #100;
A = 8'h3F; B = 8'h79; #100;
A = 8'h3F; B = 8'h7A; #100;
A = 8'h3F; B = 8'h7B; #100;
A = 8'h3F; B = 8'h7C; #100;
A = 8'h3F; B = 8'h7D; #100;
A = 8'h3F; B = 8'h7E; #100;
A = 8'h3F; B = 8'h7F; #100;
A = 8'h3F; B = 8'h80; #100;
A = 8'h3F; B = 8'h81; #100;
A = 8'h3F; B = 8'h82; #100;
A = 8'h3F; B = 8'h83; #100;
A = 8'h3F; B = 8'h84; #100;
A = 8'h3F; B = 8'h85; #100;
A = 8'h3F; B = 8'h86; #100;
A = 8'h3F; B = 8'h87; #100;
A = 8'h3F; B = 8'h88; #100;
A = 8'h3F; B = 8'h89; #100;
A = 8'h3F; B = 8'h8A; #100;
A = 8'h3F; B = 8'h8B; #100;
A = 8'h3F; B = 8'h8C; #100;
A = 8'h3F; B = 8'h8D; #100;
A = 8'h3F; B = 8'h8E; #100;
A = 8'h3F; B = 8'h8F; #100;
A = 8'h3F; B = 8'h90; #100;
A = 8'h3F; B = 8'h91; #100;
A = 8'h3F; B = 8'h92; #100;
A = 8'h3F; B = 8'h93; #100;
A = 8'h3F; B = 8'h94; #100;
A = 8'h3F; B = 8'h95; #100;
A = 8'h3F; B = 8'h96; #100;
A = 8'h3F; B = 8'h97; #100;
A = 8'h3F; B = 8'h98; #100;
A = 8'h3F; B = 8'h99; #100;
A = 8'h3F; B = 8'h9A; #100;
A = 8'h3F; B = 8'h9B; #100;
A = 8'h3F; B = 8'h9C; #100;
A = 8'h3F; B = 8'h9D; #100;
A = 8'h3F; B = 8'h9E; #100;
A = 8'h3F; B = 8'h9F; #100;
A = 8'h3F; B = 8'hA0; #100;
A = 8'h3F; B = 8'hA1; #100;
A = 8'h3F; B = 8'hA2; #100;
A = 8'h3F; B = 8'hA3; #100;
A = 8'h3F; B = 8'hA4; #100;
A = 8'h3F; B = 8'hA5; #100;
A = 8'h3F; B = 8'hA6; #100;
A = 8'h3F; B = 8'hA7; #100;
A = 8'h3F; B = 8'hA8; #100;
A = 8'h3F; B = 8'hA9; #100;
A = 8'h3F; B = 8'hAA; #100;
A = 8'h3F; B = 8'hAB; #100;
A = 8'h3F; B = 8'hAC; #100;
A = 8'h3F; B = 8'hAD; #100;
A = 8'h3F; B = 8'hAE; #100;
A = 8'h3F; B = 8'hAF; #100;
A = 8'h3F; B = 8'hB0; #100;
A = 8'h3F; B = 8'hB1; #100;
A = 8'h3F; B = 8'hB2; #100;
A = 8'h3F; B = 8'hB3; #100;
A = 8'h3F; B = 8'hB4; #100;
A = 8'h3F; B = 8'hB5; #100;
A = 8'h3F; B = 8'hB6; #100;
A = 8'h3F; B = 8'hB7; #100;
A = 8'h3F; B = 8'hB8; #100;
A = 8'h3F; B = 8'hB9; #100;
A = 8'h3F; B = 8'hBA; #100;
A = 8'h3F; B = 8'hBB; #100;
A = 8'h3F; B = 8'hBC; #100;
A = 8'h3F; B = 8'hBD; #100;
A = 8'h3F; B = 8'hBE; #100;
A = 8'h3F; B = 8'hBF; #100;
A = 8'h3F; B = 8'hC0; #100;
A = 8'h3F; B = 8'hC1; #100;
A = 8'h3F; B = 8'hC2; #100;
A = 8'h3F; B = 8'hC3; #100;
A = 8'h3F; B = 8'hC4; #100;
A = 8'h3F; B = 8'hC5; #100;
A = 8'h3F; B = 8'hC6; #100;
A = 8'h3F; B = 8'hC7; #100;
A = 8'h3F; B = 8'hC8; #100;
A = 8'h3F; B = 8'hC9; #100;
A = 8'h3F; B = 8'hCA; #100;
A = 8'h3F; B = 8'hCB; #100;
A = 8'h3F; B = 8'hCC; #100;
A = 8'h3F; B = 8'hCD; #100;
A = 8'h3F; B = 8'hCE; #100;
A = 8'h3F; B = 8'hCF; #100;
A = 8'h3F; B = 8'hD0; #100;
A = 8'h3F; B = 8'hD1; #100;
A = 8'h3F; B = 8'hD2; #100;
A = 8'h3F; B = 8'hD3; #100;
A = 8'h3F; B = 8'hD4; #100;
A = 8'h3F; B = 8'hD5; #100;
A = 8'h3F; B = 8'hD6; #100;
A = 8'h3F; B = 8'hD7; #100;
A = 8'h3F; B = 8'hD8; #100;
A = 8'h3F; B = 8'hD9; #100;
A = 8'h3F; B = 8'hDA; #100;
A = 8'h3F; B = 8'hDB; #100;
A = 8'h3F; B = 8'hDC; #100;
A = 8'h3F; B = 8'hDD; #100;
A = 8'h3F; B = 8'hDE; #100;
A = 8'h3F; B = 8'hDF; #100;
A = 8'h3F; B = 8'hE0; #100;
A = 8'h3F; B = 8'hE1; #100;
A = 8'h3F; B = 8'hE2; #100;
A = 8'h3F; B = 8'hE3; #100;
A = 8'h3F; B = 8'hE4; #100;
A = 8'h3F; B = 8'hE5; #100;
A = 8'h3F; B = 8'hE6; #100;
A = 8'h3F; B = 8'hE7; #100;
A = 8'h3F; B = 8'hE8; #100;
A = 8'h3F; B = 8'hE9; #100;
A = 8'h3F; B = 8'hEA; #100;
A = 8'h3F; B = 8'hEB; #100;
A = 8'h3F; B = 8'hEC; #100;
A = 8'h3F; B = 8'hED; #100;
A = 8'h3F; B = 8'hEE; #100;
A = 8'h3F; B = 8'hEF; #100;
A = 8'h3F; B = 8'hF0; #100;
A = 8'h3F; B = 8'hF1; #100;
A = 8'h3F; B = 8'hF2; #100;
A = 8'h3F; B = 8'hF3; #100;
A = 8'h3F; B = 8'hF4; #100;
A = 8'h3F; B = 8'hF5; #100;
A = 8'h3F; B = 8'hF6; #100;
A = 8'h3F; B = 8'hF7; #100;
A = 8'h3F; B = 8'hF8; #100;
A = 8'h3F; B = 8'hF9; #100;
A = 8'h3F; B = 8'hFA; #100;
A = 8'h3F; B = 8'hFB; #100;
A = 8'h3F; B = 8'hFC; #100;
A = 8'h3F; B = 8'hFD; #100;
A = 8'h3F; B = 8'hFE; #100;
A = 8'h3F; B = 8'hFF; #100;
A = 8'h40; B = 8'h0; #100;
A = 8'h40; B = 8'h1; #100;
A = 8'h40; B = 8'h2; #100;
A = 8'h40; B = 8'h3; #100;
A = 8'h40; B = 8'h4; #100;
A = 8'h40; B = 8'h5; #100;
A = 8'h40; B = 8'h6; #100;
A = 8'h40; B = 8'h7; #100;
A = 8'h40; B = 8'h8; #100;
A = 8'h40; B = 8'h9; #100;
A = 8'h40; B = 8'hA; #100;
A = 8'h40; B = 8'hB; #100;
A = 8'h40; B = 8'hC; #100;
A = 8'h40; B = 8'hD; #100;
A = 8'h40; B = 8'hE; #100;
A = 8'h40; B = 8'hF; #100;
A = 8'h40; B = 8'h10; #100;
A = 8'h40; B = 8'h11; #100;
A = 8'h40; B = 8'h12; #100;
A = 8'h40; B = 8'h13; #100;
A = 8'h40; B = 8'h14; #100;
A = 8'h40; B = 8'h15; #100;
A = 8'h40; B = 8'h16; #100;
A = 8'h40; B = 8'h17; #100;
A = 8'h40; B = 8'h18; #100;
A = 8'h40; B = 8'h19; #100;
A = 8'h40; B = 8'h1A; #100;
A = 8'h40; B = 8'h1B; #100;
A = 8'h40; B = 8'h1C; #100;
A = 8'h40; B = 8'h1D; #100;
A = 8'h40; B = 8'h1E; #100;
A = 8'h40; B = 8'h1F; #100;
A = 8'h40; B = 8'h20; #100;
A = 8'h40; B = 8'h21; #100;
A = 8'h40; B = 8'h22; #100;
A = 8'h40; B = 8'h23; #100;
A = 8'h40; B = 8'h24; #100;
A = 8'h40; B = 8'h25; #100;
A = 8'h40; B = 8'h26; #100;
A = 8'h40; B = 8'h27; #100;
A = 8'h40; B = 8'h28; #100;
A = 8'h40; B = 8'h29; #100;
A = 8'h40; B = 8'h2A; #100;
A = 8'h40; B = 8'h2B; #100;
A = 8'h40; B = 8'h2C; #100;
A = 8'h40; B = 8'h2D; #100;
A = 8'h40; B = 8'h2E; #100;
A = 8'h40; B = 8'h2F; #100;
A = 8'h40; B = 8'h30; #100;
A = 8'h40; B = 8'h31; #100;
A = 8'h40; B = 8'h32; #100;
A = 8'h40; B = 8'h33; #100;
A = 8'h40; B = 8'h34; #100;
A = 8'h40; B = 8'h35; #100;
A = 8'h40; B = 8'h36; #100;
A = 8'h40; B = 8'h37; #100;
A = 8'h40; B = 8'h38; #100;
A = 8'h40; B = 8'h39; #100;
A = 8'h40; B = 8'h3A; #100;
A = 8'h40; B = 8'h3B; #100;
A = 8'h40; B = 8'h3C; #100;
A = 8'h40; B = 8'h3D; #100;
A = 8'h40; B = 8'h3E; #100;
A = 8'h40; B = 8'h3F; #100;
A = 8'h40; B = 8'h40; #100;
A = 8'h40; B = 8'h41; #100;
A = 8'h40; B = 8'h42; #100;
A = 8'h40; B = 8'h43; #100;
A = 8'h40; B = 8'h44; #100;
A = 8'h40; B = 8'h45; #100;
A = 8'h40; B = 8'h46; #100;
A = 8'h40; B = 8'h47; #100;
A = 8'h40; B = 8'h48; #100;
A = 8'h40; B = 8'h49; #100;
A = 8'h40; B = 8'h4A; #100;
A = 8'h40; B = 8'h4B; #100;
A = 8'h40; B = 8'h4C; #100;
A = 8'h40; B = 8'h4D; #100;
A = 8'h40; B = 8'h4E; #100;
A = 8'h40; B = 8'h4F; #100;
A = 8'h40; B = 8'h50; #100;
A = 8'h40; B = 8'h51; #100;
A = 8'h40; B = 8'h52; #100;
A = 8'h40; B = 8'h53; #100;
A = 8'h40; B = 8'h54; #100;
A = 8'h40; B = 8'h55; #100;
A = 8'h40; B = 8'h56; #100;
A = 8'h40; B = 8'h57; #100;
A = 8'h40; B = 8'h58; #100;
A = 8'h40; B = 8'h59; #100;
A = 8'h40; B = 8'h5A; #100;
A = 8'h40; B = 8'h5B; #100;
A = 8'h40; B = 8'h5C; #100;
A = 8'h40; B = 8'h5D; #100;
A = 8'h40; B = 8'h5E; #100;
A = 8'h40; B = 8'h5F; #100;
A = 8'h40; B = 8'h60; #100;
A = 8'h40; B = 8'h61; #100;
A = 8'h40; B = 8'h62; #100;
A = 8'h40; B = 8'h63; #100;
A = 8'h40; B = 8'h64; #100;
A = 8'h40; B = 8'h65; #100;
A = 8'h40; B = 8'h66; #100;
A = 8'h40; B = 8'h67; #100;
A = 8'h40; B = 8'h68; #100;
A = 8'h40; B = 8'h69; #100;
A = 8'h40; B = 8'h6A; #100;
A = 8'h40; B = 8'h6B; #100;
A = 8'h40; B = 8'h6C; #100;
A = 8'h40; B = 8'h6D; #100;
A = 8'h40; B = 8'h6E; #100;
A = 8'h40; B = 8'h6F; #100;
A = 8'h40; B = 8'h70; #100;
A = 8'h40; B = 8'h71; #100;
A = 8'h40; B = 8'h72; #100;
A = 8'h40; B = 8'h73; #100;
A = 8'h40; B = 8'h74; #100;
A = 8'h40; B = 8'h75; #100;
A = 8'h40; B = 8'h76; #100;
A = 8'h40; B = 8'h77; #100;
A = 8'h40; B = 8'h78; #100;
A = 8'h40; B = 8'h79; #100;
A = 8'h40; B = 8'h7A; #100;
A = 8'h40; B = 8'h7B; #100;
A = 8'h40; B = 8'h7C; #100;
A = 8'h40; B = 8'h7D; #100;
A = 8'h40; B = 8'h7E; #100;
A = 8'h40; B = 8'h7F; #100;
A = 8'h40; B = 8'h80; #100;
A = 8'h40; B = 8'h81; #100;
A = 8'h40; B = 8'h82; #100;
A = 8'h40; B = 8'h83; #100;
A = 8'h40; B = 8'h84; #100;
A = 8'h40; B = 8'h85; #100;
A = 8'h40; B = 8'h86; #100;
A = 8'h40; B = 8'h87; #100;
A = 8'h40; B = 8'h88; #100;
A = 8'h40; B = 8'h89; #100;
A = 8'h40; B = 8'h8A; #100;
A = 8'h40; B = 8'h8B; #100;
A = 8'h40; B = 8'h8C; #100;
A = 8'h40; B = 8'h8D; #100;
A = 8'h40; B = 8'h8E; #100;
A = 8'h40; B = 8'h8F; #100;
A = 8'h40; B = 8'h90; #100;
A = 8'h40; B = 8'h91; #100;
A = 8'h40; B = 8'h92; #100;
A = 8'h40; B = 8'h93; #100;
A = 8'h40; B = 8'h94; #100;
A = 8'h40; B = 8'h95; #100;
A = 8'h40; B = 8'h96; #100;
A = 8'h40; B = 8'h97; #100;
A = 8'h40; B = 8'h98; #100;
A = 8'h40; B = 8'h99; #100;
A = 8'h40; B = 8'h9A; #100;
A = 8'h40; B = 8'h9B; #100;
A = 8'h40; B = 8'h9C; #100;
A = 8'h40; B = 8'h9D; #100;
A = 8'h40; B = 8'h9E; #100;
A = 8'h40; B = 8'h9F; #100;
A = 8'h40; B = 8'hA0; #100;
A = 8'h40; B = 8'hA1; #100;
A = 8'h40; B = 8'hA2; #100;
A = 8'h40; B = 8'hA3; #100;
A = 8'h40; B = 8'hA4; #100;
A = 8'h40; B = 8'hA5; #100;
A = 8'h40; B = 8'hA6; #100;
A = 8'h40; B = 8'hA7; #100;
A = 8'h40; B = 8'hA8; #100;
A = 8'h40; B = 8'hA9; #100;
A = 8'h40; B = 8'hAA; #100;
A = 8'h40; B = 8'hAB; #100;
A = 8'h40; B = 8'hAC; #100;
A = 8'h40; B = 8'hAD; #100;
A = 8'h40; B = 8'hAE; #100;
A = 8'h40; B = 8'hAF; #100;
A = 8'h40; B = 8'hB0; #100;
A = 8'h40; B = 8'hB1; #100;
A = 8'h40; B = 8'hB2; #100;
A = 8'h40; B = 8'hB3; #100;
A = 8'h40; B = 8'hB4; #100;
A = 8'h40; B = 8'hB5; #100;
A = 8'h40; B = 8'hB6; #100;
A = 8'h40; B = 8'hB7; #100;
A = 8'h40; B = 8'hB8; #100;
A = 8'h40; B = 8'hB9; #100;
A = 8'h40; B = 8'hBA; #100;
A = 8'h40; B = 8'hBB; #100;
A = 8'h40; B = 8'hBC; #100;
A = 8'h40; B = 8'hBD; #100;
A = 8'h40; B = 8'hBE; #100;
A = 8'h40; B = 8'hBF; #100;
A = 8'h40; B = 8'hC0; #100;
A = 8'h40; B = 8'hC1; #100;
A = 8'h40; B = 8'hC2; #100;
A = 8'h40; B = 8'hC3; #100;
A = 8'h40; B = 8'hC4; #100;
A = 8'h40; B = 8'hC5; #100;
A = 8'h40; B = 8'hC6; #100;
A = 8'h40; B = 8'hC7; #100;
A = 8'h40; B = 8'hC8; #100;
A = 8'h40; B = 8'hC9; #100;
A = 8'h40; B = 8'hCA; #100;
A = 8'h40; B = 8'hCB; #100;
A = 8'h40; B = 8'hCC; #100;
A = 8'h40; B = 8'hCD; #100;
A = 8'h40; B = 8'hCE; #100;
A = 8'h40; B = 8'hCF; #100;
A = 8'h40; B = 8'hD0; #100;
A = 8'h40; B = 8'hD1; #100;
A = 8'h40; B = 8'hD2; #100;
A = 8'h40; B = 8'hD3; #100;
A = 8'h40; B = 8'hD4; #100;
A = 8'h40; B = 8'hD5; #100;
A = 8'h40; B = 8'hD6; #100;
A = 8'h40; B = 8'hD7; #100;
A = 8'h40; B = 8'hD8; #100;
A = 8'h40; B = 8'hD9; #100;
A = 8'h40; B = 8'hDA; #100;
A = 8'h40; B = 8'hDB; #100;
A = 8'h40; B = 8'hDC; #100;
A = 8'h40; B = 8'hDD; #100;
A = 8'h40; B = 8'hDE; #100;
A = 8'h40; B = 8'hDF; #100;
A = 8'h40; B = 8'hE0; #100;
A = 8'h40; B = 8'hE1; #100;
A = 8'h40; B = 8'hE2; #100;
A = 8'h40; B = 8'hE3; #100;
A = 8'h40; B = 8'hE4; #100;
A = 8'h40; B = 8'hE5; #100;
A = 8'h40; B = 8'hE6; #100;
A = 8'h40; B = 8'hE7; #100;
A = 8'h40; B = 8'hE8; #100;
A = 8'h40; B = 8'hE9; #100;
A = 8'h40; B = 8'hEA; #100;
A = 8'h40; B = 8'hEB; #100;
A = 8'h40; B = 8'hEC; #100;
A = 8'h40; B = 8'hED; #100;
A = 8'h40; B = 8'hEE; #100;
A = 8'h40; B = 8'hEF; #100;
A = 8'h40; B = 8'hF0; #100;
A = 8'h40; B = 8'hF1; #100;
A = 8'h40; B = 8'hF2; #100;
A = 8'h40; B = 8'hF3; #100;
A = 8'h40; B = 8'hF4; #100;
A = 8'h40; B = 8'hF5; #100;
A = 8'h40; B = 8'hF6; #100;
A = 8'h40; B = 8'hF7; #100;
A = 8'h40; B = 8'hF8; #100;
A = 8'h40; B = 8'hF9; #100;
A = 8'h40; B = 8'hFA; #100;
A = 8'h40; B = 8'hFB; #100;
A = 8'h40; B = 8'hFC; #100;
A = 8'h40; B = 8'hFD; #100;
A = 8'h40; B = 8'hFE; #100;
A = 8'h40; B = 8'hFF; #100;
A = 8'h41; B = 8'h0; #100;
A = 8'h41; B = 8'h1; #100;
A = 8'h41; B = 8'h2; #100;
A = 8'h41; B = 8'h3; #100;
A = 8'h41; B = 8'h4; #100;
A = 8'h41; B = 8'h5; #100;
A = 8'h41; B = 8'h6; #100;
A = 8'h41; B = 8'h7; #100;
A = 8'h41; B = 8'h8; #100;
A = 8'h41; B = 8'h9; #100;
A = 8'h41; B = 8'hA; #100;
A = 8'h41; B = 8'hB; #100;
A = 8'h41; B = 8'hC; #100;
A = 8'h41; B = 8'hD; #100;
A = 8'h41; B = 8'hE; #100;
A = 8'h41; B = 8'hF; #100;
A = 8'h41; B = 8'h10; #100;
A = 8'h41; B = 8'h11; #100;
A = 8'h41; B = 8'h12; #100;
A = 8'h41; B = 8'h13; #100;
A = 8'h41; B = 8'h14; #100;
A = 8'h41; B = 8'h15; #100;
A = 8'h41; B = 8'h16; #100;
A = 8'h41; B = 8'h17; #100;
A = 8'h41; B = 8'h18; #100;
A = 8'h41; B = 8'h19; #100;
A = 8'h41; B = 8'h1A; #100;
A = 8'h41; B = 8'h1B; #100;
A = 8'h41; B = 8'h1C; #100;
A = 8'h41; B = 8'h1D; #100;
A = 8'h41; B = 8'h1E; #100;
A = 8'h41; B = 8'h1F; #100;
A = 8'h41; B = 8'h20; #100;
A = 8'h41; B = 8'h21; #100;
A = 8'h41; B = 8'h22; #100;
A = 8'h41; B = 8'h23; #100;
A = 8'h41; B = 8'h24; #100;
A = 8'h41; B = 8'h25; #100;
A = 8'h41; B = 8'h26; #100;
A = 8'h41; B = 8'h27; #100;
A = 8'h41; B = 8'h28; #100;
A = 8'h41; B = 8'h29; #100;
A = 8'h41; B = 8'h2A; #100;
A = 8'h41; B = 8'h2B; #100;
A = 8'h41; B = 8'h2C; #100;
A = 8'h41; B = 8'h2D; #100;
A = 8'h41; B = 8'h2E; #100;
A = 8'h41; B = 8'h2F; #100;
A = 8'h41; B = 8'h30; #100;
A = 8'h41; B = 8'h31; #100;
A = 8'h41; B = 8'h32; #100;
A = 8'h41; B = 8'h33; #100;
A = 8'h41; B = 8'h34; #100;
A = 8'h41; B = 8'h35; #100;
A = 8'h41; B = 8'h36; #100;
A = 8'h41; B = 8'h37; #100;
A = 8'h41; B = 8'h38; #100;
A = 8'h41; B = 8'h39; #100;
A = 8'h41; B = 8'h3A; #100;
A = 8'h41; B = 8'h3B; #100;
A = 8'h41; B = 8'h3C; #100;
A = 8'h41; B = 8'h3D; #100;
A = 8'h41; B = 8'h3E; #100;
A = 8'h41; B = 8'h3F; #100;
A = 8'h41; B = 8'h40; #100;
A = 8'h41; B = 8'h41; #100;
A = 8'h41; B = 8'h42; #100;
A = 8'h41; B = 8'h43; #100;
A = 8'h41; B = 8'h44; #100;
A = 8'h41; B = 8'h45; #100;
A = 8'h41; B = 8'h46; #100;
A = 8'h41; B = 8'h47; #100;
A = 8'h41; B = 8'h48; #100;
A = 8'h41; B = 8'h49; #100;
A = 8'h41; B = 8'h4A; #100;
A = 8'h41; B = 8'h4B; #100;
A = 8'h41; B = 8'h4C; #100;
A = 8'h41; B = 8'h4D; #100;
A = 8'h41; B = 8'h4E; #100;
A = 8'h41; B = 8'h4F; #100;
A = 8'h41; B = 8'h50; #100;
A = 8'h41; B = 8'h51; #100;
A = 8'h41; B = 8'h52; #100;
A = 8'h41; B = 8'h53; #100;
A = 8'h41; B = 8'h54; #100;
A = 8'h41; B = 8'h55; #100;
A = 8'h41; B = 8'h56; #100;
A = 8'h41; B = 8'h57; #100;
A = 8'h41; B = 8'h58; #100;
A = 8'h41; B = 8'h59; #100;
A = 8'h41; B = 8'h5A; #100;
A = 8'h41; B = 8'h5B; #100;
A = 8'h41; B = 8'h5C; #100;
A = 8'h41; B = 8'h5D; #100;
A = 8'h41; B = 8'h5E; #100;
A = 8'h41; B = 8'h5F; #100;
A = 8'h41; B = 8'h60; #100;
A = 8'h41; B = 8'h61; #100;
A = 8'h41; B = 8'h62; #100;
A = 8'h41; B = 8'h63; #100;
A = 8'h41; B = 8'h64; #100;
A = 8'h41; B = 8'h65; #100;
A = 8'h41; B = 8'h66; #100;
A = 8'h41; B = 8'h67; #100;
A = 8'h41; B = 8'h68; #100;
A = 8'h41; B = 8'h69; #100;
A = 8'h41; B = 8'h6A; #100;
A = 8'h41; B = 8'h6B; #100;
A = 8'h41; B = 8'h6C; #100;
A = 8'h41; B = 8'h6D; #100;
A = 8'h41; B = 8'h6E; #100;
A = 8'h41; B = 8'h6F; #100;
A = 8'h41; B = 8'h70; #100;
A = 8'h41; B = 8'h71; #100;
A = 8'h41; B = 8'h72; #100;
A = 8'h41; B = 8'h73; #100;
A = 8'h41; B = 8'h74; #100;
A = 8'h41; B = 8'h75; #100;
A = 8'h41; B = 8'h76; #100;
A = 8'h41; B = 8'h77; #100;
A = 8'h41; B = 8'h78; #100;
A = 8'h41; B = 8'h79; #100;
A = 8'h41; B = 8'h7A; #100;
A = 8'h41; B = 8'h7B; #100;
A = 8'h41; B = 8'h7C; #100;
A = 8'h41; B = 8'h7D; #100;
A = 8'h41; B = 8'h7E; #100;
A = 8'h41; B = 8'h7F; #100;
A = 8'h41; B = 8'h80; #100;
A = 8'h41; B = 8'h81; #100;
A = 8'h41; B = 8'h82; #100;
A = 8'h41; B = 8'h83; #100;
A = 8'h41; B = 8'h84; #100;
A = 8'h41; B = 8'h85; #100;
A = 8'h41; B = 8'h86; #100;
A = 8'h41; B = 8'h87; #100;
A = 8'h41; B = 8'h88; #100;
A = 8'h41; B = 8'h89; #100;
A = 8'h41; B = 8'h8A; #100;
A = 8'h41; B = 8'h8B; #100;
A = 8'h41; B = 8'h8C; #100;
A = 8'h41; B = 8'h8D; #100;
A = 8'h41; B = 8'h8E; #100;
A = 8'h41; B = 8'h8F; #100;
A = 8'h41; B = 8'h90; #100;
A = 8'h41; B = 8'h91; #100;
A = 8'h41; B = 8'h92; #100;
A = 8'h41; B = 8'h93; #100;
A = 8'h41; B = 8'h94; #100;
A = 8'h41; B = 8'h95; #100;
A = 8'h41; B = 8'h96; #100;
A = 8'h41; B = 8'h97; #100;
A = 8'h41; B = 8'h98; #100;
A = 8'h41; B = 8'h99; #100;
A = 8'h41; B = 8'h9A; #100;
A = 8'h41; B = 8'h9B; #100;
A = 8'h41; B = 8'h9C; #100;
A = 8'h41; B = 8'h9D; #100;
A = 8'h41; B = 8'h9E; #100;
A = 8'h41; B = 8'h9F; #100;
A = 8'h41; B = 8'hA0; #100;
A = 8'h41; B = 8'hA1; #100;
A = 8'h41; B = 8'hA2; #100;
A = 8'h41; B = 8'hA3; #100;
A = 8'h41; B = 8'hA4; #100;
A = 8'h41; B = 8'hA5; #100;
A = 8'h41; B = 8'hA6; #100;
A = 8'h41; B = 8'hA7; #100;
A = 8'h41; B = 8'hA8; #100;
A = 8'h41; B = 8'hA9; #100;
A = 8'h41; B = 8'hAA; #100;
A = 8'h41; B = 8'hAB; #100;
A = 8'h41; B = 8'hAC; #100;
A = 8'h41; B = 8'hAD; #100;
A = 8'h41; B = 8'hAE; #100;
A = 8'h41; B = 8'hAF; #100;
A = 8'h41; B = 8'hB0; #100;
A = 8'h41; B = 8'hB1; #100;
A = 8'h41; B = 8'hB2; #100;
A = 8'h41; B = 8'hB3; #100;
A = 8'h41; B = 8'hB4; #100;
A = 8'h41; B = 8'hB5; #100;
A = 8'h41; B = 8'hB6; #100;
A = 8'h41; B = 8'hB7; #100;
A = 8'h41; B = 8'hB8; #100;
A = 8'h41; B = 8'hB9; #100;
A = 8'h41; B = 8'hBA; #100;
A = 8'h41; B = 8'hBB; #100;
A = 8'h41; B = 8'hBC; #100;
A = 8'h41; B = 8'hBD; #100;
A = 8'h41; B = 8'hBE; #100;
A = 8'h41; B = 8'hBF; #100;
A = 8'h41; B = 8'hC0; #100;
A = 8'h41; B = 8'hC1; #100;
A = 8'h41; B = 8'hC2; #100;
A = 8'h41; B = 8'hC3; #100;
A = 8'h41; B = 8'hC4; #100;
A = 8'h41; B = 8'hC5; #100;
A = 8'h41; B = 8'hC6; #100;
A = 8'h41; B = 8'hC7; #100;
A = 8'h41; B = 8'hC8; #100;
A = 8'h41; B = 8'hC9; #100;
A = 8'h41; B = 8'hCA; #100;
A = 8'h41; B = 8'hCB; #100;
A = 8'h41; B = 8'hCC; #100;
A = 8'h41; B = 8'hCD; #100;
A = 8'h41; B = 8'hCE; #100;
A = 8'h41; B = 8'hCF; #100;
A = 8'h41; B = 8'hD0; #100;
A = 8'h41; B = 8'hD1; #100;
A = 8'h41; B = 8'hD2; #100;
A = 8'h41; B = 8'hD3; #100;
A = 8'h41; B = 8'hD4; #100;
A = 8'h41; B = 8'hD5; #100;
A = 8'h41; B = 8'hD6; #100;
A = 8'h41; B = 8'hD7; #100;
A = 8'h41; B = 8'hD8; #100;
A = 8'h41; B = 8'hD9; #100;
A = 8'h41; B = 8'hDA; #100;
A = 8'h41; B = 8'hDB; #100;
A = 8'h41; B = 8'hDC; #100;
A = 8'h41; B = 8'hDD; #100;
A = 8'h41; B = 8'hDE; #100;
A = 8'h41; B = 8'hDF; #100;
A = 8'h41; B = 8'hE0; #100;
A = 8'h41; B = 8'hE1; #100;
A = 8'h41; B = 8'hE2; #100;
A = 8'h41; B = 8'hE3; #100;
A = 8'h41; B = 8'hE4; #100;
A = 8'h41; B = 8'hE5; #100;
A = 8'h41; B = 8'hE6; #100;
A = 8'h41; B = 8'hE7; #100;
A = 8'h41; B = 8'hE8; #100;
A = 8'h41; B = 8'hE9; #100;
A = 8'h41; B = 8'hEA; #100;
A = 8'h41; B = 8'hEB; #100;
A = 8'h41; B = 8'hEC; #100;
A = 8'h41; B = 8'hED; #100;
A = 8'h41; B = 8'hEE; #100;
A = 8'h41; B = 8'hEF; #100;
A = 8'h41; B = 8'hF0; #100;
A = 8'h41; B = 8'hF1; #100;
A = 8'h41; B = 8'hF2; #100;
A = 8'h41; B = 8'hF3; #100;
A = 8'h41; B = 8'hF4; #100;
A = 8'h41; B = 8'hF5; #100;
A = 8'h41; B = 8'hF6; #100;
A = 8'h41; B = 8'hF7; #100;
A = 8'h41; B = 8'hF8; #100;
A = 8'h41; B = 8'hF9; #100;
A = 8'h41; B = 8'hFA; #100;
A = 8'h41; B = 8'hFB; #100;
A = 8'h41; B = 8'hFC; #100;
A = 8'h41; B = 8'hFD; #100;
A = 8'h41; B = 8'hFE; #100;
A = 8'h41; B = 8'hFF; #100;
A = 8'h42; B = 8'h0; #100;
A = 8'h42; B = 8'h1; #100;
A = 8'h42; B = 8'h2; #100;
A = 8'h42; B = 8'h3; #100;
A = 8'h42; B = 8'h4; #100;
A = 8'h42; B = 8'h5; #100;
A = 8'h42; B = 8'h6; #100;
A = 8'h42; B = 8'h7; #100;
A = 8'h42; B = 8'h8; #100;
A = 8'h42; B = 8'h9; #100;
A = 8'h42; B = 8'hA; #100;
A = 8'h42; B = 8'hB; #100;
A = 8'h42; B = 8'hC; #100;
A = 8'h42; B = 8'hD; #100;
A = 8'h42; B = 8'hE; #100;
A = 8'h42; B = 8'hF; #100;
A = 8'h42; B = 8'h10; #100;
A = 8'h42; B = 8'h11; #100;
A = 8'h42; B = 8'h12; #100;
A = 8'h42; B = 8'h13; #100;
A = 8'h42; B = 8'h14; #100;
A = 8'h42; B = 8'h15; #100;
A = 8'h42; B = 8'h16; #100;
A = 8'h42; B = 8'h17; #100;
A = 8'h42; B = 8'h18; #100;
A = 8'h42; B = 8'h19; #100;
A = 8'h42; B = 8'h1A; #100;
A = 8'h42; B = 8'h1B; #100;
A = 8'h42; B = 8'h1C; #100;
A = 8'h42; B = 8'h1D; #100;
A = 8'h42; B = 8'h1E; #100;
A = 8'h42; B = 8'h1F; #100;
A = 8'h42; B = 8'h20; #100;
A = 8'h42; B = 8'h21; #100;
A = 8'h42; B = 8'h22; #100;
A = 8'h42; B = 8'h23; #100;
A = 8'h42; B = 8'h24; #100;
A = 8'h42; B = 8'h25; #100;
A = 8'h42; B = 8'h26; #100;
A = 8'h42; B = 8'h27; #100;
A = 8'h42; B = 8'h28; #100;
A = 8'h42; B = 8'h29; #100;
A = 8'h42; B = 8'h2A; #100;
A = 8'h42; B = 8'h2B; #100;
A = 8'h42; B = 8'h2C; #100;
A = 8'h42; B = 8'h2D; #100;
A = 8'h42; B = 8'h2E; #100;
A = 8'h42; B = 8'h2F; #100;
A = 8'h42; B = 8'h30; #100;
A = 8'h42; B = 8'h31; #100;
A = 8'h42; B = 8'h32; #100;
A = 8'h42; B = 8'h33; #100;
A = 8'h42; B = 8'h34; #100;
A = 8'h42; B = 8'h35; #100;
A = 8'h42; B = 8'h36; #100;
A = 8'h42; B = 8'h37; #100;
A = 8'h42; B = 8'h38; #100;
A = 8'h42; B = 8'h39; #100;
A = 8'h42; B = 8'h3A; #100;
A = 8'h42; B = 8'h3B; #100;
A = 8'h42; B = 8'h3C; #100;
A = 8'h42; B = 8'h3D; #100;
A = 8'h42; B = 8'h3E; #100;
A = 8'h42; B = 8'h3F; #100;
A = 8'h42; B = 8'h40; #100;
A = 8'h42; B = 8'h41; #100;
A = 8'h42; B = 8'h42; #100;
A = 8'h42; B = 8'h43; #100;
A = 8'h42; B = 8'h44; #100;
A = 8'h42; B = 8'h45; #100;
A = 8'h42; B = 8'h46; #100;
A = 8'h42; B = 8'h47; #100;
A = 8'h42; B = 8'h48; #100;
A = 8'h42; B = 8'h49; #100;
A = 8'h42; B = 8'h4A; #100;
A = 8'h42; B = 8'h4B; #100;
A = 8'h42; B = 8'h4C; #100;
A = 8'h42; B = 8'h4D; #100;
A = 8'h42; B = 8'h4E; #100;
A = 8'h42; B = 8'h4F; #100;
A = 8'h42; B = 8'h50; #100;
A = 8'h42; B = 8'h51; #100;
A = 8'h42; B = 8'h52; #100;
A = 8'h42; B = 8'h53; #100;
A = 8'h42; B = 8'h54; #100;
A = 8'h42; B = 8'h55; #100;
A = 8'h42; B = 8'h56; #100;
A = 8'h42; B = 8'h57; #100;
A = 8'h42; B = 8'h58; #100;
A = 8'h42; B = 8'h59; #100;
A = 8'h42; B = 8'h5A; #100;
A = 8'h42; B = 8'h5B; #100;
A = 8'h42; B = 8'h5C; #100;
A = 8'h42; B = 8'h5D; #100;
A = 8'h42; B = 8'h5E; #100;
A = 8'h42; B = 8'h5F; #100;
A = 8'h42; B = 8'h60; #100;
A = 8'h42; B = 8'h61; #100;
A = 8'h42; B = 8'h62; #100;
A = 8'h42; B = 8'h63; #100;
A = 8'h42; B = 8'h64; #100;
A = 8'h42; B = 8'h65; #100;
A = 8'h42; B = 8'h66; #100;
A = 8'h42; B = 8'h67; #100;
A = 8'h42; B = 8'h68; #100;
A = 8'h42; B = 8'h69; #100;
A = 8'h42; B = 8'h6A; #100;
A = 8'h42; B = 8'h6B; #100;
A = 8'h42; B = 8'h6C; #100;
A = 8'h42; B = 8'h6D; #100;
A = 8'h42; B = 8'h6E; #100;
A = 8'h42; B = 8'h6F; #100;
A = 8'h42; B = 8'h70; #100;
A = 8'h42; B = 8'h71; #100;
A = 8'h42; B = 8'h72; #100;
A = 8'h42; B = 8'h73; #100;
A = 8'h42; B = 8'h74; #100;
A = 8'h42; B = 8'h75; #100;
A = 8'h42; B = 8'h76; #100;
A = 8'h42; B = 8'h77; #100;
A = 8'h42; B = 8'h78; #100;
A = 8'h42; B = 8'h79; #100;
A = 8'h42; B = 8'h7A; #100;
A = 8'h42; B = 8'h7B; #100;
A = 8'h42; B = 8'h7C; #100;
A = 8'h42; B = 8'h7D; #100;
A = 8'h42; B = 8'h7E; #100;
A = 8'h42; B = 8'h7F; #100;
A = 8'h42; B = 8'h80; #100;
A = 8'h42; B = 8'h81; #100;
A = 8'h42; B = 8'h82; #100;
A = 8'h42; B = 8'h83; #100;
A = 8'h42; B = 8'h84; #100;
A = 8'h42; B = 8'h85; #100;
A = 8'h42; B = 8'h86; #100;
A = 8'h42; B = 8'h87; #100;
A = 8'h42; B = 8'h88; #100;
A = 8'h42; B = 8'h89; #100;
A = 8'h42; B = 8'h8A; #100;
A = 8'h42; B = 8'h8B; #100;
A = 8'h42; B = 8'h8C; #100;
A = 8'h42; B = 8'h8D; #100;
A = 8'h42; B = 8'h8E; #100;
A = 8'h42; B = 8'h8F; #100;
A = 8'h42; B = 8'h90; #100;
A = 8'h42; B = 8'h91; #100;
A = 8'h42; B = 8'h92; #100;
A = 8'h42; B = 8'h93; #100;
A = 8'h42; B = 8'h94; #100;
A = 8'h42; B = 8'h95; #100;
A = 8'h42; B = 8'h96; #100;
A = 8'h42; B = 8'h97; #100;
A = 8'h42; B = 8'h98; #100;
A = 8'h42; B = 8'h99; #100;
A = 8'h42; B = 8'h9A; #100;
A = 8'h42; B = 8'h9B; #100;
A = 8'h42; B = 8'h9C; #100;
A = 8'h42; B = 8'h9D; #100;
A = 8'h42; B = 8'h9E; #100;
A = 8'h42; B = 8'h9F; #100;
A = 8'h42; B = 8'hA0; #100;
A = 8'h42; B = 8'hA1; #100;
A = 8'h42; B = 8'hA2; #100;
A = 8'h42; B = 8'hA3; #100;
A = 8'h42; B = 8'hA4; #100;
A = 8'h42; B = 8'hA5; #100;
A = 8'h42; B = 8'hA6; #100;
A = 8'h42; B = 8'hA7; #100;
A = 8'h42; B = 8'hA8; #100;
A = 8'h42; B = 8'hA9; #100;
A = 8'h42; B = 8'hAA; #100;
A = 8'h42; B = 8'hAB; #100;
A = 8'h42; B = 8'hAC; #100;
A = 8'h42; B = 8'hAD; #100;
A = 8'h42; B = 8'hAE; #100;
A = 8'h42; B = 8'hAF; #100;
A = 8'h42; B = 8'hB0; #100;
A = 8'h42; B = 8'hB1; #100;
A = 8'h42; B = 8'hB2; #100;
A = 8'h42; B = 8'hB3; #100;
A = 8'h42; B = 8'hB4; #100;
A = 8'h42; B = 8'hB5; #100;
A = 8'h42; B = 8'hB6; #100;
A = 8'h42; B = 8'hB7; #100;
A = 8'h42; B = 8'hB8; #100;
A = 8'h42; B = 8'hB9; #100;
A = 8'h42; B = 8'hBA; #100;
A = 8'h42; B = 8'hBB; #100;
A = 8'h42; B = 8'hBC; #100;
A = 8'h42; B = 8'hBD; #100;
A = 8'h42; B = 8'hBE; #100;
A = 8'h42; B = 8'hBF; #100;
A = 8'h42; B = 8'hC0; #100;
A = 8'h42; B = 8'hC1; #100;
A = 8'h42; B = 8'hC2; #100;
A = 8'h42; B = 8'hC3; #100;
A = 8'h42; B = 8'hC4; #100;
A = 8'h42; B = 8'hC5; #100;
A = 8'h42; B = 8'hC6; #100;
A = 8'h42; B = 8'hC7; #100;
A = 8'h42; B = 8'hC8; #100;
A = 8'h42; B = 8'hC9; #100;
A = 8'h42; B = 8'hCA; #100;
A = 8'h42; B = 8'hCB; #100;
A = 8'h42; B = 8'hCC; #100;
A = 8'h42; B = 8'hCD; #100;
A = 8'h42; B = 8'hCE; #100;
A = 8'h42; B = 8'hCF; #100;
A = 8'h42; B = 8'hD0; #100;
A = 8'h42; B = 8'hD1; #100;
A = 8'h42; B = 8'hD2; #100;
A = 8'h42; B = 8'hD3; #100;
A = 8'h42; B = 8'hD4; #100;
A = 8'h42; B = 8'hD5; #100;
A = 8'h42; B = 8'hD6; #100;
A = 8'h42; B = 8'hD7; #100;
A = 8'h42; B = 8'hD8; #100;
A = 8'h42; B = 8'hD9; #100;
A = 8'h42; B = 8'hDA; #100;
A = 8'h42; B = 8'hDB; #100;
A = 8'h42; B = 8'hDC; #100;
A = 8'h42; B = 8'hDD; #100;
A = 8'h42; B = 8'hDE; #100;
A = 8'h42; B = 8'hDF; #100;
A = 8'h42; B = 8'hE0; #100;
A = 8'h42; B = 8'hE1; #100;
A = 8'h42; B = 8'hE2; #100;
A = 8'h42; B = 8'hE3; #100;
A = 8'h42; B = 8'hE4; #100;
A = 8'h42; B = 8'hE5; #100;
A = 8'h42; B = 8'hE6; #100;
A = 8'h42; B = 8'hE7; #100;
A = 8'h42; B = 8'hE8; #100;
A = 8'h42; B = 8'hE9; #100;
A = 8'h42; B = 8'hEA; #100;
A = 8'h42; B = 8'hEB; #100;
A = 8'h42; B = 8'hEC; #100;
A = 8'h42; B = 8'hED; #100;
A = 8'h42; B = 8'hEE; #100;
A = 8'h42; B = 8'hEF; #100;
A = 8'h42; B = 8'hF0; #100;
A = 8'h42; B = 8'hF1; #100;
A = 8'h42; B = 8'hF2; #100;
A = 8'h42; B = 8'hF3; #100;
A = 8'h42; B = 8'hF4; #100;
A = 8'h42; B = 8'hF5; #100;
A = 8'h42; B = 8'hF6; #100;
A = 8'h42; B = 8'hF7; #100;
A = 8'h42; B = 8'hF8; #100;
A = 8'h42; B = 8'hF9; #100;
A = 8'h42; B = 8'hFA; #100;
A = 8'h42; B = 8'hFB; #100;
A = 8'h42; B = 8'hFC; #100;
A = 8'h42; B = 8'hFD; #100;
A = 8'h42; B = 8'hFE; #100;
A = 8'h42; B = 8'hFF; #100;
A = 8'h43; B = 8'h0; #100;
A = 8'h43; B = 8'h1; #100;
A = 8'h43; B = 8'h2; #100;
A = 8'h43; B = 8'h3; #100;
A = 8'h43; B = 8'h4; #100;
A = 8'h43; B = 8'h5; #100;
A = 8'h43; B = 8'h6; #100;
A = 8'h43; B = 8'h7; #100;
A = 8'h43; B = 8'h8; #100;
A = 8'h43; B = 8'h9; #100;
A = 8'h43; B = 8'hA; #100;
A = 8'h43; B = 8'hB; #100;
A = 8'h43; B = 8'hC; #100;
A = 8'h43; B = 8'hD; #100;
A = 8'h43; B = 8'hE; #100;
A = 8'h43; B = 8'hF; #100;
A = 8'h43; B = 8'h10; #100;
A = 8'h43; B = 8'h11; #100;
A = 8'h43; B = 8'h12; #100;
A = 8'h43; B = 8'h13; #100;
A = 8'h43; B = 8'h14; #100;
A = 8'h43; B = 8'h15; #100;
A = 8'h43; B = 8'h16; #100;
A = 8'h43; B = 8'h17; #100;
A = 8'h43; B = 8'h18; #100;
A = 8'h43; B = 8'h19; #100;
A = 8'h43; B = 8'h1A; #100;
A = 8'h43; B = 8'h1B; #100;
A = 8'h43; B = 8'h1C; #100;
A = 8'h43; B = 8'h1D; #100;
A = 8'h43; B = 8'h1E; #100;
A = 8'h43; B = 8'h1F; #100;
A = 8'h43; B = 8'h20; #100;
A = 8'h43; B = 8'h21; #100;
A = 8'h43; B = 8'h22; #100;
A = 8'h43; B = 8'h23; #100;
A = 8'h43; B = 8'h24; #100;
A = 8'h43; B = 8'h25; #100;
A = 8'h43; B = 8'h26; #100;
A = 8'h43; B = 8'h27; #100;
A = 8'h43; B = 8'h28; #100;
A = 8'h43; B = 8'h29; #100;
A = 8'h43; B = 8'h2A; #100;
A = 8'h43; B = 8'h2B; #100;
A = 8'h43; B = 8'h2C; #100;
A = 8'h43; B = 8'h2D; #100;
A = 8'h43; B = 8'h2E; #100;
A = 8'h43; B = 8'h2F; #100;
A = 8'h43; B = 8'h30; #100;
A = 8'h43; B = 8'h31; #100;
A = 8'h43; B = 8'h32; #100;
A = 8'h43; B = 8'h33; #100;
A = 8'h43; B = 8'h34; #100;
A = 8'h43; B = 8'h35; #100;
A = 8'h43; B = 8'h36; #100;
A = 8'h43; B = 8'h37; #100;
A = 8'h43; B = 8'h38; #100;
A = 8'h43; B = 8'h39; #100;
A = 8'h43; B = 8'h3A; #100;
A = 8'h43; B = 8'h3B; #100;
A = 8'h43; B = 8'h3C; #100;
A = 8'h43; B = 8'h3D; #100;
A = 8'h43; B = 8'h3E; #100;
A = 8'h43; B = 8'h3F; #100;
A = 8'h43; B = 8'h40; #100;
A = 8'h43; B = 8'h41; #100;
A = 8'h43; B = 8'h42; #100;
A = 8'h43; B = 8'h43; #100;
A = 8'h43; B = 8'h44; #100;
A = 8'h43; B = 8'h45; #100;
A = 8'h43; B = 8'h46; #100;
A = 8'h43; B = 8'h47; #100;
A = 8'h43; B = 8'h48; #100;
A = 8'h43; B = 8'h49; #100;
A = 8'h43; B = 8'h4A; #100;
A = 8'h43; B = 8'h4B; #100;
A = 8'h43; B = 8'h4C; #100;
A = 8'h43; B = 8'h4D; #100;
A = 8'h43; B = 8'h4E; #100;
A = 8'h43; B = 8'h4F; #100;
A = 8'h43; B = 8'h50; #100;
A = 8'h43; B = 8'h51; #100;
A = 8'h43; B = 8'h52; #100;
A = 8'h43; B = 8'h53; #100;
A = 8'h43; B = 8'h54; #100;
A = 8'h43; B = 8'h55; #100;
A = 8'h43; B = 8'h56; #100;
A = 8'h43; B = 8'h57; #100;
A = 8'h43; B = 8'h58; #100;
A = 8'h43; B = 8'h59; #100;
A = 8'h43; B = 8'h5A; #100;
A = 8'h43; B = 8'h5B; #100;
A = 8'h43; B = 8'h5C; #100;
A = 8'h43; B = 8'h5D; #100;
A = 8'h43; B = 8'h5E; #100;
A = 8'h43; B = 8'h5F; #100;
A = 8'h43; B = 8'h60; #100;
A = 8'h43; B = 8'h61; #100;
A = 8'h43; B = 8'h62; #100;
A = 8'h43; B = 8'h63; #100;
A = 8'h43; B = 8'h64; #100;
A = 8'h43; B = 8'h65; #100;
A = 8'h43; B = 8'h66; #100;
A = 8'h43; B = 8'h67; #100;
A = 8'h43; B = 8'h68; #100;
A = 8'h43; B = 8'h69; #100;
A = 8'h43; B = 8'h6A; #100;
A = 8'h43; B = 8'h6B; #100;
A = 8'h43; B = 8'h6C; #100;
A = 8'h43; B = 8'h6D; #100;
A = 8'h43; B = 8'h6E; #100;
A = 8'h43; B = 8'h6F; #100;
A = 8'h43; B = 8'h70; #100;
A = 8'h43; B = 8'h71; #100;
A = 8'h43; B = 8'h72; #100;
A = 8'h43; B = 8'h73; #100;
A = 8'h43; B = 8'h74; #100;
A = 8'h43; B = 8'h75; #100;
A = 8'h43; B = 8'h76; #100;
A = 8'h43; B = 8'h77; #100;
A = 8'h43; B = 8'h78; #100;
A = 8'h43; B = 8'h79; #100;
A = 8'h43; B = 8'h7A; #100;
A = 8'h43; B = 8'h7B; #100;
A = 8'h43; B = 8'h7C; #100;
A = 8'h43; B = 8'h7D; #100;
A = 8'h43; B = 8'h7E; #100;
A = 8'h43; B = 8'h7F; #100;
A = 8'h43; B = 8'h80; #100;
A = 8'h43; B = 8'h81; #100;
A = 8'h43; B = 8'h82; #100;
A = 8'h43; B = 8'h83; #100;
A = 8'h43; B = 8'h84; #100;
A = 8'h43; B = 8'h85; #100;
A = 8'h43; B = 8'h86; #100;
A = 8'h43; B = 8'h87; #100;
A = 8'h43; B = 8'h88; #100;
A = 8'h43; B = 8'h89; #100;
A = 8'h43; B = 8'h8A; #100;
A = 8'h43; B = 8'h8B; #100;
A = 8'h43; B = 8'h8C; #100;
A = 8'h43; B = 8'h8D; #100;
A = 8'h43; B = 8'h8E; #100;
A = 8'h43; B = 8'h8F; #100;
A = 8'h43; B = 8'h90; #100;
A = 8'h43; B = 8'h91; #100;
A = 8'h43; B = 8'h92; #100;
A = 8'h43; B = 8'h93; #100;
A = 8'h43; B = 8'h94; #100;
A = 8'h43; B = 8'h95; #100;
A = 8'h43; B = 8'h96; #100;
A = 8'h43; B = 8'h97; #100;
A = 8'h43; B = 8'h98; #100;
A = 8'h43; B = 8'h99; #100;
A = 8'h43; B = 8'h9A; #100;
A = 8'h43; B = 8'h9B; #100;
A = 8'h43; B = 8'h9C; #100;
A = 8'h43; B = 8'h9D; #100;
A = 8'h43; B = 8'h9E; #100;
A = 8'h43; B = 8'h9F; #100;
A = 8'h43; B = 8'hA0; #100;
A = 8'h43; B = 8'hA1; #100;
A = 8'h43; B = 8'hA2; #100;
A = 8'h43; B = 8'hA3; #100;
A = 8'h43; B = 8'hA4; #100;
A = 8'h43; B = 8'hA5; #100;
A = 8'h43; B = 8'hA6; #100;
A = 8'h43; B = 8'hA7; #100;
A = 8'h43; B = 8'hA8; #100;
A = 8'h43; B = 8'hA9; #100;
A = 8'h43; B = 8'hAA; #100;
A = 8'h43; B = 8'hAB; #100;
A = 8'h43; B = 8'hAC; #100;
A = 8'h43; B = 8'hAD; #100;
A = 8'h43; B = 8'hAE; #100;
A = 8'h43; B = 8'hAF; #100;
A = 8'h43; B = 8'hB0; #100;
A = 8'h43; B = 8'hB1; #100;
A = 8'h43; B = 8'hB2; #100;
A = 8'h43; B = 8'hB3; #100;
A = 8'h43; B = 8'hB4; #100;
A = 8'h43; B = 8'hB5; #100;
A = 8'h43; B = 8'hB6; #100;
A = 8'h43; B = 8'hB7; #100;
A = 8'h43; B = 8'hB8; #100;
A = 8'h43; B = 8'hB9; #100;
A = 8'h43; B = 8'hBA; #100;
A = 8'h43; B = 8'hBB; #100;
A = 8'h43; B = 8'hBC; #100;
A = 8'h43; B = 8'hBD; #100;
A = 8'h43; B = 8'hBE; #100;
A = 8'h43; B = 8'hBF; #100;
A = 8'h43; B = 8'hC0; #100;
A = 8'h43; B = 8'hC1; #100;
A = 8'h43; B = 8'hC2; #100;
A = 8'h43; B = 8'hC3; #100;
A = 8'h43; B = 8'hC4; #100;
A = 8'h43; B = 8'hC5; #100;
A = 8'h43; B = 8'hC6; #100;
A = 8'h43; B = 8'hC7; #100;
A = 8'h43; B = 8'hC8; #100;
A = 8'h43; B = 8'hC9; #100;
A = 8'h43; B = 8'hCA; #100;
A = 8'h43; B = 8'hCB; #100;
A = 8'h43; B = 8'hCC; #100;
A = 8'h43; B = 8'hCD; #100;
A = 8'h43; B = 8'hCE; #100;
A = 8'h43; B = 8'hCF; #100;
A = 8'h43; B = 8'hD0; #100;
A = 8'h43; B = 8'hD1; #100;
A = 8'h43; B = 8'hD2; #100;
A = 8'h43; B = 8'hD3; #100;
A = 8'h43; B = 8'hD4; #100;
A = 8'h43; B = 8'hD5; #100;
A = 8'h43; B = 8'hD6; #100;
A = 8'h43; B = 8'hD7; #100;
A = 8'h43; B = 8'hD8; #100;
A = 8'h43; B = 8'hD9; #100;
A = 8'h43; B = 8'hDA; #100;
A = 8'h43; B = 8'hDB; #100;
A = 8'h43; B = 8'hDC; #100;
A = 8'h43; B = 8'hDD; #100;
A = 8'h43; B = 8'hDE; #100;
A = 8'h43; B = 8'hDF; #100;
A = 8'h43; B = 8'hE0; #100;
A = 8'h43; B = 8'hE1; #100;
A = 8'h43; B = 8'hE2; #100;
A = 8'h43; B = 8'hE3; #100;
A = 8'h43; B = 8'hE4; #100;
A = 8'h43; B = 8'hE5; #100;
A = 8'h43; B = 8'hE6; #100;
A = 8'h43; B = 8'hE7; #100;
A = 8'h43; B = 8'hE8; #100;
A = 8'h43; B = 8'hE9; #100;
A = 8'h43; B = 8'hEA; #100;
A = 8'h43; B = 8'hEB; #100;
A = 8'h43; B = 8'hEC; #100;
A = 8'h43; B = 8'hED; #100;
A = 8'h43; B = 8'hEE; #100;
A = 8'h43; B = 8'hEF; #100;
A = 8'h43; B = 8'hF0; #100;
A = 8'h43; B = 8'hF1; #100;
A = 8'h43; B = 8'hF2; #100;
A = 8'h43; B = 8'hF3; #100;
A = 8'h43; B = 8'hF4; #100;
A = 8'h43; B = 8'hF5; #100;
A = 8'h43; B = 8'hF6; #100;
A = 8'h43; B = 8'hF7; #100;
A = 8'h43; B = 8'hF8; #100;
A = 8'h43; B = 8'hF9; #100;
A = 8'h43; B = 8'hFA; #100;
A = 8'h43; B = 8'hFB; #100;
A = 8'h43; B = 8'hFC; #100;
A = 8'h43; B = 8'hFD; #100;
A = 8'h43; B = 8'hFE; #100;
A = 8'h43; B = 8'hFF; #100;
A = 8'h44; B = 8'h0; #100;
A = 8'h44; B = 8'h1; #100;
A = 8'h44; B = 8'h2; #100;
A = 8'h44; B = 8'h3; #100;
A = 8'h44; B = 8'h4; #100;
A = 8'h44; B = 8'h5; #100;
A = 8'h44; B = 8'h6; #100;
A = 8'h44; B = 8'h7; #100;
A = 8'h44; B = 8'h8; #100;
A = 8'h44; B = 8'h9; #100;
A = 8'h44; B = 8'hA; #100;
A = 8'h44; B = 8'hB; #100;
A = 8'h44; B = 8'hC; #100;
A = 8'h44; B = 8'hD; #100;
A = 8'h44; B = 8'hE; #100;
A = 8'h44; B = 8'hF; #100;
A = 8'h44; B = 8'h10; #100;
A = 8'h44; B = 8'h11; #100;
A = 8'h44; B = 8'h12; #100;
A = 8'h44; B = 8'h13; #100;
A = 8'h44; B = 8'h14; #100;
A = 8'h44; B = 8'h15; #100;
A = 8'h44; B = 8'h16; #100;
A = 8'h44; B = 8'h17; #100;
A = 8'h44; B = 8'h18; #100;
A = 8'h44; B = 8'h19; #100;
A = 8'h44; B = 8'h1A; #100;
A = 8'h44; B = 8'h1B; #100;
A = 8'h44; B = 8'h1C; #100;
A = 8'h44; B = 8'h1D; #100;
A = 8'h44; B = 8'h1E; #100;
A = 8'h44; B = 8'h1F; #100;
A = 8'h44; B = 8'h20; #100;
A = 8'h44; B = 8'h21; #100;
A = 8'h44; B = 8'h22; #100;
A = 8'h44; B = 8'h23; #100;
A = 8'h44; B = 8'h24; #100;
A = 8'h44; B = 8'h25; #100;
A = 8'h44; B = 8'h26; #100;
A = 8'h44; B = 8'h27; #100;
A = 8'h44; B = 8'h28; #100;
A = 8'h44; B = 8'h29; #100;
A = 8'h44; B = 8'h2A; #100;
A = 8'h44; B = 8'h2B; #100;
A = 8'h44; B = 8'h2C; #100;
A = 8'h44; B = 8'h2D; #100;
A = 8'h44; B = 8'h2E; #100;
A = 8'h44; B = 8'h2F; #100;
A = 8'h44; B = 8'h30; #100;
A = 8'h44; B = 8'h31; #100;
A = 8'h44; B = 8'h32; #100;
A = 8'h44; B = 8'h33; #100;
A = 8'h44; B = 8'h34; #100;
A = 8'h44; B = 8'h35; #100;
A = 8'h44; B = 8'h36; #100;
A = 8'h44; B = 8'h37; #100;
A = 8'h44; B = 8'h38; #100;
A = 8'h44; B = 8'h39; #100;
A = 8'h44; B = 8'h3A; #100;
A = 8'h44; B = 8'h3B; #100;
A = 8'h44; B = 8'h3C; #100;
A = 8'h44; B = 8'h3D; #100;
A = 8'h44; B = 8'h3E; #100;
A = 8'h44; B = 8'h3F; #100;
A = 8'h44; B = 8'h40; #100;
A = 8'h44; B = 8'h41; #100;
A = 8'h44; B = 8'h42; #100;
A = 8'h44; B = 8'h43; #100;
A = 8'h44; B = 8'h44; #100;
A = 8'h44; B = 8'h45; #100;
A = 8'h44; B = 8'h46; #100;
A = 8'h44; B = 8'h47; #100;
A = 8'h44; B = 8'h48; #100;
A = 8'h44; B = 8'h49; #100;
A = 8'h44; B = 8'h4A; #100;
A = 8'h44; B = 8'h4B; #100;
A = 8'h44; B = 8'h4C; #100;
A = 8'h44; B = 8'h4D; #100;
A = 8'h44; B = 8'h4E; #100;
A = 8'h44; B = 8'h4F; #100;
A = 8'h44; B = 8'h50; #100;
A = 8'h44; B = 8'h51; #100;
A = 8'h44; B = 8'h52; #100;
A = 8'h44; B = 8'h53; #100;
A = 8'h44; B = 8'h54; #100;
A = 8'h44; B = 8'h55; #100;
A = 8'h44; B = 8'h56; #100;
A = 8'h44; B = 8'h57; #100;
A = 8'h44; B = 8'h58; #100;
A = 8'h44; B = 8'h59; #100;
A = 8'h44; B = 8'h5A; #100;
A = 8'h44; B = 8'h5B; #100;
A = 8'h44; B = 8'h5C; #100;
A = 8'h44; B = 8'h5D; #100;
A = 8'h44; B = 8'h5E; #100;
A = 8'h44; B = 8'h5F; #100;
A = 8'h44; B = 8'h60; #100;
A = 8'h44; B = 8'h61; #100;
A = 8'h44; B = 8'h62; #100;
A = 8'h44; B = 8'h63; #100;
A = 8'h44; B = 8'h64; #100;
A = 8'h44; B = 8'h65; #100;
A = 8'h44; B = 8'h66; #100;
A = 8'h44; B = 8'h67; #100;
A = 8'h44; B = 8'h68; #100;
A = 8'h44; B = 8'h69; #100;
A = 8'h44; B = 8'h6A; #100;
A = 8'h44; B = 8'h6B; #100;
A = 8'h44; B = 8'h6C; #100;
A = 8'h44; B = 8'h6D; #100;
A = 8'h44; B = 8'h6E; #100;
A = 8'h44; B = 8'h6F; #100;
A = 8'h44; B = 8'h70; #100;
A = 8'h44; B = 8'h71; #100;
A = 8'h44; B = 8'h72; #100;
A = 8'h44; B = 8'h73; #100;
A = 8'h44; B = 8'h74; #100;
A = 8'h44; B = 8'h75; #100;
A = 8'h44; B = 8'h76; #100;
A = 8'h44; B = 8'h77; #100;
A = 8'h44; B = 8'h78; #100;
A = 8'h44; B = 8'h79; #100;
A = 8'h44; B = 8'h7A; #100;
A = 8'h44; B = 8'h7B; #100;
A = 8'h44; B = 8'h7C; #100;
A = 8'h44; B = 8'h7D; #100;
A = 8'h44; B = 8'h7E; #100;
A = 8'h44; B = 8'h7F; #100;
A = 8'h44; B = 8'h80; #100;
A = 8'h44; B = 8'h81; #100;
A = 8'h44; B = 8'h82; #100;
A = 8'h44; B = 8'h83; #100;
A = 8'h44; B = 8'h84; #100;
A = 8'h44; B = 8'h85; #100;
A = 8'h44; B = 8'h86; #100;
A = 8'h44; B = 8'h87; #100;
A = 8'h44; B = 8'h88; #100;
A = 8'h44; B = 8'h89; #100;
A = 8'h44; B = 8'h8A; #100;
A = 8'h44; B = 8'h8B; #100;
A = 8'h44; B = 8'h8C; #100;
A = 8'h44; B = 8'h8D; #100;
A = 8'h44; B = 8'h8E; #100;
A = 8'h44; B = 8'h8F; #100;
A = 8'h44; B = 8'h90; #100;
A = 8'h44; B = 8'h91; #100;
A = 8'h44; B = 8'h92; #100;
A = 8'h44; B = 8'h93; #100;
A = 8'h44; B = 8'h94; #100;
A = 8'h44; B = 8'h95; #100;
A = 8'h44; B = 8'h96; #100;
A = 8'h44; B = 8'h97; #100;
A = 8'h44; B = 8'h98; #100;
A = 8'h44; B = 8'h99; #100;
A = 8'h44; B = 8'h9A; #100;
A = 8'h44; B = 8'h9B; #100;
A = 8'h44; B = 8'h9C; #100;
A = 8'h44; B = 8'h9D; #100;
A = 8'h44; B = 8'h9E; #100;
A = 8'h44; B = 8'h9F; #100;
A = 8'h44; B = 8'hA0; #100;
A = 8'h44; B = 8'hA1; #100;
A = 8'h44; B = 8'hA2; #100;
A = 8'h44; B = 8'hA3; #100;
A = 8'h44; B = 8'hA4; #100;
A = 8'h44; B = 8'hA5; #100;
A = 8'h44; B = 8'hA6; #100;
A = 8'h44; B = 8'hA7; #100;
A = 8'h44; B = 8'hA8; #100;
A = 8'h44; B = 8'hA9; #100;
A = 8'h44; B = 8'hAA; #100;
A = 8'h44; B = 8'hAB; #100;
A = 8'h44; B = 8'hAC; #100;
A = 8'h44; B = 8'hAD; #100;
A = 8'h44; B = 8'hAE; #100;
A = 8'h44; B = 8'hAF; #100;
A = 8'h44; B = 8'hB0; #100;
A = 8'h44; B = 8'hB1; #100;
A = 8'h44; B = 8'hB2; #100;
A = 8'h44; B = 8'hB3; #100;
A = 8'h44; B = 8'hB4; #100;
A = 8'h44; B = 8'hB5; #100;
A = 8'h44; B = 8'hB6; #100;
A = 8'h44; B = 8'hB7; #100;
A = 8'h44; B = 8'hB8; #100;
A = 8'h44; B = 8'hB9; #100;
A = 8'h44; B = 8'hBA; #100;
A = 8'h44; B = 8'hBB; #100;
A = 8'h44; B = 8'hBC; #100;
A = 8'h44; B = 8'hBD; #100;
A = 8'h44; B = 8'hBE; #100;
A = 8'h44; B = 8'hBF; #100;
A = 8'h44; B = 8'hC0; #100;
A = 8'h44; B = 8'hC1; #100;
A = 8'h44; B = 8'hC2; #100;
A = 8'h44; B = 8'hC3; #100;
A = 8'h44; B = 8'hC4; #100;
A = 8'h44; B = 8'hC5; #100;
A = 8'h44; B = 8'hC6; #100;
A = 8'h44; B = 8'hC7; #100;
A = 8'h44; B = 8'hC8; #100;
A = 8'h44; B = 8'hC9; #100;
A = 8'h44; B = 8'hCA; #100;
A = 8'h44; B = 8'hCB; #100;
A = 8'h44; B = 8'hCC; #100;
A = 8'h44; B = 8'hCD; #100;
A = 8'h44; B = 8'hCE; #100;
A = 8'h44; B = 8'hCF; #100;
A = 8'h44; B = 8'hD0; #100;
A = 8'h44; B = 8'hD1; #100;
A = 8'h44; B = 8'hD2; #100;
A = 8'h44; B = 8'hD3; #100;
A = 8'h44; B = 8'hD4; #100;
A = 8'h44; B = 8'hD5; #100;
A = 8'h44; B = 8'hD6; #100;
A = 8'h44; B = 8'hD7; #100;
A = 8'h44; B = 8'hD8; #100;
A = 8'h44; B = 8'hD9; #100;
A = 8'h44; B = 8'hDA; #100;
A = 8'h44; B = 8'hDB; #100;
A = 8'h44; B = 8'hDC; #100;
A = 8'h44; B = 8'hDD; #100;
A = 8'h44; B = 8'hDE; #100;
A = 8'h44; B = 8'hDF; #100;
A = 8'h44; B = 8'hE0; #100;
A = 8'h44; B = 8'hE1; #100;
A = 8'h44; B = 8'hE2; #100;
A = 8'h44; B = 8'hE3; #100;
A = 8'h44; B = 8'hE4; #100;
A = 8'h44; B = 8'hE5; #100;
A = 8'h44; B = 8'hE6; #100;
A = 8'h44; B = 8'hE7; #100;
A = 8'h44; B = 8'hE8; #100;
A = 8'h44; B = 8'hE9; #100;
A = 8'h44; B = 8'hEA; #100;
A = 8'h44; B = 8'hEB; #100;
A = 8'h44; B = 8'hEC; #100;
A = 8'h44; B = 8'hED; #100;
A = 8'h44; B = 8'hEE; #100;
A = 8'h44; B = 8'hEF; #100;
A = 8'h44; B = 8'hF0; #100;
A = 8'h44; B = 8'hF1; #100;
A = 8'h44; B = 8'hF2; #100;
A = 8'h44; B = 8'hF3; #100;
A = 8'h44; B = 8'hF4; #100;
A = 8'h44; B = 8'hF5; #100;
A = 8'h44; B = 8'hF6; #100;
A = 8'h44; B = 8'hF7; #100;
A = 8'h44; B = 8'hF8; #100;
A = 8'h44; B = 8'hF9; #100;
A = 8'h44; B = 8'hFA; #100;
A = 8'h44; B = 8'hFB; #100;
A = 8'h44; B = 8'hFC; #100;
A = 8'h44; B = 8'hFD; #100;
A = 8'h44; B = 8'hFE; #100;
A = 8'h44; B = 8'hFF; #100;
A = 8'h45; B = 8'h0; #100;
A = 8'h45; B = 8'h1; #100;
A = 8'h45; B = 8'h2; #100;
A = 8'h45; B = 8'h3; #100;
A = 8'h45; B = 8'h4; #100;
A = 8'h45; B = 8'h5; #100;
A = 8'h45; B = 8'h6; #100;
A = 8'h45; B = 8'h7; #100;
A = 8'h45; B = 8'h8; #100;
A = 8'h45; B = 8'h9; #100;
A = 8'h45; B = 8'hA; #100;
A = 8'h45; B = 8'hB; #100;
A = 8'h45; B = 8'hC; #100;
A = 8'h45; B = 8'hD; #100;
A = 8'h45; B = 8'hE; #100;
A = 8'h45; B = 8'hF; #100;
A = 8'h45; B = 8'h10; #100;
A = 8'h45; B = 8'h11; #100;
A = 8'h45; B = 8'h12; #100;
A = 8'h45; B = 8'h13; #100;
A = 8'h45; B = 8'h14; #100;
A = 8'h45; B = 8'h15; #100;
A = 8'h45; B = 8'h16; #100;
A = 8'h45; B = 8'h17; #100;
A = 8'h45; B = 8'h18; #100;
A = 8'h45; B = 8'h19; #100;
A = 8'h45; B = 8'h1A; #100;
A = 8'h45; B = 8'h1B; #100;
A = 8'h45; B = 8'h1C; #100;
A = 8'h45; B = 8'h1D; #100;
A = 8'h45; B = 8'h1E; #100;
A = 8'h45; B = 8'h1F; #100;
A = 8'h45; B = 8'h20; #100;
A = 8'h45; B = 8'h21; #100;
A = 8'h45; B = 8'h22; #100;
A = 8'h45; B = 8'h23; #100;
A = 8'h45; B = 8'h24; #100;
A = 8'h45; B = 8'h25; #100;
A = 8'h45; B = 8'h26; #100;
A = 8'h45; B = 8'h27; #100;
A = 8'h45; B = 8'h28; #100;
A = 8'h45; B = 8'h29; #100;
A = 8'h45; B = 8'h2A; #100;
A = 8'h45; B = 8'h2B; #100;
A = 8'h45; B = 8'h2C; #100;
A = 8'h45; B = 8'h2D; #100;
A = 8'h45; B = 8'h2E; #100;
A = 8'h45; B = 8'h2F; #100;
A = 8'h45; B = 8'h30; #100;
A = 8'h45; B = 8'h31; #100;
A = 8'h45; B = 8'h32; #100;
A = 8'h45; B = 8'h33; #100;
A = 8'h45; B = 8'h34; #100;
A = 8'h45; B = 8'h35; #100;
A = 8'h45; B = 8'h36; #100;
A = 8'h45; B = 8'h37; #100;
A = 8'h45; B = 8'h38; #100;
A = 8'h45; B = 8'h39; #100;
A = 8'h45; B = 8'h3A; #100;
A = 8'h45; B = 8'h3B; #100;
A = 8'h45; B = 8'h3C; #100;
A = 8'h45; B = 8'h3D; #100;
A = 8'h45; B = 8'h3E; #100;
A = 8'h45; B = 8'h3F; #100;
A = 8'h45; B = 8'h40; #100;
A = 8'h45; B = 8'h41; #100;
A = 8'h45; B = 8'h42; #100;
A = 8'h45; B = 8'h43; #100;
A = 8'h45; B = 8'h44; #100;
A = 8'h45; B = 8'h45; #100;
A = 8'h45; B = 8'h46; #100;
A = 8'h45; B = 8'h47; #100;
A = 8'h45; B = 8'h48; #100;
A = 8'h45; B = 8'h49; #100;
A = 8'h45; B = 8'h4A; #100;
A = 8'h45; B = 8'h4B; #100;
A = 8'h45; B = 8'h4C; #100;
A = 8'h45; B = 8'h4D; #100;
A = 8'h45; B = 8'h4E; #100;
A = 8'h45; B = 8'h4F; #100;
A = 8'h45; B = 8'h50; #100;
A = 8'h45; B = 8'h51; #100;
A = 8'h45; B = 8'h52; #100;
A = 8'h45; B = 8'h53; #100;
A = 8'h45; B = 8'h54; #100;
A = 8'h45; B = 8'h55; #100;
A = 8'h45; B = 8'h56; #100;
A = 8'h45; B = 8'h57; #100;
A = 8'h45; B = 8'h58; #100;
A = 8'h45; B = 8'h59; #100;
A = 8'h45; B = 8'h5A; #100;
A = 8'h45; B = 8'h5B; #100;
A = 8'h45; B = 8'h5C; #100;
A = 8'h45; B = 8'h5D; #100;
A = 8'h45; B = 8'h5E; #100;
A = 8'h45; B = 8'h5F; #100;
A = 8'h45; B = 8'h60; #100;
A = 8'h45; B = 8'h61; #100;
A = 8'h45; B = 8'h62; #100;
A = 8'h45; B = 8'h63; #100;
A = 8'h45; B = 8'h64; #100;
A = 8'h45; B = 8'h65; #100;
A = 8'h45; B = 8'h66; #100;
A = 8'h45; B = 8'h67; #100;
A = 8'h45; B = 8'h68; #100;
A = 8'h45; B = 8'h69; #100;
A = 8'h45; B = 8'h6A; #100;
A = 8'h45; B = 8'h6B; #100;
A = 8'h45; B = 8'h6C; #100;
A = 8'h45; B = 8'h6D; #100;
A = 8'h45; B = 8'h6E; #100;
A = 8'h45; B = 8'h6F; #100;
A = 8'h45; B = 8'h70; #100;
A = 8'h45; B = 8'h71; #100;
A = 8'h45; B = 8'h72; #100;
A = 8'h45; B = 8'h73; #100;
A = 8'h45; B = 8'h74; #100;
A = 8'h45; B = 8'h75; #100;
A = 8'h45; B = 8'h76; #100;
A = 8'h45; B = 8'h77; #100;
A = 8'h45; B = 8'h78; #100;
A = 8'h45; B = 8'h79; #100;
A = 8'h45; B = 8'h7A; #100;
A = 8'h45; B = 8'h7B; #100;
A = 8'h45; B = 8'h7C; #100;
A = 8'h45; B = 8'h7D; #100;
A = 8'h45; B = 8'h7E; #100;
A = 8'h45; B = 8'h7F; #100;
A = 8'h45; B = 8'h80; #100;
A = 8'h45; B = 8'h81; #100;
A = 8'h45; B = 8'h82; #100;
A = 8'h45; B = 8'h83; #100;
A = 8'h45; B = 8'h84; #100;
A = 8'h45; B = 8'h85; #100;
A = 8'h45; B = 8'h86; #100;
A = 8'h45; B = 8'h87; #100;
A = 8'h45; B = 8'h88; #100;
A = 8'h45; B = 8'h89; #100;
A = 8'h45; B = 8'h8A; #100;
A = 8'h45; B = 8'h8B; #100;
A = 8'h45; B = 8'h8C; #100;
A = 8'h45; B = 8'h8D; #100;
A = 8'h45; B = 8'h8E; #100;
A = 8'h45; B = 8'h8F; #100;
A = 8'h45; B = 8'h90; #100;
A = 8'h45; B = 8'h91; #100;
A = 8'h45; B = 8'h92; #100;
A = 8'h45; B = 8'h93; #100;
A = 8'h45; B = 8'h94; #100;
A = 8'h45; B = 8'h95; #100;
A = 8'h45; B = 8'h96; #100;
A = 8'h45; B = 8'h97; #100;
A = 8'h45; B = 8'h98; #100;
A = 8'h45; B = 8'h99; #100;
A = 8'h45; B = 8'h9A; #100;
A = 8'h45; B = 8'h9B; #100;
A = 8'h45; B = 8'h9C; #100;
A = 8'h45; B = 8'h9D; #100;
A = 8'h45; B = 8'h9E; #100;
A = 8'h45; B = 8'h9F; #100;
A = 8'h45; B = 8'hA0; #100;
A = 8'h45; B = 8'hA1; #100;
A = 8'h45; B = 8'hA2; #100;
A = 8'h45; B = 8'hA3; #100;
A = 8'h45; B = 8'hA4; #100;
A = 8'h45; B = 8'hA5; #100;
A = 8'h45; B = 8'hA6; #100;
A = 8'h45; B = 8'hA7; #100;
A = 8'h45; B = 8'hA8; #100;
A = 8'h45; B = 8'hA9; #100;
A = 8'h45; B = 8'hAA; #100;
A = 8'h45; B = 8'hAB; #100;
A = 8'h45; B = 8'hAC; #100;
A = 8'h45; B = 8'hAD; #100;
A = 8'h45; B = 8'hAE; #100;
A = 8'h45; B = 8'hAF; #100;
A = 8'h45; B = 8'hB0; #100;
A = 8'h45; B = 8'hB1; #100;
A = 8'h45; B = 8'hB2; #100;
A = 8'h45; B = 8'hB3; #100;
A = 8'h45; B = 8'hB4; #100;
A = 8'h45; B = 8'hB5; #100;
A = 8'h45; B = 8'hB6; #100;
A = 8'h45; B = 8'hB7; #100;
A = 8'h45; B = 8'hB8; #100;
A = 8'h45; B = 8'hB9; #100;
A = 8'h45; B = 8'hBA; #100;
A = 8'h45; B = 8'hBB; #100;
A = 8'h45; B = 8'hBC; #100;
A = 8'h45; B = 8'hBD; #100;
A = 8'h45; B = 8'hBE; #100;
A = 8'h45; B = 8'hBF; #100;
A = 8'h45; B = 8'hC0; #100;
A = 8'h45; B = 8'hC1; #100;
A = 8'h45; B = 8'hC2; #100;
A = 8'h45; B = 8'hC3; #100;
A = 8'h45; B = 8'hC4; #100;
A = 8'h45; B = 8'hC5; #100;
A = 8'h45; B = 8'hC6; #100;
A = 8'h45; B = 8'hC7; #100;
A = 8'h45; B = 8'hC8; #100;
A = 8'h45; B = 8'hC9; #100;
A = 8'h45; B = 8'hCA; #100;
A = 8'h45; B = 8'hCB; #100;
A = 8'h45; B = 8'hCC; #100;
A = 8'h45; B = 8'hCD; #100;
A = 8'h45; B = 8'hCE; #100;
A = 8'h45; B = 8'hCF; #100;
A = 8'h45; B = 8'hD0; #100;
A = 8'h45; B = 8'hD1; #100;
A = 8'h45; B = 8'hD2; #100;
A = 8'h45; B = 8'hD3; #100;
A = 8'h45; B = 8'hD4; #100;
A = 8'h45; B = 8'hD5; #100;
A = 8'h45; B = 8'hD6; #100;
A = 8'h45; B = 8'hD7; #100;
A = 8'h45; B = 8'hD8; #100;
A = 8'h45; B = 8'hD9; #100;
A = 8'h45; B = 8'hDA; #100;
A = 8'h45; B = 8'hDB; #100;
A = 8'h45; B = 8'hDC; #100;
A = 8'h45; B = 8'hDD; #100;
A = 8'h45; B = 8'hDE; #100;
A = 8'h45; B = 8'hDF; #100;
A = 8'h45; B = 8'hE0; #100;
A = 8'h45; B = 8'hE1; #100;
A = 8'h45; B = 8'hE2; #100;
A = 8'h45; B = 8'hE3; #100;
A = 8'h45; B = 8'hE4; #100;
A = 8'h45; B = 8'hE5; #100;
A = 8'h45; B = 8'hE6; #100;
A = 8'h45; B = 8'hE7; #100;
A = 8'h45; B = 8'hE8; #100;
A = 8'h45; B = 8'hE9; #100;
A = 8'h45; B = 8'hEA; #100;
A = 8'h45; B = 8'hEB; #100;
A = 8'h45; B = 8'hEC; #100;
A = 8'h45; B = 8'hED; #100;
A = 8'h45; B = 8'hEE; #100;
A = 8'h45; B = 8'hEF; #100;
A = 8'h45; B = 8'hF0; #100;
A = 8'h45; B = 8'hF1; #100;
A = 8'h45; B = 8'hF2; #100;
A = 8'h45; B = 8'hF3; #100;
A = 8'h45; B = 8'hF4; #100;
A = 8'h45; B = 8'hF5; #100;
A = 8'h45; B = 8'hF6; #100;
A = 8'h45; B = 8'hF7; #100;
A = 8'h45; B = 8'hF8; #100;
A = 8'h45; B = 8'hF9; #100;
A = 8'h45; B = 8'hFA; #100;
A = 8'h45; B = 8'hFB; #100;
A = 8'h45; B = 8'hFC; #100;
A = 8'h45; B = 8'hFD; #100;
A = 8'h45; B = 8'hFE; #100;
A = 8'h45; B = 8'hFF; #100;
A = 8'h46; B = 8'h0; #100;
A = 8'h46; B = 8'h1; #100;
A = 8'h46; B = 8'h2; #100;
A = 8'h46; B = 8'h3; #100;
A = 8'h46; B = 8'h4; #100;
A = 8'h46; B = 8'h5; #100;
A = 8'h46; B = 8'h6; #100;
A = 8'h46; B = 8'h7; #100;
A = 8'h46; B = 8'h8; #100;
A = 8'h46; B = 8'h9; #100;
A = 8'h46; B = 8'hA; #100;
A = 8'h46; B = 8'hB; #100;
A = 8'h46; B = 8'hC; #100;
A = 8'h46; B = 8'hD; #100;
A = 8'h46; B = 8'hE; #100;
A = 8'h46; B = 8'hF; #100;
A = 8'h46; B = 8'h10; #100;
A = 8'h46; B = 8'h11; #100;
A = 8'h46; B = 8'h12; #100;
A = 8'h46; B = 8'h13; #100;
A = 8'h46; B = 8'h14; #100;
A = 8'h46; B = 8'h15; #100;
A = 8'h46; B = 8'h16; #100;
A = 8'h46; B = 8'h17; #100;
A = 8'h46; B = 8'h18; #100;
A = 8'h46; B = 8'h19; #100;
A = 8'h46; B = 8'h1A; #100;
A = 8'h46; B = 8'h1B; #100;
A = 8'h46; B = 8'h1C; #100;
A = 8'h46; B = 8'h1D; #100;
A = 8'h46; B = 8'h1E; #100;
A = 8'h46; B = 8'h1F; #100;
A = 8'h46; B = 8'h20; #100;
A = 8'h46; B = 8'h21; #100;
A = 8'h46; B = 8'h22; #100;
A = 8'h46; B = 8'h23; #100;
A = 8'h46; B = 8'h24; #100;
A = 8'h46; B = 8'h25; #100;
A = 8'h46; B = 8'h26; #100;
A = 8'h46; B = 8'h27; #100;
A = 8'h46; B = 8'h28; #100;
A = 8'h46; B = 8'h29; #100;
A = 8'h46; B = 8'h2A; #100;
A = 8'h46; B = 8'h2B; #100;
A = 8'h46; B = 8'h2C; #100;
A = 8'h46; B = 8'h2D; #100;
A = 8'h46; B = 8'h2E; #100;
A = 8'h46; B = 8'h2F; #100;
A = 8'h46; B = 8'h30; #100;
A = 8'h46; B = 8'h31; #100;
A = 8'h46; B = 8'h32; #100;
A = 8'h46; B = 8'h33; #100;
A = 8'h46; B = 8'h34; #100;
A = 8'h46; B = 8'h35; #100;
A = 8'h46; B = 8'h36; #100;
A = 8'h46; B = 8'h37; #100;
A = 8'h46; B = 8'h38; #100;
A = 8'h46; B = 8'h39; #100;
A = 8'h46; B = 8'h3A; #100;
A = 8'h46; B = 8'h3B; #100;
A = 8'h46; B = 8'h3C; #100;
A = 8'h46; B = 8'h3D; #100;
A = 8'h46; B = 8'h3E; #100;
A = 8'h46; B = 8'h3F; #100;
A = 8'h46; B = 8'h40; #100;
A = 8'h46; B = 8'h41; #100;
A = 8'h46; B = 8'h42; #100;
A = 8'h46; B = 8'h43; #100;
A = 8'h46; B = 8'h44; #100;
A = 8'h46; B = 8'h45; #100;
A = 8'h46; B = 8'h46; #100;
A = 8'h46; B = 8'h47; #100;
A = 8'h46; B = 8'h48; #100;
A = 8'h46; B = 8'h49; #100;
A = 8'h46; B = 8'h4A; #100;
A = 8'h46; B = 8'h4B; #100;
A = 8'h46; B = 8'h4C; #100;
A = 8'h46; B = 8'h4D; #100;
A = 8'h46; B = 8'h4E; #100;
A = 8'h46; B = 8'h4F; #100;
A = 8'h46; B = 8'h50; #100;
A = 8'h46; B = 8'h51; #100;
A = 8'h46; B = 8'h52; #100;
A = 8'h46; B = 8'h53; #100;
A = 8'h46; B = 8'h54; #100;
A = 8'h46; B = 8'h55; #100;
A = 8'h46; B = 8'h56; #100;
A = 8'h46; B = 8'h57; #100;
A = 8'h46; B = 8'h58; #100;
A = 8'h46; B = 8'h59; #100;
A = 8'h46; B = 8'h5A; #100;
A = 8'h46; B = 8'h5B; #100;
A = 8'h46; B = 8'h5C; #100;
A = 8'h46; B = 8'h5D; #100;
A = 8'h46; B = 8'h5E; #100;
A = 8'h46; B = 8'h5F; #100;
A = 8'h46; B = 8'h60; #100;
A = 8'h46; B = 8'h61; #100;
A = 8'h46; B = 8'h62; #100;
A = 8'h46; B = 8'h63; #100;
A = 8'h46; B = 8'h64; #100;
A = 8'h46; B = 8'h65; #100;
A = 8'h46; B = 8'h66; #100;
A = 8'h46; B = 8'h67; #100;
A = 8'h46; B = 8'h68; #100;
A = 8'h46; B = 8'h69; #100;
A = 8'h46; B = 8'h6A; #100;
A = 8'h46; B = 8'h6B; #100;
A = 8'h46; B = 8'h6C; #100;
A = 8'h46; B = 8'h6D; #100;
A = 8'h46; B = 8'h6E; #100;
A = 8'h46; B = 8'h6F; #100;
A = 8'h46; B = 8'h70; #100;
A = 8'h46; B = 8'h71; #100;
A = 8'h46; B = 8'h72; #100;
A = 8'h46; B = 8'h73; #100;
A = 8'h46; B = 8'h74; #100;
A = 8'h46; B = 8'h75; #100;
A = 8'h46; B = 8'h76; #100;
A = 8'h46; B = 8'h77; #100;
A = 8'h46; B = 8'h78; #100;
A = 8'h46; B = 8'h79; #100;
A = 8'h46; B = 8'h7A; #100;
A = 8'h46; B = 8'h7B; #100;
A = 8'h46; B = 8'h7C; #100;
A = 8'h46; B = 8'h7D; #100;
A = 8'h46; B = 8'h7E; #100;
A = 8'h46; B = 8'h7F; #100;
A = 8'h46; B = 8'h80; #100;
A = 8'h46; B = 8'h81; #100;
A = 8'h46; B = 8'h82; #100;
A = 8'h46; B = 8'h83; #100;
A = 8'h46; B = 8'h84; #100;
A = 8'h46; B = 8'h85; #100;
A = 8'h46; B = 8'h86; #100;
A = 8'h46; B = 8'h87; #100;
A = 8'h46; B = 8'h88; #100;
A = 8'h46; B = 8'h89; #100;
A = 8'h46; B = 8'h8A; #100;
A = 8'h46; B = 8'h8B; #100;
A = 8'h46; B = 8'h8C; #100;
A = 8'h46; B = 8'h8D; #100;
A = 8'h46; B = 8'h8E; #100;
A = 8'h46; B = 8'h8F; #100;
A = 8'h46; B = 8'h90; #100;
A = 8'h46; B = 8'h91; #100;
A = 8'h46; B = 8'h92; #100;
A = 8'h46; B = 8'h93; #100;
A = 8'h46; B = 8'h94; #100;
A = 8'h46; B = 8'h95; #100;
A = 8'h46; B = 8'h96; #100;
A = 8'h46; B = 8'h97; #100;
A = 8'h46; B = 8'h98; #100;
A = 8'h46; B = 8'h99; #100;
A = 8'h46; B = 8'h9A; #100;
A = 8'h46; B = 8'h9B; #100;
A = 8'h46; B = 8'h9C; #100;
A = 8'h46; B = 8'h9D; #100;
A = 8'h46; B = 8'h9E; #100;
A = 8'h46; B = 8'h9F; #100;
A = 8'h46; B = 8'hA0; #100;
A = 8'h46; B = 8'hA1; #100;
A = 8'h46; B = 8'hA2; #100;
A = 8'h46; B = 8'hA3; #100;
A = 8'h46; B = 8'hA4; #100;
A = 8'h46; B = 8'hA5; #100;
A = 8'h46; B = 8'hA6; #100;
A = 8'h46; B = 8'hA7; #100;
A = 8'h46; B = 8'hA8; #100;
A = 8'h46; B = 8'hA9; #100;
A = 8'h46; B = 8'hAA; #100;
A = 8'h46; B = 8'hAB; #100;
A = 8'h46; B = 8'hAC; #100;
A = 8'h46; B = 8'hAD; #100;
A = 8'h46; B = 8'hAE; #100;
A = 8'h46; B = 8'hAF; #100;
A = 8'h46; B = 8'hB0; #100;
A = 8'h46; B = 8'hB1; #100;
A = 8'h46; B = 8'hB2; #100;
A = 8'h46; B = 8'hB3; #100;
A = 8'h46; B = 8'hB4; #100;
A = 8'h46; B = 8'hB5; #100;
A = 8'h46; B = 8'hB6; #100;
A = 8'h46; B = 8'hB7; #100;
A = 8'h46; B = 8'hB8; #100;
A = 8'h46; B = 8'hB9; #100;
A = 8'h46; B = 8'hBA; #100;
A = 8'h46; B = 8'hBB; #100;
A = 8'h46; B = 8'hBC; #100;
A = 8'h46; B = 8'hBD; #100;
A = 8'h46; B = 8'hBE; #100;
A = 8'h46; B = 8'hBF; #100;
A = 8'h46; B = 8'hC0; #100;
A = 8'h46; B = 8'hC1; #100;
A = 8'h46; B = 8'hC2; #100;
A = 8'h46; B = 8'hC3; #100;
A = 8'h46; B = 8'hC4; #100;
A = 8'h46; B = 8'hC5; #100;
A = 8'h46; B = 8'hC6; #100;
A = 8'h46; B = 8'hC7; #100;
A = 8'h46; B = 8'hC8; #100;
A = 8'h46; B = 8'hC9; #100;
A = 8'h46; B = 8'hCA; #100;
A = 8'h46; B = 8'hCB; #100;
A = 8'h46; B = 8'hCC; #100;
A = 8'h46; B = 8'hCD; #100;
A = 8'h46; B = 8'hCE; #100;
A = 8'h46; B = 8'hCF; #100;
A = 8'h46; B = 8'hD0; #100;
A = 8'h46; B = 8'hD1; #100;
A = 8'h46; B = 8'hD2; #100;
A = 8'h46; B = 8'hD3; #100;
A = 8'h46; B = 8'hD4; #100;
A = 8'h46; B = 8'hD5; #100;
A = 8'h46; B = 8'hD6; #100;
A = 8'h46; B = 8'hD7; #100;
A = 8'h46; B = 8'hD8; #100;
A = 8'h46; B = 8'hD9; #100;
A = 8'h46; B = 8'hDA; #100;
A = 8'h46; B = 8'hDB; #100;
A = 8'h46; B = 8'hDC; #100;
A = 8'h46; B = 8'hDD; #100;
A = 8'h46; B = 8'hDE; #100;
A = 8'h46; B = 8'hDF; #100;
A = 8'h46; B = 8'hE0; #100;
A = 8'h46; B = 8'hE1; #100;
A = 8'h46; B = 8'hE2; #100;
A = 8'h46; B = 8'hE3; #100;
A = 8'h46; B = 8'hE4; #100;
A = 8'h46; B = 8'hE5; #100;
A = 8'h46; B = 8'hE6; #100;
A = 8'h46; B = 8'hE7; #100;
A = 8'h46; B = 8'hE8; #100;
A = 8'h46; B = 8'hE9; #100;
A = 8'h46; B = 8'hEA; #100;
A = 8'h46; B = 8'hEB; #100;
A = 8'h46; B = 8'hEC; #100;
A = 8'h46; B = 8'hED; #100;
A = 8'h46; B = 8'hEE; #100;
A = 8'h46; B = 8'hEF; #100;
A = 8'h46; B = 8'hF0; #100;
A = 8'h46; B = 8'hF1; #100;
A = 8'h46; B = 8'hF2; #100;
A = 8'h46; B = 8'hF3; #100;
A = 8'h46; B = 8'hF4; #100;
A = 8'h46; B = 8'hF5; #100;
A = 8'h46; B = 8'hF6; #100;
A = 8'h46; B = 8'hF7; #100;
A = 8'h46; B = 8'hF8; #100;
A = 8'h46; B = 8'hF9; #100;
A = 8'h46; B = 8'hFA; #100;
A = 8'h46; B = 8'hFB; #100;
A = 8'h46; B = 8'hFC; #100;
A = 8'h46; B = 8'hFD; #100;
A = 8'h46; B = 8'hFE; #100;
A = 8'h46; B = 8'hFF; #100;
A = 8'h47; B = 8'h0; #100;
A = 8'h47; B = 8'h1; #100;
A = 8'h47; B = 8'h2; #100;
A = 8'h47; B = 8'h3; #100;
A = 8'h47; B = 8'h4; #100;
A = 8'h47; B = 8'h5; #100;
A = 8'h47; B = 8'h6; #100;
A = 8'h47; B = 8'h7; #100;
A = 8'h47; B = 8'h8; #100;
A = 8'h47; B = 8'h9; #100;
A = 8'h47; B = 8'hA; #100;
A = 8'h47; B = 8'hB; #100;
A = 8'h47; B = 8'hC; #100;
A = 8'h47; B = 8'hD; #100;
A = 8'h47; B = 8'hE; #100;
A = 8'h47; B = 8'hF; #100;
A = 8'h47; B = 8'h10; #100;
A = 8'h47; B = 8'h11; #100;
A = 8'h47; B = 8'h12; #100;
A = 8'h47; B = 8'h13; #100;
A = 8'h47; B = 8'h14; #100;
A = 8'h47; B = 8'h15; #100;
A = 8'h47; B = 8'h16; #100;
A = 8'h47; B = 8'h17; #100;
A = 8'h47; B = 8'h18; #100;
A = 8'h47; B = 8'h19; #100;
A = 8'h47; B = 8'h1A; #100;
A = 8'h47; B = 8'h1B; #100;
A = 8'h47; B = 8'h1C; #100;
A = 8'h47; B = 8'h1D; #100;
A = 8'h47; B = 8'h1E; #100;
A = 8'h47; B = 8'h1F; #100;
A = 8'h47; B = 8'h20; #100;
A = 8'h47; B = 8'h21; #100;
A = 8'h47; B = 8'h22; #100;
A = 8'h47; B = 8'h23; #100;
A = 8'h47; B = 8'h24; #100;
A = 8'h47; B = 8'h25; #100;
A = 8'h47; B = 8'h26; #100;
A = 8'h47; B = 8'h27; #100;
A = 8'h47; B = 8'h28; #100;
A = 8'h47; B = 8'h29; #100;
A = 8'h47; B = 8'h2A; #100;
A = 8'h47; B = 8'h2B; #100;
A = 8'h47; B = 8'h2C; #100;
A = 8'h47; B = 8'h2D; #100;
A = 8'h47; B = 8'h2E; #100;
A = 8'h47; B = 8'h2F; #100;
A = 8'h47; B = 8'h30; #100;
A = 8'h47; B = 8'h31; #100;
A = 8'h47; B = 8'h32; #100;
A = 8'h47; B = 8'h33; #100;
A = 8'h47; B = 8'h34; #100;
A = 8'h47; B = 8'h35; #100;
A = 8'h47; B = 8'h36; #100;
A = 8'h47; B = 8'h37; #100;
A = 8'h47; B = 8'h38; #100;
A = 8'h47; B = 8'h39; #100;
A = 8'h47; B = 8'h3A; #100;
A = 8'h47; B = 8'h3B; #100;
A = 8'h47; B = 8'h3C; #100;
A = 8'h47; B = 8'h3D; #100;
A = 8'h47; B = 8'h3E; #100;
A = 8'h47; B = 8'h3F; #100;
A = 8'h47; B = 8'h40; #100;
A = 8'h47; B = 8'h41; #100;
A = 8'h47; B = 8'h42; #100;
A = 8'h47; B = 8'h43; #100;
A = 8'h47; B = 8'h44; #100;
A = 8'h47; B = 8'h45; #100;
A = 8'h47; B = 8'h46; #100;
A = 8'h47; B = 8'h47; #100;
A = 8'h47; B = 8'h48; #100;
A = 8'h47; B = 8'h49; #100;
A = 8'h47; B = 8'h4A; #100;
A = 8'h47; B = 8'h4B; #100;
A = 8'h47; B = 8'h4C; #100;
A = 8'h47; B = 8'h4D; #100;
A = 8'h47; B = 8'h4E; #100;
A = 8'h47; B = 8'h4F; #100;
A = 8'h47; B = 8'h50; #100;
A = 8'h47; B = 8'h51; #100;
A = 8'h47; B = 8'h52; #100;
A = 8'h47; B = 8'h53; #100;
A = 8'h47; B = 8'h54; #100;
A = 8'h47; B = 8'h55; #100;
A = 8'h47; B = 8'h56; #100;
A = 8'h47; B = 8'h57; #100;
A = 8'h47; B = 8'h58; #100;
A = 8'h47; B = 8'h59; #100;
A = 8'h47; B = 8'h5A; #100;
A = 8'h47; B = 8'h5B; #100;
A = 8'h47; B = 8'h5C; #100;
A = 8'h47; B = 8'h5D; #100;
A = 8'h47; B = 8'h5E; #100;
A = 8'h47; B = 8'h5F; #100;
A = 8'h47; B = 8'h60; #100;
A = 8'h47; B = 8'h61; #100;
A = 8'h47; B = 8'h62; #100;
A = 8'h47; B = 8'h63; #100;
A = 8'h47; B = 8'h64; #100;
A = 8'h47; B = 8'h65; #100;
A = 8'h47; B = 8'h66; #100;
A = 8'h47; B = 8'h67; #100;
A = 8'h47; B = 8'h68; #100;
A = 8'h47; B = 8'h69; #100;
A = 8'h47; B = 8'h6A; #100;
A = 8'h47; B = 8'h6B; #100;
A = 8'h47; B = 8'h6C; #100;
A = 8'h47; B = 8'h6D; #100;
A = 8'h47; B = 8'h6E; #100;
A = 8'h47; B = 8'h6F; #100;
A = 8'h47; B = 8'h70; #100;
A = 8'h47; B = 8'h71; #100;
A = 8'h47; B = 8'h72; #100;
A = 8'h47; B = 8'h73; #100;
A = 8'h47; B = 8'h74; #100;
A = 8'h47; B = 8'h75; #100;
A = 8'h47; B = 8'h76; #100;
A = 8'h47; B = 8'h77; #100;
A = 8'h47; B = 8'h78; #100;
A = 8'h47; B = 8'h79; #100;
A = 8'h47; B = 8'h7A; #100;
A = 8'h47; B = 8'h7B; #100;
A = 8'h47; B = 8'h7C; #100;
A = 8'h47; B = 8'h7D; #100;
A = 8'h47; B = 8'h7E; #100;
A = 8'h47; B = 8'h7F; #100;
A = 8'h47; B = 8'h80; #100;
A = 8'h47; B = 8'h81; #100;
A = 8'h47; B = 8'h82; #100;
A = 8'h47; B = 8'h83; #100;
A = 8'h47; B = 8'h84; #100;
A = 8'h47; B = 8'h85; #100;
A = 8'h47; B = 8'h86; #100;
A = 8'h47; B = 8'h87; #100;
A = 8'h47; B = 8'h88; #100;
A = 8'h47; B = 8'h89; #100;
A = 8'h47; B = 8'h8A; #100;
A = 8'h47; B = 8'h8B; #100;
A = 8'h47; B = 8'h8C; #100;
A = 8'h47; B = 8'h8D; #100;
A = 8'h47; B = 8'h8E; #100;
A = 8'h47; B = 8'h8F; #100;
A = 8'h47; B = 8'h90; #100;
A = 8'h47; B = 8'h91; #100;
A = 8'h47; B = 8'h92; #100;
A = 8'h47; B = 8'h93; #100;
A = 8'h47; B = 8'h94; #100;
A = 8'h47; B = 8'h95; #100;
A = 8'h47; B = 8'h96; #100;
A = 8'h47; B = 8'h97; #100;
A = 8'h47; B = 8'h98; #100;
A = 8'h47; B = 8'h99; #100;
A = 8'h47; B = 8'h9A; #100;
A = 8'h47; B = 8'h9B; #100;
A = 8'h47; B = 8'h9C; #100;
A = 8'h47; B = 8'h9D; #100;
A = 8'h47; B = 8'h9E; #100;
A = 8'h47; B = 8'h9F; #100;
A = 8'h47; B = 8'hA0; #100;
A = 8'h47; B = 8'hA1; #100;
A = 8'h47; B = 8'hA2; #100;
A = 8'h47; B = 8'hA3; #100;
A = 8'h47; B = 8'hA4; #100;
A = 8'h47; B = 8'hA5; #100;
A = 8'h47; B = 8'hA6; #100;
A = 8'h47; B = 8'hA7; #100;
A = 8'h47; B = 8'hA8; #100;
A = 8'h47; B = 8'hA9; #100;
A = 8'h47; B = 8'hAA; #100;
A = 8'h47; B = 8'hAB; #100;
A = 8'h47; B = 8'hAC; #100;
A = 8'h47; B = 8'hAD; #100;
A = 8'h47; B = 8'hAE; #100;
A = 8'h47; B = 8'hAF; #100;
A = 8'h47; B = 8'hB0; #100;
A = 8'h47; B = 8'hB1; #100;
A = 8'h47; B = 8'hB2; #100;
A = 8'h47; B = 8'hB3; #100;
A = 8'h47; B = 8'hB4; #100;
A = 8'h47; B = 8'hB5; #100;
A = 8'h47; B = 8'hB6; #100;
A = 8'h47; B = 8'hB7; #100;
A = 8'h47; B = 8'hB8; #100;
A = 8'h47; B = 8'hB9; #100;
A = 8'h47; B = 8'hBA; #100;
A = 8'h47; B = 8'hBB; #100;
A = 8'h47; B = 8'hBC; #100;
A = 8'h47; B = 8'hBD; #100;
A = 8'h47; B = 8'hBE; #100;
A = 8'h47; B = 8'hBF; #100;
A = 8'h47; B = 8'hC0; #100;
A = 8'h47; B = 8'hC1; #100;
A = 8'h47; B = 8'hC2; #100;
A = 8'h47; B = 8'hC3; #100;
A = 8'h47; B = 8'hC4; #100;
A = 8'h47; B = 8'hC5; #100;
A = 8'h47; B = 8'hC6; #100;
A = 8'h47; B = 8'hC7; #100;
A = 8'h47; B = 8'hC8; #100;
A = 8'h47; B = 8'hC9; #100;
A = 8'h47; B = 8'hCA; #100;
A = 8'h47; B = 8'hCB; #100;
A = 8'h47; B = 8'hCC; #100;
A = 8'h47; B = 8'hCD; #100;
A = 8'h47; B = 8'hCE; #100;
A = 8'h47; B = 8'hCF; #100;
A = 8'h47; B = 8'hD0; #100;
A = 8'h47; B = 8'hD1; #100;
A = 8'h47; B = 8'hD2; #100;
A = 8'h47; B = 8'hD3; #100;
A = 8'h47; B = 8'hD4; #100;
A = 8'h47; B = 8'hD5; #100;
A = 8'h47; B = 8'hD6; #100;
A = 8'h47; B = 8'hD7; #100;
A = 8'h47; B = 8'hD8; #100;
A = 8'h47; B = 8'hD9; #100;
A = 8'h47; B = 8'hDA; #100;
A = 8'h47; B = 8'hDB; #100;
A = 8'h47; B = 8'hDC; #100;
A = 8'h47; B = 8'hDD; #100;
A = 8'h47; B = 8'hDE; #100;
A = 8'h47; B = 8'hDF; #100;
A = 8'h47; B = 8'hE0; #100;
A = 8'h47; B = 8'hE1; #100;
A = 8'h47; B = 8'hE2; #100;
A = 8'h47; B = 8'hE3; #100;
A = 8'h47; B = 8'hE4; #100;
A = 8'h47; B = 8'hE5; #100;
A = 8'h47; B = 8'hE6; #100;
A = 8'h47; B = 8'hE7; #100;
A = 8'h47; B = 8'hE8; #100;
A = 8'h47; B = 8'hE9; #100;
A = 8'h47; B = 8'hEA; #100;
A = 8'h47; B = 8'hEB; #100;
A = 8'h47; B = 8'hEC; #100;
A = 8'h47; B = 8'hED; #100;
A = 8'h47; B = 8'hEE; #100;
A = 8'h47; B = 8'hEF; #100;
A = 8'h47; B = 8'hF0; #100;
A = 8'h47; B = 8'hF1; #100;
A = 8'h47; B = 8'hF2; #100;
A = 8'h47; B = 8'hF3; #100;
A = 8'h47; B = 8'hF4; #100;
A = 8'h47; B = 8'hF5; #100;
A = 8'h47; B = 8'hF6; #100;
A = 8'h47; B = 8'hF7; #100;
A = 8'h47; B = 8'hF8; #100;
A = 8'h47; B = 8'hF9; #100;
A = 8'h47; B = 8'hFA; #100;
A = 8'h47; B = 8'hFB; #100;
A = 8'h47; B = 8'hFC; #100;
A = 8'h47; B = 8'hFD; #100;
A = 8'h47; B = 8'hFE; #100;
A = 8'h47; B = 8'hFF; #100;
A = 8'h48; B = 8'h0; #100;
A = 8'h48; B = 8'h1; #100;
A = 8'h48; B = 8'h2; #100;
A = 8'h48; B = 8'h3; #100;
A = 8'h48; B = 8'h4; #100;
A = 8'h48; B = 8'h5; #100;
A = 8'h48; B = 8'h6; #100;
A = 8'h48; B = 8'h7; #100;
A = 8'h48; B = 8'h8; #100;
A = 8'h48; B = 8'h9; #100;
A = 8'h48; B = 8'hA; #100;
A = 8'h48; B = 8'hB; #100;
A = 8'h48; B = 8'hC; #100;
A = 8'h48; B = 8'hD; #100;
A = 8'h48; B = 8'hE; #100;
A = 8'h48; B = 8'hF; #100;
A = 8'h48; B = 8'h10; #100;
A = 8'h48; B = 8'h11; #100;
A = 8'h48; B = 8'h12; #100;
A = 8'h48; B = 8'h13; #100;
A = 8'h48; B = 8'h14; #100;
A = 8'h48; B = 8'h15; #100;
A = 8'h48; B = 8'h16; #100;
A = 8'h48; B = 8'h17; #100;
A = 8'h48; B = 8'h18; #100;
A = 8'h48; B = 8'h19; #100;
A = 8'h48; B = 8'h1A; #100;
A = 8'h48; B = 8'h1B; #100;
A = 8'h48; B = 8'h1C; #100;
A = 8'h48; B = 8'h1D; #100;
A = 8'h48; B = 8'h1E; #100;
A = 8'h48; B = 8'h1F; #100;
A = 8'h48; B = 8'h20; #100;
A = 8'h48; B = 8'h21; #100;
A = 8'h48; B = 8'h22; #100;
A = 8'h48; B = 8'h23; #100;
A = 8'h48; B = 8'h24; #100;
A = 8'h48; B = 8'h25; #100;
A = 8'h48; B = 8'h26; #100;
A = 8'h48; B = 8'h27; #100;
A = 8'h48; B = 8'h28; #100;
A = 8'h48; B = 8'h29; #100;
A = 8'h48; B = 8'h2A; #100;
A = 8'h48; B = 8'h2B; #100;
A = 8'h48; B = 8'h2C; #100;
A = 8'h48; B = 8'h2D; #100;
A = 8'h48; B = 8'h2E; #100;
A = 8'h48; B = 8'h2F; #100;
A = 8'h48; B = 8'h30; #100;
A = 8'h48; B = 8'h31; #100;
A = 8'h48; B = 8'h32; #100;
A = 8'h48; B = 8'h33; #100;
A = 8'h48; B = 8'h34; #100;
A = 8'h48; B = 8'h35; #100;
A = 8'h48; B = 8'h36; #100;
A = 8'h48; B = 8'h37; #100;
A = 8'h48; B = 8'h38; #100;
A = 8'h48; B = 8'h39; #100;
A = 8'h48; B = 8'h3A; #100;
A = 8'h48; B = 8'h3B; #100;
A = 8'h48; B = 8'h3C; #100;
A = 8'h48; B = 8'h3D; #100;
A = 8'h48; B = 8'h3E; #100;
A = 8'h48; B = 8'h3F; #100;
A = 8'h48; B = 8'h40; #100;
A = 8'h48; B = 8'h41; #100;
A = 8'h48; B = 8'h42; #100;
A = 8'h48; B = 8'h43; #100;
A = 8'h48; B = 8'h44; #100;
A = 8'h48; B = 8'h45; #100;
A = 8'h48; B = 8'h46; #100;
A = 8'h48; B = 8'h47; #100;
A = 8'h48; B = 8'h48; #100;
A = 8'h48; B = 8'h49; #100;
A = 8'h48; B = 8'h4A; #100;
A = 8'h48; B = 8'h4B; #100;
A = 8'h48; B = 8'h4C; #100;
A = 8'h48; B = 8'h4D; #100;
A = 8'h48; B = 8'h4E; #100;
A = 8'h48; B = 8'h4F; #100;
A = 8'h48; B = 8'h50; #100;
A = 8'h48; B = 8'h51; #100;
A = 8'h48; B = 8'h52; #100;
A = 8'h48; B = 8'h53; #100;
A = 8'h48; B = 8'h54; #100;
A = 8'h48; B = 8'h55; #100;
A = 8'h48; B = 8'h56; #100;
A = 8'h48; B = 8'h57; #100;
A = 8'h48; B = 8'h58; #100;
A = 8'h48; B = 8'h59; #100;
A = 8'h48; B = 8'h5A; #100;
A = 8'h48; B = 8'h5B; #100;
A = 8'h48; B = 8'h5C; #100;
A = 8'h48; B = 8'h5D; #100;
A = 8'h48; B = 8'h5E; #100;
A = 8'h48; B = 8'h5F; #100;
A = 8'h48; B = 8'h60; #100;
A = 8'h48; B = 8'h61; #100;
A = 8'h48; B = 8'h62; #100;
A = 8'h48; B = 8'h63; #100;
A = 8'h48; B = 8'h64; #100;
A = 8'h48; B = 8'h65; #100;
A = 8'h48; B = 8'h66; #100;
A = 8'h48; B = 8'h67; #100;
A = 8'h48; B = 8'h68; #100;
A = 8'h48; B = 8'h69; #100;
A = 8'h48; B = 8'h6A; #100;
A = 8'h48; B = 8'h6B; #100;
A = 8'h48; B = 8'h6C; #100;
A = 8'h48; B = 8'h6D; #100;
A = 8'h48; B = 8'h6E; #100;
A = 8'h48; B = 8'h6F; #100;
A = 8'h48; B = 8'h70; #100;
A = 8'h48; B = 8'h71; #100;
A = 8'h48; B = 8'h72; #100;
A = 8'h48; B = 8'h73; #100;
A = 8'h48; B = 8'h74; #100;
A = 8'h48; B = 8'h75; #100;
A = 8'h48; B = 8'h76; #100;
A = 8'h48; B = 8'h77; #100;
A = 8'h48; B = 8'h78; #100;
A = 8'h48; B = 8'h79; #100;
A = 8'h48; B = 8'h7A; #100;
A = 8'h48; B = 8'h7B; #100;
A = 8'h48; B = 8'h7C; #100;
A = 8'h48; B = 8'h7D; #100;
A = 8'h48; B = 8'h7E; #100;
A = 8'h48; B = 8'h7F; #100;
A = 8'h48; B = 8'h80; #100;
A = 8'h48; B = 8'h81; #100;
A = 8'h48; B = 8'h82; #100;
A = 8'h48; B = 8'h83; #100;
A = 8'h48; B = 8'h84; #100;
A = 8'h48; B = 8'h85; #100;
A = 8'h48; B = 8'h86; #100;
A = 8'h48; B = 8'h87; #100;
A = 8'h48; B = 8'h88; #100;
A = 8'h48; B = 8'h89; #100;
A = 8'h48; B = 8'h8A; #100;
A = 8'h48; B = 8'h8B; #100;
A = 8'h48; B = 8'h8C; #100;
A = 8'h48; B = 8'h8D; #100;
A = 8'h48; B = 8'h8E; #100;
A = 8'h48; B = 8'h8F; #100;
A = 8'h48; B = 8'h90; #100;
A = 8'h48; B = 8'h91; #100;
A = 8'h48; B = 8'h92; #100;
A = 8'h48; B = 8'h93; #100;
A = 8'h48; B = 8'h94; #100;
A = 8'h48; B = 8'h95; #100;
A = 8'h48; B = 8'h96; #100;
A = 8'h48; B = 8'h97; #100;
A = 8'h48; B = 8'h98; #100;
A = 8'h48; B = 8'h99; #100;
A = 8'h48; B = 8'h9A; #100;
A = 8'h48; B = 8'h9B; #100;
A = 8'h48; B = 8'h9C; #100;
A = 8'h48; B = 8'h9D; #100;
A = 8'h48; B = 8'h9E; #100;
A = 8'h48; B = 8'h9F; #100;
A = 8'h48; B = 8'hA0; #100;
A = 8'h48; B = 8'hA1; #100;
A = 8'h48; B = 8'hA2; #100;
A = 8'h48; B = 8'hA3; #100;
A = 8'h48; B = 8'hA4; #100;
A = 8'h48; B = 8'hA5; #100;
A = 8'h48; B = 8'hA6; #100;
A = 8'h48; B = 8'hA7; #100;
A = 8'h48; B = 8'hA8; #100;
A = 8'h48; B = 8'hA9; #100;
A = 8'h48; B = 8'hAA; #100;
A = 8'h48; B = 8'hAB; #100;
A = 8'h48; B = 8'hAC; #100;
A = 8'h48; B = 8'hAD; #100;
A = 8'h48; B = 8'hAE; #100;
A = 8'h48; B = 8'hAF; #100;
A = 8'h48; B = 8'hB0; #100;
A = 8'h48; B = 8'hB1; #100;
A = 8'h48; B = 8'hB2; #100;
A = 8'h48; B = 8'hB3; #100;
A = 8'h48; B = 8'hB4; #100;
A = 8'h48; B = 8'hB5; #100;
A = 8'h48; B = 8'hB6; #100;
A = 8'h48; B = 8'hB7; #100;
A = 8'h48; B = 8'hB8; #100;
A = 8'h48; B = 8'hB9; #100;
A = 8'h48; B = 8'hBA; #100;
A = 8'h48; B = 8'hBB; #100;
A = 8'h48; B = 8'hBC; #100;
A = 8'h48; B = 8'hBD; #100;
A = 8'h48; B = 8'hBE; #100;
A = 8'h48; B = 8'hBF; #100;
A = 8'h48; B = 8'hC0; #100;
A = 8'h48; B = 8'hC1; #100;
A = 8'h48; B = 8'hC2; #100;
A = 8'h48; B = 8'hC3; #100;
A = 8'h48; B = 8'hC4; #100;
A = 8'h48; B = 8'hC5; #100;
A = 8'h48; B = 8'hC6; #100;
A = 8'h48; B = 8'hC7; #100;
A = 8'h48; B = 8'hC8; #100;
A = 8'h48; B = 8'hC9; #100;
A = 8'h48; B = 8'hCA; #100;
A = 8'h48; B = 8'hCB; #100;
A = 8'h48; B = 8'hCC; #100;
A = 8'h48; B = 8'hCD; #100;
A = 8'h48; B = 8'hCE; #100;
A = 8'h48; B = 8'hCF; #100;
A = 8'h48; B = 8'hD0; #100;
A = 8'h48; B = 8'hD1; #100;
A = 8'h48; B = 8'hD2; #100;
A = 8'h48; B = 8'hD3; #100;
A = 8'h48; B = 8'hD4; #100;
A = 8'h48; B = 8'hD5; #100;
A = 8'h48; B = 8'hD6; #100;
A = 8'h48; B = 8'hD7; #100;
A = 8'h48; B = 8'hD8; #100;
A = 8'h48; B = 8'hD9; #100;
A = 8'h48; B = 8'hDA; #100;
A = 8'h48; B = 8'hDB; #100;
A = 8'h48; B = 8'hDC; #100;
A = 8'h48; B = 8'hDD; #100;
A = 8'h48; B = 8'hDE; #100;
A = 8'h48; B = 8'hDF; #100;
A = 8'h48; B = 8'hE0; #100;
A = 8'h48; B = 8'hE1; #100;
A = 8'h48; B = 8'hE2; #100;
A = 8'h48; B = 8'hE3; #100;
A = 8'h48; B = 8'hE4; #100;
A = 8'h48; B = 8'hE5; #100;
A = 8'h48; B = 8'hE6; #100;
A = 8'h48; B = 8'hE7; #100;
A = 8'h48; B = 8'hE8; #100;
A = 8'h48; B = 8'hE9; #100;
A = 8'h48; B = 8'hEA; #100;
A = 8'h48; B = 8'hEB; #100;
A = 8'h48; B = 8'hEC; #100;
A = 8'h48; B = 8'hED; #100;
A = 8'h48; B = 8'hEE; #100;
A = 8'h48; B = 8'hEF; #100;
A = 8'h48; B = 8'hF0; #100;
A = 8'h48; B = 8'hF1; #100;
A = 8'h48; B = 8'hF2; #100;
A = 8'h48; B = 8'hF3; #100;
A = 8'h48; B = 8'hF4; #100;
A = 8'h48; B = 8'hF5; #100;
A = 8'h48; B = 8'hF6; #100;
A = 8'h48; B = 8'hF7; #100;
A = 8'h48; B = 8'hF8; #100;
A = 8'h48; B = 8'hF9; #100;
A = 8'h48; B = 8'hFA; #100;
A = 8'h48; B = 8'hFB; #100;
A = 8'h48; B = 8'hFC; #100;
A = 8'h48; B = 8'hFD; #100;
A = 8'h48; B = 8'hFE; #100;
A = 8'h48; B = 8'hFF; #100;
A = 8'h49; B = 8'h0; #100;
A = 8'h49; B = 8'h1; #100;
A = 8'h49; B = 8'h2; #100;
A = 8'h49; B = 8'h3; #100;
A = 8'h49; B = 8'h4; #100;
A = 8'h49; B = 8'h5; #100;
A = 8'h49; B = 8'h6; #100;
A = 8'h49; B = 8'h7; #100;
A = 8'h49; B = 8'h8; #100;
A = 8'h49; B = 8'h9; #100;
A = 8'h49; B = 8'hA; #100;
A = 8'h49; B = 8'hB; #100;
A = 8'h49; B = 8'hC; #100;
A = 8'h49; B = 8'hD; #100;
A = 8'h49; B = 8'hE; #100;
A = 8'h49; B = 8'hF; #100;
A = 8'h49; B = 8'h10; #100;
A = 8'h49; B = 8'h11; #100;
A = 8'h49; B = 8'h12; #100;
A = 8'h49; B = 8'h13; #100;
A = 8'h49; B = 8'h14; #100;
A = 8'h49; B = 8'h15; #100;
A = 8'h49; B = 8'h16; #100;
A = 8'h49; B = 8'h17; #100;
A = 8'h49; B = 8'h18; #100;
A = 8'h49; B = 8'h19; #100;
A = 8'h49; B = 8'h1A; #100;
A = 8'h49; B = 8'h1B; #100;
A = 8'h49; B = 8'h1C; #100;
A = 8'h49; B = 8'h1D; #100;
A = 8'h49; B = 8'h1E; #100;
A = 8'h49; B = 8'h1F; #100;
A = 8'h49; B = 8'h20; #100;
A = 8'h49; B = 8'h21; #100;
A = 8'h49; B = 8'h22; #100;
A = 8'h49; B = 8'h23; #100;
A = 8'h49; B = 8'h24; #100;
A = 8'h49; B = 8'h25; #100;
A = 8'h49; B = 8'h26; #100;
A = 8'h49; B = 8'h27; #100;
A = 8'h49; B = 8'h28; #100;
A = 8'h49; B = 8'h29; #100;
A = 8'h49; B = 8'h2A; #100;
A = 8'h49; B = 8'h2B; #100;
A = 8'h49; B = 8'h2C; #100;
A = 8'h49; B = 8'h2D; #100;
A = 8'h49; B = 8'h2E; #100;
A = 8'h49; B = 8'h2F; #100;
A = 8'h49; B = 8'h30; #100;
A = 8'h49; B = 8'h31; #100;
A = 8'h49; B = 8'h32; #100;
A = 8'h49; B = 8'h33; #100;
A = 8'h49; B = 8'h34; #100;
A = 8'h49; B = 8'h35; #100;
A = 8'h49; B = 8'h36; #100;
A = 8'h49; B = 8'h37; #100;
A = 8'h49; B = 8'h38; #100;
A = 8'h49; B = 8'h39; #100;
A = 8'h49; B = 8'h3A; #100;
A = 8'h49; B = 8'h3B; #100;
A = 8'h49; B = 8'h3C; #100;
A = 8'h49; B = 8'h3D; #100;
A = 8'h49; B = 8'h3E; #100;
A = 8'h49; B = 8'h3F; #100;
A = 8'h49; B = 8'h40; #100;
A = 8'h49; B = 8'h41; #100;
A = 8'h49; B = 8'h42; #100;
A = 8'h49; B = 8'h43; #100;
A = 8'h49; B = 8'h44; #100;
A = 8'h49; B = 8'h45; #100;
A = 8'h49; B = 8'h46; #100;
A = 8'h49; B = 8'h47; #100;
A = 8'h49; B = 8'h48; #100;
A = 8'h49; B = 8'h49; #100;
A = 8'h49; B = 8'h4A; #100;
A = 8'h49; B = 8'h4B; #100;
A = 8'h49; B = 8'h4C; #100;
A = 8'h49; B = 8'h4D; #100;
A = 8'h49; B = 8'h4E; #100;
A = 8'h49; B = 8'h4F; #100;
A = 8'h49; B = 8'h50; #100;
A = 8'h49; B = 8'h51; #100;
A = 8'h49; B = 8'h52; #100;
A = 8'h49; B = 8'h53; #100;
A = 8'h49; B = 8'h54; #100;
A = 8'h49; B = 8'h55; #100;
A = 8'h49; B = 8'h56; #100;
A = 8'h49; B = 8'h57; #100;
A = 8'h49; B = 8'h58; #100;
A = 8'h49; B = 8'h59; #100;
A = 8'h49; B = 8'h5A; #100;
A = 8'h49; B = 8'h5B; #100;
A = 8'h49; B = 8'h5C; #100;
A = 8'h49; B = 8'h5D; #100;
A = 8'h49; B = 8'h5E; #100;
A = 8'h49; B = 8'h5F; #100;
A = 8'h49; B = 8'h60; #100;
A = 8'h49; B = 8'h61; #100;
A = 8'h49; B = 8'h62; #100;
A = 8'h49; B = 8'h63; #100;
A = 8'h49; B = 8'h64; #100;
A = 8'h49; B = 8'h65; #100;
A = 8'h49; B = 8'h66; #100;
A = 8'h49; B = 8'h67; #100;
A = 8'h49; B = 8'h68; #100;
A = 8'h49; B = 8'h69; #100;
A = 8'h49; B = 8'h6A; #100;
A = 8'h49; B = 8'h6B; #100;
A = 8'h49; B = 8'h6C; #100;
A = 8'h49; B = 8'h6D; #100;
A = 8'h49; B = 8'h6E; #100;
A = 8'h49; B = 8'h6F; #100;
A = 8'h49; B = 8'h70; #100;
A = 8'h49; B = 8'h71; #100;
A = 8'h49; B = 8'h72; #100;
A = 8'h49; B = 8'h73; #100;
A = 8'h49; B = 8'h74; #100;
A = 8'h49; B = 8'h75; #100;
A = 8'h49; B = 8'h76; #100;
A = 8'h49; B = 8'h77; #100;
A = 8'h49; B = 8'h78; #100;
A = 8'h49; B = 8'h79; #100;
A = 8'h49; B = 8'h7A; #100;
A = 8'h49; B = 8'h7B; #100;
A = 8'h49; B = 8'h7C; #100;
A = 8'h49; B = 8'h7D; #100;
A = 8'h49; B = 8'h7E; #100;
A = 8'h49; B = 8'h7F; #100;
A = 8'h49; B = 8'h80; #100;
A = 8'h49; B = 8'h81; #100;
A = 8'h49; B = 8'h82; #100;
A = 8'h49; B = 8'h83; #100;
A = 8'h49; B = 8'h84; #100;
A = 8'h49; B = 8'h85; #100;
A = 8'h49; B = 8'h86; #100;
A = 8'h49; B = 8'h87; #100;
A = 8'h49; B = 8'h88; #100;
A = 8'h49; B = 8'h89; #100;
A = 8'h49; B = 8'h8A; #100;
A = 8'h49; B = 8'h8B; #100;
A = 8'h49; B = 8'h8C; #100;
A = 8'h49; B = 8'h8D; #100;
A = 8'h49; B = 8'h8E; #100;
A = 8'h49; B = 8'h8F; #100;
A = 8'h49; B = 8'h90; #100;
A = 8'h49; B = 8'h91; #100;
A = 8'h49; B = 8'h92; #100;
A = 8'h49; B = 8'h93; #100;
A = 8'h49; B = 8'h94; #100;
A = 8'h49; B = 8'h95; #100;
A = 8'h49; B = 8'h96; #100;
A = 8'h49; B = 8'h97; #100;
A = 8'h49; B = 8'h98; #100;
A = 8'h49; B = 8'h99; #100;
A = 8'h49; B = 8'h9A; #100;
A = 8'h49; B = 8'h9B; #100;
A = 8'h49; B = 8'h9C; #100;
A = 8'h49; B = 8'h9D; #100;
A = 8'h49; B = 8'h9E; #100;
A = 8'h49; B = 8'h9F; #100;
A = 8'h49; B = 8'hA0; #100;
A = 8'h49; B = 8'hA1; #100;
A = 8'h49; B = 8'hA2; #100;
A = 8'h49; B = 8'hA3; #100;
A = 8'h49; B = 8'hA4; #100;
A = 8'h49; B = 8'hA5; #100;
A = 8'h49; B = 8'hA6; #100;
A = 8'h49; B = 8'hA7; #100;
A = 8'h49; B = 8'hA8; #100;
A = 8'h49; B = 8'hA9; #100;
A = 8'h49; B = 8'hAA; #100;
A = 8'h49; B = 8'hAB; #100;
A = 8'h49; B = 8'hAC; #100;
A = 8'h49; B = 8'hAD; #100;
A = 8'h49; B = 8'hAE; #100;
A = 8'h49; B = 8'hAF; #100;
A = 8'h49; B = 8'hB0; #100;
A = 8'h49; B = 8'hB1; #100;
A = 8'h49; B = 8'hB2; #100;
A = 8'h49; B = 8'hB3; #100;
A = 8'h49; B = 8'hB4; #100;
A = 8'h49; B = 8'hB5; #100;
A = 8'h49; B = 8'hB6; #100;
A = 8'h49; B = 8'hB7; #100;
A = 8'h49; B = 8'hB8; #100;
A = 8'h49; B = 8'hB9; #100;
A = 8'h49; B = 8'hBA; #100;
A = 8'h49; B = 8'hBB; #100;
A = 8'h49; B = 8'hBC; #100;
A = 8'h49; B = 8'hBD; #100;
A = 8'h49; B = 8'hBE; #100;
A = 8'h49; B = 8'hBF; #100;
A = 8'h49; B = 8'hC0; #100;
A = 8'h49; B = 8'hC1; #100;
A = 8'h49; B = 8'hC2; #100;
A = 8'h49; B = 8'hC3; #100;
A = 8'h49; B = 8'hC4; #100;
A = 8'h49; B = 8'hC5; #100;
A = 8'h49; B = 8'hC6; #100;
A = 8'h49; B = 8'hC7; #100;
A = 8'h49; B = 8'hC8; #100;
A = 8'h49; B = 8'hC9; #100;
A = 8'h49; B = 8'hCA; #100;
A = 8'h49; B = 8'hCB; #100;
A = 8'h49; B = 8'hCC; #100;
A = 8'h49; B = 8'hCD; #100;
A = 8'h49; B = 8'hCE; #100;
A = 8'h49; B = 8'hCF; #100;
A = 8'h49; B = 8'hD0; #100;
A = 8'h49; B = 8'hD1; #100;
A = 8'h49; B = 8'hD2; #100;
A = 8'h49; B = 8'hD3; #100;
A = 8'h49; B = 8'hD4; #100;
A = 8'h49; B = 8'hD5; #100;
A = 8'h49; B = 8'hD6; #100;
A = 8'h49; B = 8'hD7; #100;
A = 8'h49; B = 8'hD8; #100;
A = 8'h49; B = 8'hD9; #100;
A = 8'h49; B = 8'hDA; #100;
A = 8'h49; B = 8'hDB; #100;
A = 8'h49; B = 8'hDC; #100;
A = 8'h49; B = 8'hDD; #100;
A = 8'h49; B = 8'hDE; #100;
A = 8'h49; B = 8'hDF; #100;
A = 8'h49; B = 8'hE0; #100;
A = 8'h49; B = 8'hE1; #100;
A = 8'h49; B = 8'hE2; #100;
A = 8'h49; B = 8'hE3; #100;
A = 8'h49; B = 8'hE4; #100;
A = 8'h49; B = 8'hE5; #100;
A = 8'h49; B = 8'hE6; #100;
A = 8'h49; B = 8'hE7; #100;
A = 8'h49; B = 8'hE8; #100;
A = 8'h49; B = 8'hE9; #100;
A = 8'h49; B = 8'hEA; #100;
A = 8'h49; B = 8'hEB; #100;
A = 8'h49; B = 8'hEC; #100;
A = 8'h49; B = 8'hED; #100;
A = 8'h49; B = 8'hEE; #100;
A = 8'h49; B = 8'hEF; #100;
A = 8'h49; B = 8'hF0; #100;
A = 8'h49; B = 8'hF1; #100;
A = 8'h49; B = 8'hF2; #100;
A = 8'h49; B = 8'hF3; #100;
A = 8'h49; B = 8'hF4; #100;
A = 8'h49; B = 8'hF5; #100;
A = 8'h49; B = 8'hF6; #100;
A = 8'h49; B = 8'hF7; #100;
A = 8'h49; B = 8'hF8; #100;
A = 8'h49; B = 8'hF9; #100;
A = 8'h49; B = 8'hFA; #100;
A = 8'h49; B = 8'hFB; #100;
A = 8'h49; B = 8'hFC; #100;
A = 8'h49; B = 8'hFD; #100;
A = 8'h49; B = 8'hFE; #100;
A = 8'h49; B = 8'hFF; #100;
A = 8'h4A; B = 8'h0; #100;
A = 8'h4A; B = 8'h1; #100;
A = 8'h4A; B = 8'h2; #100;
A = 8'h4A; B = 8'h3; #100;
A = 8'h4A; B = 8'h4; #100;
A = 8'h4A; B = 8'h5; #100;
A = 8'h4A; B = 8'h6; #100;
A = 8'h4A; B = 8'h7; #100;
A = 8'h4A; B = 8'h8; #100;
A = 8'h4A; B = 8'h9; #100;
A = 8'h4A; B = 8'hA; #100;
A = 8'h4A; B = 8'hB; #100;
A = 8'h4A; B = 8'hC; #100;
A = 8'h4A; B = 8'hD; #100;
A = 8'h4A; B = 8'hE; #100;
A = 8'h4A; B = 8'hF; #100;
A = 8'h4A; B = 8'h10; #100;
A = 8'h4A; B = 8'h11; #100;
A = 8'h4A; B = 8'h12; #100;
A = 8'h4A; B = 8'h13; #100;
A = 8'h4A; B = 8'h14; #100;
A = 8'h4A; B = 8'h15; #100;
A = 8'h4A; B = 8'h16; #100;
A = 8'h4A; B = 8'h17; #100;
A = 8'h4A; B = 8'h18; #100;
A = 8'h4A; B = 8'h19; #100;
A = 8'h4A; B = 8'h1A; #100;
A = 8'h4A; B = 8'h1B; #100;
A = 8'h4A; B = 8'h1C; #100;
A = 8'h4A; B = 8'h1D; #100;
A = 8'h4A; B = 8'h1E; #100;
A = 8'h4A; B = 8'h1F; #100;
A = 8'h4A; B = 8'h20; #100;
A = 8'h4A; B = 8'h21; #100;
A = 8'h4A; B = 8'h22; #100;
A = 8'h4A; B = 8'h23; #100;
A = 8'h4A; B = 8'h24; #100;
A = 8'h4A; B = 8'h25; #100;
A = 8'h4A; B = 8'h26; #100;
A = 8'h4A; B = 8'h27; #100;
A = 8'h4A; B = 8'h28; #100;
A = 8'h4A; B = 8'h29; #100;
A = 8'h4A; B = 8'h2A; #100;
A = 8'h4A; B = 8'h2B; #100;
A = 8'h4A; B = 8'h2C; #100;
A = 8'h4A; B = 8'h2D; #100;
A = 8'h4A; B = 8'h2E; #100;
A = 8'h4A; B = 8'h2F; #100;
A = 8'h4A; B = 8'h30; #100;
A = 8'h4A; B = 8'h31; #100;
A = 8'h4A; B = 8'h32; #100;
A = 8'h4A; B = 8'h33; #100;
A = 8'h4A; B = 8'h34; #100;
A = 8'h4A; B = 8'h35; #100;
A = 8'h4A; B = 8'h36; #100;
A = 8'h4A; B = 8'h37; #100;
A = 8'h4A; B = 8'h38; #100;
A = 8'h4A; B = 8'h39; #100;
A = 8'h4A; B = 8'h3A; #100;
A = 8'h4A; B = 8'h3B; #100;
A = 8'h4A; B = 8'h3C; #100;
A = 8'h4A; B = 8'h3D; #100;
A = 8'h4A; B = 8'h3E; #100;
A = 8'h4A; B = 8'h3F; #100;
A = 8'h4A; B = 8'h40; #100;
A = 8'h4A; B = 8'h41; #100;
A = 8'h4A; B = 8'h42; #100;
A = 8'h4A; B = 8'h43; #100;
A = 8'h4A; B = 8'h44; #100;
A = 8'h4A; B = 8'h45; #100;
A = 8'h4A; B = 8'h46; #100;
A = 8'h4A; B = 8'h47; #100;
A = 8'h4A; B = 8'h48; #100;
A = 8'h4A; B = 8'h49; #100;
A = 8'h4A; B = 8'h4A; #100;
A = 8'h4A; B = 8'h4B; #100;
A = 8'h4A; B = 8'h4C; #100;
A = 8'h4A; B = 8'h4D; #100;
A = 8'h4A; B = 8'h4E; #100;
A = 8'h4A; B = 8'h4F; #100;
A = 8'h4A; B = 8'h50; #100;
A = 8'h4A; B = 8'h51; #100;
A = 8'h4A; B = 8'h52; #100;
A = 8'h4A; B = 8'h53; #100;
A = 8'h4A; B = 8'h54; #100;
A = 8'h4A; B = 8'h55; #100;
A = 8'h4A; B = 8'h56; #100;
A = 8'h4A; B = 8'h57; #100;
A = 8'h4A; B = 8'h58; #100;
A = 8'h4A; B = 8'h59; #100;
A = 8'h4A; B = 8'h5A; #100;
A = 8'h4A; B = 8'h5B; #100;
A = 8'h4A; B = 8'h5C; #100;
A = 8'h4A; B = 8'h5D; #100;
A = 8'h4A; B = 8'h5E; #100;
A = 8'h4A; B = 8'h5F; #100;
A = 8'h4A; B = 8'h60; #100;
A = 8'h4A; B = 8'h61; #100;
A = 8'h4A; B = 8'h62; #100;
A = 8'h4A; B = 8'h63; #100;
A = 8'h4A; B = 8'h64; #100;
A = 8'h4A; B = 8'h65; #100;
A = 8'h4A; B = 8'h66; #100;
A = 8'h4A; B = 8'h67; #100;
A = 8'h4A; B = 8'h68; #100;
A = 8'h4A; B = 8'h69; #100;
A = 8'h4A; B = 8'h6A; #100;
A = 8'h4A; B = 8'h6B; #100;
A = 8'h4A; B = 8'h6C; #100;
A = 8'h4A; B = 8'h6D; #100;
A = 8'h4A; B = 8'h6E; #100;
A = 8'h4A; B = 8'h6F; #100;
A = 8'h4A; B = 8'h70; #100;
A = 8'h4A; B = 8'h71; #100;
A = 8'h4A; B = 8'h72; #100;
A = 8'h4A; B = 8'h73; #100;
A = 8'h4A; B = 8'h74; #100;
A = 8'h4A; B = 8'h75; #100;
A = 8'h4A; B = 8'h76; #100;
A = 8'h4A; B = 8'h77; #100;
A = 8'h4A; B = 8'h78; #100;
A = 8'h4A; B = 8'h79; #100;
A = 8'h4A; B = 8'h7A; #100;
A = 8'h4A; B = 8'h7B; #100;
A = 8'h4A; B = 8'h7C; #100;
A = 8'h4A; B = 8'h7D; #100;
A = 8'h4A; B = 8'h7E; #100;
A = 8'h4A; B = 8'h7F; #100;
A = 8'h4A; B = 8'h80; #100;
A = 8'h4A; B = 8'h81; #100;
A = 8'h4A; B = 8'h82; #100;
A = 8'h4A; B = 8'h83; #100;
A = 8'h4A; B = 8'h84; #100;
A = 8'h4A; B = 8'h85; #100;
A = 8'h4A; B = 8'h86; #100;
A = 8'h4A; B = 8'h87; #100;
A = 8'h4A; B = 8'h88; #100;
A = 8'h4A; B = 8'h89; #100;
A = 8'h4A; B = 8'h8A; #100;
A = 8'h4A; B = 8'h8B; #100;
A = 8'h4A; B = 8'h8C; #100;
A = 8'h4A; B = 8'h8D; #100;
A = 8'h4A; B = 8'h8E; #100;
A = 8'h4A; B = 8'h8F; #100;
A = 8'h4A; B = 8'h90; #100;
A = 8'h4A; B = 8'h91; #100;
A = 8'h4A; B = 8'h92; #100;
A = 8'h4A; B = 8'h93; #100;
A = 8'h4A; B = 8'h94; #100;
A = 8'h4A; B = 8'h95; #100;
A = 8'h4A; B = 8'h96; #100;
A = 8'h4A; B = 8'h97; #100;
A = 8'h4A; B = 8'h98; #100;
A = 8'h4A; B = 8'h99; #100;
A = 8'h4A; B = 8'h9A; #100;
A = 8'h4A; B = 8'h9B; #100;
A = 8'h4A; B = 8'h9C; #100;
A = 8'h4A; B = 8'h9D; #100;
A = 8'h4A; B = 8'h9E; #100;
A = 8'h4A; B = 8'h9F; #100;
A = 8'h4A; B = 8'hA0; #100;
A = 8'h4A; B = 8'hA1; #100;
A = 8'h4A; B = 8'hA2; #100;
A = 8'h4A; B = 8'hA3; #100;
A = 8'h4A; B = 8'hA4; #100;
A = 8'h4A; B = 8'hA5; #100;
A = 8'h4A; B = 8'hA6; #100;
A = 8'h4A; B = 8'hA7; #100;
A = 8'h4A; B = 8'hA8; #100;
A = 8'h4A; B = 8'hA9; #100;
A = 8'h4A; B = 8'hAA; #100;
A = 8'h4A; B = 8'hAB; #100;
A = 8'h4A; B = 8'hAC; #100;
A = 8'h4A; B = 8'hAD; #100;
A = 8'h4A; B = 8'hAE; #100;
A = 8'h4A; B = 8'hAF; #100;
A = 8'h4A; B = 8'hB0; #100;
A = 8'h4A; B = 8'hB1; #100;
A = 8'h4A; B = 8'hB2; #100;
A = 8'h4A; B = 8'hB3; #100;
A = 8'h4A; B = 8'hB4; #100;
A = 8'h4A; B = 8'hB5; #100;
A = 8'h4A; B = 8'hB6; #100;
A = 8'h4A; B = 8'hB7; #100;
A = 8'h4A; B = 8'hB8; #100;
A = 8'h4A; B = 8'hB9; #100;
A = 8'h4A; B = 8'hBA; #100;
A = 8'h4A; B = 8'hBB; #100;
A = 8'h4A; B = 8'hBC; #100;
A = 8'h4A; B = 8'hBD; #100;
A = 8'h4A; B = 8'hBE; #100;
A = 8'h4A; B = 8'hBF; #100;
A = 8'h4A; B = 8'hC0; #100;
A = 8'h4A; B = 8'hC1; #100;
A = 8'h4A; B = 8'hC2; #100;
A = 8'h4A; B = 8'hC3; #100;
A = 8'h4A; B = 8'hC4; #100;
A = 8'h4A; B = 8'hC5; #100;
A = 8'h4A; B = 8'hC6; #100;
A = 8'h4A; B = 8'hC7; #100;
A = 8'h4A; B = 8'hC8; #100;
A = 8'h4A; B = 8'hC9; #100;
A = 8'h4A; B = 8'hCA; #100;
A = 8'h4A; B = 8'hCB; #100;
A = 8'h4A; B = 8'hCC; #100;
A = 8'h4A; B = 8'hCD; #100;
A = 8'h4A; B = 8'hCE; #100;
A = 8'h4A; B = 8'hCF; #100;
A = 8'h4A; B = 8'hD0; #100;
A = 8'h4A; B = 8'hD1; #100;
A = 8'h4A; B = 8'hD2; #100;
A = 8'h4A; B = 8'hD3; #100;
A = 8'h4A; B = 8'hD4; #100;
A = 8'h4A; B = 8'hD5; #100;
A = 8'h4A; B = 8'hD6; #100;
A = 8'h4A; B = 8'hD7; #100;
A = 8'h4A; B = 8'hD8; #100;
A = 8'h4A; B = 8'hD9; #100;
A = 8'h4A; B = 8'hDA; #100;
A = 8'h4A; B = 8'hDB; #100;
A = 8'h4A; B = 8'hDC; #100;
A = 8'h4A; B = 8'hDD; #100;
A = 8'h4A; B = 8'hDE; #100;
A = 8'h4A; B = 8'hDF; #100;
A = 8'h4A; B = 8'hE0; #100;
A = 8'h4A; B = 8'hE1; #100;
A = 8'h4A; B = 8'hE2; #100;
A = 8'h4A; B = 8'hE3; #100;
A = 8'h4A; B = 8'hE4; #100;
A = 8'h4A; B = 8'hE5; #100;
A = 8'h4A; B = 8'hE6; #100;
A = 8'h4A; B = 8'hE7; #100;
A = 8'h4A; B = 8'hE8; #100;
A = 8'h4A; B = 8'hE9; #100;
A = 8'h4A; B = 8'hEA; #100;
A = 8'h4A; B = 8'hEB; #100;
A = 8'h4A; B = 8'hEC; #100;
A = 8'h4A; B = 8'hED; #100;
A = 8'h4A; B = 8'hEE; #100;
A = 8'h4A; B = 8'hEF; #100;
A = 8'h4A; B = 8'hF0; #100;
A = 8'h4A; B = 8'hF1; #100;
A = 8'h4A; B = 8'hF2; #100;
A = 8'h4A; B = 8'hF3; #100;
A = 8'h4A; B = 8'hF4; #100;
A = 8'h4A; B = 8'hF5; #100;
A = 8'h4A; B = 8'hF6; #100;
A = 8'h4A; B = 8'hF7; #100;
A = 8'h4A; B = 8'hF8; #100;
A = 8'h4A; B = 8'hF9; #100;
A = 8'h4A; B = 8'hFA; #100;
A = 8'h4A; B = 8'hFB; #100;
A = 8'h4A; B = 8'hFC; #100;
A = 8'h4A; B = 8'hFD; #100;
A = 8'h4A; B = 8'hFE; #100;
A = 8'h4A; B = 8'hFF; #100;
A = 8'h4B; B = 8'h0; #100;
A = 8'h4B; B = 8'h1; #100;
A = 8'h4B; B = 8'h2; #100;
A = 8'h4B; B = 8'h3; #100;
A = 8'h4B; B = 8'h4; #100;
A = 8'h4B; B = 8'h5; #100;
A = 8'h4B; B = 8'h6; #100;
A = 8'h4B; B = 8'h7; #100;
A = 8'h4B; B = 8'h8; #100;
A = 8'h4B; B = 8'h9; #100;
A = 8'h4B; B = 8'hA; #100;
A = 8'h4B; B = 8'hB; #100;
A = 8'h4B; B = 8'hC; #100;
A = 8'h4B; B = 8'hD; #100;
A = 8'h4B; B = 8'hE; #100;
A = 8'h4B; B = 8'hF; #100;
A = 8'h4B; B = 8'h10; #100;
A = 8'h4B; B = 8'h11; #100;
A = 8'h4B; B = 8'h12; #100;
A = 8'h4B; B = 8'h13; #100;
A = 8'h4B; B = 8'h14; #100;
A = 8'h4B; B = 8'h15; #100;
A = 8'h4B; B = 8'h16; #100;
A = 8'h4B; B = 8'h17; #100;
A = 8'h4B; B = 8'h18; #100;
A = 8'h4B; B = 8'h19; #100;
A = 8'h4B; B = 8'h1A; #100;
A = 8'h4B; B = 8'h1B; #100;
A = 8'h4B; B = 8'h1C; #100;
A = 8'h4B; B = 8'h1D; #100;
A = 8'h4B; B = 8'h1E; #100;
A = 8'h4B; B = 8'h1F; #100;
A = 8'h4B; B = 8'h20; #100;
A = 8'h4B; B = 8'h21; #100;
A = 8'h4B; B = 8'h22; #100;
A = 8'h4B; B = 8'h23; #100;
A = 8'h4B; B = 8'h24; #100;
A = 8'h4B; B = 8'h25; #100;
A = 8'h4B; B = 8'h26; #100;
A = 8'h4B; B = 8'h27; #100;
A = 8'h4B; B = 8'h28; #100;
A = 8'h4B; B = 8'h29; #100;
A = 8'h4B; B = 8'h2A; #100;
A = 8'h4B; B = 8'h2B; #100;
A = 8'h4B; B = 8'h2C; #100;
A = 8'h4B; B = 8'h2D; #100;
A = 8'h4B; B = 8'h2E; #100;
A = 8'h4B; B = 8'h2F; #100;
A = 8'h4B; B = 8'h30; #100;
A = 8'h4B; B = 8'h31; #100;
A = 8'h4B; B = 8'h32; #100;
A = 8'h4B; B = 8'h33; #100;
A = 8'h4B; B = 8'h34; #100;
A = 8'h4B; B = 8'h35; #100;
A = 8'h4B; B = 8'h36; #100;
A = 8'h4B; B = 8'h37; #100;
A = 8'h4B; B = 8'h38; #100;
A = 8'h4B; B = 8'h39; #100;
A = 8'h4B; B = 8'h3A; #100;
A = 8'h4B; B = 8'h3B; #100;
A = 8'h4B; B = 8'h3C; #100;
A = 8'h4B; B = 8'h3D; #100;
A = 8'h4B; B = 8'h3E; #100;
A = 8'h4B; B = 8'h3F; #100;
A = 8'h4B; B = 8'h40; #100;
A = 8'h4B; B = 8'h41; #100;
A = 8'h4B; B = 8'h42; #100;
A = 8'h4B; B = 8'h43; #100;
A = 8'h4B; B = 8'h44; #100;
A = 8'h4B; B = 8'h45; #100;
A = 8'h4B; B = 8'h46; #100;
A = 8'h4B; B = 8'h47; #100;
A = 8'h4B; B = 8'h48; #100;
A = 8'h4B; B = 8'h49; #100;
A = 8'h4B; B = 8'h4A; #100;
A = 8'h4B; B = 8'h4B; #100;
A = 8'h4B; B = 8'h4C; #100;
A = 8'h4B; B = 8'h4D; #100;
A = 8'h4B; B = 8'h4E; #100;
A = 8'h4B; B = 8'h4F; #100;
A = 8'h4B; B = 8'h50; #100;
A = 8'h4B; B = 8'h51; #100;
A = 8'h4B; B = 8'h52; #100;
A = 8'h4B; B = 8'h53; #100;
A = 8'h4B; B = 8'h54; #100;
A = 8'h4B; B = 8'h55; #100;
A = 8'h4B; B = 8'h56; #100;
A = 8'h4B; B = 8'h57; #100;
A = 8'h4B; B = 8'h58; #100;
A = 8'h4B; B = 8'h59; #100;
A = 8'h4B; B = 8'h5A; #100;
A = 8'h4B; B = 8'h5B; #100;
A = 8'h4B; B = 8'h5C; #100;
A = 8'h4B; B = 8'h5D; #100;
A = 8'h4B; B = 8'h5E; #100;
A = 8'h4B; B = 8'h5F; #100;
A = 8'h4B; B = 8'h60; #100;
A = 8'h4B; B = 8'h61; #100;
A = 8'h4B; B = 8'h62; #100;
A = 8'h4B; B = 8'h63; #100;
A = 8'h4B; B = 8'h64; #100;
A = 8'h4B; B = 8'h65; #100;
A = 8'h4B; B = 8'h66; #100;
A = 8'h4B; B = 8'h67; #100;
A = 8'h4B; B = 8'h68; #100;
A = 8'h4B; B = 8'h69; #100;
A = 8'h4B; B = 8'h6A; #100;
A = 8'h4B; B = 8'h6B; #100;
A = 8'h4B; B = 8'h6C; #100;
A = 8'h4B; B = 8'h6D; #100;
A = 8'h4B; B = 8'h6E; #100;
A = 8'h4B; B = 8'h6F; #100;
A = 8'h4B; B = 8'h70; #100;
A = 8'h4B; B = 8'h71; #100;
A = 8'h4B; B = 8'h72; #100;
A = 8'h4B; B = 8'h73; #100;
A = 8'h4B; B = 8'h74; #100;
A = 8'h4B; B = 8'h75; #100;
A = 8'h4B; B = 8'h76; #100;
A = 8'h4B; B = 8'h77; #100;
A = 8'h4B; B = 8'h78; #100;
A = 8'h4B; B = 8'h79; #100;
A = 8'h4B; B = 8'h7A; #100;
A = 8'h4B; B = 8'h7B; #100;
A = 8'h4B; B = 8'h7C; #100;
A = 8'h4B; B = 8'h7D; #100;
A = 8'h4B; B = 8'h7E; #100;
A = 8'h4B; B = 8'h7F; #100;
A = 8'h4B; B = 8'h80; #100;
A = 8'h4B; B = 8'h81; #100;
A = 8'h4B; B = 8'h82; #100;
A = 8'h4B; B = 8'h83; #100;
A = 8'h4B; B = 8'h84; #100;
A = 8'h4B; B = 8'h85; #100;
A = 8'h4B; B = 8'h86; #100;
A = 8'h4B; B = 8'h87; #100;
A = 8'h4B; B = 8'h88; #100;
A = 8'h4B; B = 8'h89; #100;
A = 8'h4B; B = 8'h8A; #100;
A = 8'h4B; B = 8'h8B; #100;
A = 8'h4B; B = 8'h8C; #100;
A = 8'h4B; B = 8'h8D; #100;
A = 8'h4B; B = 8'h8E; #100;
A = 8'h4B; B = 8'h8F; #100;
A = 8'h4B; B = 8'h90; #100;
A = 8'h4B; B = 8'h91; #100;
A = 8'h4B; B = 8'h92; #100;
A = 8'h4B; B = 8'h93; #100;
A = 8'h4B; B = 8'h94; #100;
A = 8'h4B; B = 8'h95; #100;
A = 8'h4B; B = 8'h96; #100;
A = 8'h4B; B = 8'h97; #100;
A = 8'h4B; B = 8'h98; #100;
A = 8'h4B; B = 8'h99; #100;
A = 8'h4B; B = 8'h9A; #100;
A = 8'h4B; B = 8'h9B; #100;
A = 8'h4B; B = 8'h9C; #100;
A = 8'h4B; B = 8'h9D; #100;
A = 8'h4B; B = 8'h9E; #100;
A = 8'h4B; B = 8'h9F; #100;
A = 8'h4B; B = 8'hA0; #100;
A = 8'h4B; B = 8'hA1; #100;
A = 8'h4B; B = 8'hA2; #100;
A = 8'h4B; B = 8'hA3; #100;
A = 8'h4B; B = 8'hA4; #100;
A = 8'h4B; B = 8'hA5; #100;
A = 8'h4B; B = 8'hA6; #100;
A = 8'h4B; B = 8'hA7; #100;
A = 8'h4B; B = 8'hA8; #100;
A = 8'h4B; B = 8'hA9; #100;
A = 8'h4B; B = 8'hAA; #100;
A = 8'h4B; B = 8'hAB; #100;
A = 8'h4B; B = 8'hAC; #100;
A = 8'h4B; B = 8'hAD; #100;
A = 8'h4B; B = 8'hAE; #100;
A = 8'h4B; B = 8'hAF; #100;
A = 8'h4B; B = 8'hB0; #100;
A = 8'h4B; B = 8'hB1; #100;
A = 8'h4B; B = 8'hB2; #100;
A = 8'h4B; B = 8'hB3; #100;
A = 8'h4B; B = 8'hB4; #100;
A = 8'h4B; B = 8'hB5; #100;
A = 8'h4B; B = 8'hB6; #100;
A = 8'h4B; B = 8'hB7; #100;
A = 8'h4B; B = 8'hB8; #100;
A = 8'h4B; B = 8'hB9; #100;
A = 8'h4B; B = 8'hBA; #100;
A = 8'h4B; B = 8'hBB; #100;
A = 8'h4B; B = 8'hBC; #100;
A = 8'h4B; B = 8'hBD; #100;
A = 8'h4B; B = 8'hBE; #100;
A = 8'h4B; B = 8'hBF; #100;
A = 8'h4B; B = 8'hC0; #100;
A = 8'h4B; B = 8'hC1; #100;
A = 8'h4B; B = 8'hC2; #100;
A = 8'h4B; B = 8'hC3; #100;
A = 8'h4B; B = 8'hC4; #100;
A = 8'h4B; B = 8'hC5; #100;
A = 8'h4B; B = 8'hC6; #100;
A = 8'h4B; B = 8'hC7; #100;
A = 8'h4B; B = 8'hC8; #100;
A = 8'h4B; B = 8'hC9; #100;
A = 8'h4B; B = 8'hCA; #100;
A = 8'h4B; B = 8'hCB; #100;
A = 8'h4B; B = 8'hCC; #100;
A = 8'h4B; B = 8'hCD; #100;
A = 8'h4B; B = 8'hCE; #100;
A = 8'h4B; B = 8'hCF; #100;
A = 8'h4B; B = 8'hD0; #100;
A = 8'h4B; B = 8'hD1; #100;
A = 8'h4B; B = 8'hD2; #100;
A = 8'h4B; B = 8'hD3; #100;
A = 8'h4B; B = 8'hD4; #100;
A = 8'h4B; B = 8'hD5; #100;
A = 8'h4B; B = 8'hD6; #100;
A = 8'h4B; B = 8'hD7; #100;
A = 8'h4B; B = 8'hD8; #100;
A = 8'h4B; B = 8'hD9; #100;
A = 8'h4B; B = 8'hDA; #100;
A = 8'h4B; B = 8'hDB; #100;
A = 8'h4B; B = 8'hDC; #100;
A = 8'h4B; B = 8'hDD; #100;
A = 8'h4B; B = 8'hDE; #100;
A = 8'h4B; B = 8'hDF; #100;
A = 8'h4B; B = 8'hE0; #100;
A = 8'h4B; B = 8'hE1; #100;
A = 8'h4B; B = 8'hE2; #100;
A = 8'h4B; B = 8'hE3; #100;
A = 8'h4B; B = 8'hE4; #100;
A = 8'h4B; B = 8'hE5; #100;
A = 8'h4B; B = 8'hE6; #100;
A = 8'h4B; B = 8'hE7; #100;
A = 8'h4B; B = 8'hE8; #100;
A = 8'h4B; B = 8'hE9; #100;
A = 8'h4B; B = 8'hEA; #100;
A = 8'h4B; B = 8'hEB; #100;
A = 8'h4B; B = 8'hEC; #100;
A = 8'h4B; B = 8'hED; #100;
A = 8'h4B; B = 8'hEE; #100;
A = 8'h4B; B = 8'hEF; #100;
A = 8'h4B; B = 8'hF0; #100;
A = 8'h4B; B = 8'hF1; #100;
A = 8'h4B; B = 8'hF2; #100;
A = 8'h4B; B = 8'hF3; #100;
A = 8'h4B; B = 8'hF4; #100;
A = 8'h4B; B = 8'hF5; #100;
A = 8'h4B; B = 8'hF6; #100;
A = 8'h4B; B = 8'hF7; #100;
A = 8'h4B; B = 8'hF8; #100;
A = 8'h4B; B = 8'hF9; #100;
A = 8'h4B; B = 8'hFA; #100;
A = 8'h4B; B = 8'hFB; #100;
A = 8'h4B; B = 8'hFC; #100;
A = 8'h4B; B = 8'hFD; #100;
A = 8'h4B; B = 8'hFE; #100;
A = 8'h4B; B = 8'hFF; #100;
A = 8'h4C; B = 8'h0; #100;
A = 8'h4C; B = 8'h1; #100;
A = 8'h4C; B = 8'h2; #100;
A = 8'h4C; B = 8'h3; #100;
A = 8'h4C; B = 8'h4; #100;
A = 8'h4C; B = 8'h5; #100;
A = 8'h4C; B = 8'h6; #100;
A = 8'h4C; B = 8'h7; #100;
A = 8'h4C; B = 8'h8; #100;
A = 8'h4C; B = 8'h9; #100;
A = 8'h4C; B = 8'hA; #100;
A = 8'h4C; B = 8'hB; #100;
A = 8'h4C; B = 8'hC; #100;
A = 8'h4C; B = 8'hD; #100;
A = 8'h4C; B = 8'hE; #100;
A = 8'h4C; B = 8'hF; #100;
A = 8'h4C; B = 8'h10; #100;
A = 8'h4C; B = 8'h11; #100;
A = 8'h4C; B = 8'h12; #100;
A = 8'h4C; B = 8'h13; #100;
A = 8'h4C; B = 8'h14; #100;
A = 8'h4C; B = 8'h15; #100;
A = 8'h4C; B = 8'h16; #100;
A = 8'h4C; B = 8'h17; #100;
A = 8'h4C; B = 8'h18; #100;
A = 8'h4C; B = 8'h19; #100;
A = 8'h4C; B = 8'h1A; #100;
A = 8'h4C; B = 8'h1B; #100;
A = 8'h4C; B = 8'h1C; #100;
A = 8'h4C; B = 8'h1D; #100;
A = 8'h4C; B = 8'h1E; #100;
A = 8'h4C; B = 8'h1F; #100;
A = 8'h4C; B = 8'h20; #100;
A = 8'h4C; B = 8'h21; #100;
A = 8'h4C; B = 8'h22; #100;
A = 8'h4C; B = 8'h23; #100;
A = 8'h4C; B = 8'h24; #100;
A = 8'h4C; B = 8'h25; #100;
A = 8'h4C; B = 8'h26; #100;
A = 8'h4C; B = 8'h27; #100;
A = 8'h4C; B = 8'h28; #100;
A = 8'h4C; B = 8'h29; #100;
A = 8'h4C; B = 8'h2A; #100;
A = 8'h4C; B = 8'h2B; #100;
A = 8'h4C; B = 8'h2C; #100;
A = 8'h4C; B = 8'h2D; #100;
A = 8'h4C; B = 8'h2E; #100;
A = 8'h4C; B = 8'h2F; #100;
A = 8'h4C; B = 8'h30; #100;
A = 8'h4C; B = 8'h31; #100;
A = 8'h4C; B = 8'h32; #100;
A = 8'h4C; B = 8'h33; #100;
A = 8'h4C; B = 8'h34; #100;
A = 8'h4C; B = 8'h35; #100;
A = 8'h4C; B = 8'h36; #100;
A = 8'h4C; B = 8'h37; #100;
A = 8'h4C; B = 8'h38; #100;
A = 8'h4C; B = 8'h39; #100;
A = 8'h4C; B = 8'h3A; #100;
A = 8'h4C; B = 8'h3B; #100;
A = 8'h4C; B = 8'h3C; #100;
A = 8'h4C; B = 8'h3D; #100;
A = 8'h4C; B = 8'h3E; #100;
A = 8'h4C; B = 8'h3F; #100;
A = 8'h4C; B = 8'h40; #100;
A = 8'h4C; B = 8'h41; #100;
A = 8'h4C; B = 8'h42; #100;
A = 8'h4C; B = 8'h43; #100;
A = 8'h4C; B = 8'h44; #100;
A = 8'h4C; B = 8'h45; #100;
A = 8'h4C; B = 8'h46; #100;
A = 8'h4C; B = 8'h47; #100;
A = 8'h4C; B = 8'h48; #100;
A = 8'h4C; B = 8'h49; #100;
A = 8'h4C; B = 8'h4A; #100;
A = 8'h4C; B = 8'h4B; #100;
A = 8'h4C; B = 8'h4C; #100;
A = 8'h4C; B = 8'h4D; #100;
A = 8'h4C; B = 8'h4E; #100;
A = 8'h4C; B = 8'h4F; #100;
A = 8'h4C; B = 8'h50; #100;
A = 8'h4C; B = 8'h51; #100;
A = 8'h4C; B = 8'h52; #100;
A = 8'h4C; B = 8'h53; #100;
A = 8'h4C; B = 8'h54; #100;
A = 8'h4C; B = 8'h55; #100;
A = 8'h4C; B = 8'h56; #100;
A = 8'h4C; B = 8'h57; #100;
A = 8'h4C; B = 8'h58; #100;
A = 8'h4C; B = 8'h59; #100;
A = 8'h4C; B = 8'h5A; #100;
A = 8'h4C; B = 8'h5B; #100;
A = 8'h4C; B = 8'h5C; #100;
A = 8'h4C; B = 8'h5D; #100;
A = 8'h4C; B = 8'h5E; #100;
A = 8'h4C; B = 8'h5F; #100;
A = 8'h4C; B = 8'h60; #100;
A = 8'h4C; B = 8'h61; #100;
A = 8'h4C; B = 8'h62; #100;
A = 8'h4C; B = 8'h63; #100;
A = 8'h4C; B = 8'h64; #100;
A = 8'h4C; B = 8'h65; #100;
A = 8'h4C; B = 8'h66; #100;
A = 8'h4C; B = 8'h67; #100;
A = 8'h4C; B = 8'h68; #100;
A = 8'h4C; B = 8'h69; #100;
A = 8'h4C; B = 8'h6A; #100;
A = 8'h4C; B = 8'h6B; #100;
A = 8'h4C; B = 8'h6C; #100;
A = 8'h4C; B = 8'h6D; #100;
A = 8'h4C; B = 8'h6E; #100;
A = 8'h4C; B = 8'h6F; #100;
A = 8'h4C; B = 8'h70; #100;
A = 8'h4C; B = 8'h71; #100;
A = 8'h4C; B = 8'h72; #100;
A = 8'h4C; B = 8'h73; #100;
A = 8'h4C; B = 8'h74; #100;
A = 8'h4C; B = 8'h75; #100;
A = 8'h4C; B = 8'h76; #100;
A = 8'h4C; B = 8'h77; #100;
A = 8'h4C; B = 8'h78; #100;
A = 8'h4C; B = 8'h79; #100;
A = 8'h4C; B = 8'h7A; #100;
A = 8'h4C; B = 8'h7B; #100;
A = 8'h4C; B = 8'h7C; #100;
A = 8'h4C; B = 8'h7D; #100;
A = 8'h4C; B = 8'h7E; #100;
A = 8'h4C; B = 8'h7F; #100;
A = 8'h4C; B = 8'h80; #100;
A = 8'h4C; B = 8'h81; #100;
A = 8'h4C; B = 8'h82; #100;
A = 8'h4C; B = 8'h83; #100;
A = 8'h4C; B = 8'h84; #100;
A = 8'h4C; B = 8'h85; #100;
A = 8'h4C; B = 8'h86; #100;
A = 8'h4C; B = 8'h87; #100;
A = 8'h4C; B = 8'h88; #100;
A = 8'h4C; B = 8'h89; #100;
A = 8'h4C; B = 8'h8A; #100;
A = 8'h4C; B = 8'h8B; #100;
A = 8'h4C; B = 8'h8C; #100;
A = 8'h4C; B = 8'h8D; #100;
A = 8'h4C; B = 8'h8E; #100;
A = 8'h4C; B = 8'h8F; #100;
A = 8'h4C; B = 8'h90; #100;
A = 8'h4C; B = 8'h91; #100;
A = 8'h4C; B = 8'h92; #100;
A = 8'h4C; B = 8'h93; #100;
A = 8'h4C; B = 8'h94; #100;
A = 8'h4C; B = 8'h95; #100;
A = 8'h4C; B = 8'h96; #100;
A = 8'h4C; B = 8'h97; #100;
A = 8'h4C; B = 8'h98; #100;
A = 8'h4C; B = 8'h99; #100;
A = 8'h4C; B = 8'h9A; #100;
A = 8'h4C; B = 8'h9B; #100;
A = 8'h4C; B = 8'h9C; #100;
A = 8'h4C; B = 8'h9D; #100;
A = 8'h4C; B = 8'h9E; #100;
A = 8'h4C; B = 8'h9F; #100;
A = 8'h4C; B = 8'hA0; #100;
A = 8'h4C; B = 8'hA1; #100;
A = 8'h4C; B = 8'hA2; #100;
A = 8'h4C; B = 8'hA3; #100;
A = 8'h4C; B = 8'hA4; #100;
A = 8'h4C; B = 8'hA5; #100;
A = 8'h4C; B = 8'hA6; #100;
A = 8'h4C; B = 8'hA7; #100;
A = 8'h4C; B = 8'hA8; #100;
A = 8'h4C; B = 8'hA9; #100;
A = 8'h4C; B = 8'hAA; #100;
A = 8'h4C; B = 8'hAB; #100;
A = 8'h4C; B = 8'hAC; #100;
A = 8'h4C; B = 8'hAD; #100;
A = 8'h4C; B = 8'hAE; #100;
A = 8'h4C; B = 8'hAF; #100;
A = 8'h4C; B = 8'hB0; #100;
A = 8'h4C; B = 8'hB1; #100;
A = 8'h4C; B = 8'hB2; #100;
A = 8'h4C; B = 8'hB3; #100;
A = 8'h4C; B = 8'hB4; #100;
A = 8'h4C; B = 8'hB5; #100;
A = 8'h4C; B = 8'hB6; #100;
A = 8'h4C; B = 8'hB7; #100;
A = 8'h4C; B = 8'hB8; #100;
A = 8'h4C; B = 8'hB9; #100;
A = 8'h4C; B = 8'hBA; #100;
A = 8'h4C; B = 8'hBB; #100;
A = 8'h4C; B = 8'hBC; #100;
A = 8'h4C; B = 8'hBD; #100;
A = 8'h4C; B = 8'hBE; #100;
A = 8'h4C; B = 8'hBF; #100;
A = 8'h4C; B = 8'hC0; #100;
A = 8'h4C; B = 8'hC1; #100;
A = 8'h4C; B = 8'hC2; #100;
A = 8'h4C; B = 8'hC3; #100;
A = 8'h4C; B = 8'hC4; #100;
A = 8'h4C; B = 8'hC5; #100;
A = 8'h4C; B = 8'hC6; #100;
A = 8'h4C; B = 8'hC7; #100;
A = 8'h4C; B = 8'hC8; #100;
A = 8'h4C; B = 8'hC9; #100;
A = 8'h4C; B = 8'hCA; #100;
A = 8'h4C; B = 8'hCB; #100;
A = 8'h4C; B = 8'hCC; #100;
A = 8'h4C; B = 8'hCD; #100;
A = 8'h4C; B = 8'hCE; #100;
A = 8'h4C; B = 8'hCF; #100;
A = 8'h4C; B = 8'hD0; #100;
A = 8'h4C; B = 8'hD1; #100;
A = 8'h4C; B = 8'hD2; #100;
A = 8'h4C; B = 8'hD3; #100;
A = 8'h4C; B = 8'hD4; #100;
A = 8'h4C; B = 8'hD5; #100;
A = 8'h4C; B = 8'hD6; #100;
A = 8'h4C; B = 8'hD7; #100;
A = 8'h4C; B = 8'hD8; #100;
A = 8'h4C; B = 8'hD9; #100;
A = 8'h4C; B = 8'hDA; #100;
A = 8'h4C; B = 8'hDB; #100;
A = 8'h4C; B = 8'hDC; #100;
A = 8'h4C; B = 8'hDD; #100;
A = 8'h4C; B = 8'hDE; #100;
A = 8'h4C; B = 8'hDF; #100;
A = 8'h4C; B = 8'hE0; #100;
A = 8'h4C; B = 8'hE1; #100;
A = 8'h4C; B = 8'hE2; #100;
A = 8'h4C; B = 8'hE3; #100;
A = 8'h4C; B = 8'hE4; #100;
A = 8'h4C; B = 8'hE5; #100;
A = 8'h4C; B = 8'hE6; #100;
A = 8'h4C; B = 8'hE7; #100;
A = 8'h4C; B = 8'hE8; #100;
A = 8'h4C; B = 8'hE9; #100;
A = 8'h4C; B = 8'hEA; #100;
A = 8'h4C; B = 8'hEB; #100;
A = 8'h4C; B = 8'hEC; #100;
A = 8'h4C; B = 8'hED; #100;
A = 8'h4C; B = 8'hEE; #100;
A = 8'h4C; B = 8'hEF; #100;
A = 8'h4C; B = 8'hF0; #100;
A = 8'h4C; B = 8'hF1; #100;
A = 8'h4C; B = 8'hF2; #100;
A = 8'h4C; B = 8'hF3; #100;
A = 8'h4C; B = 8'hF4; #100;
A = 8'h4C; B = 8'hF5; #100;
A = 8'h4C; B = 8'hF6; #100;
A = 8'h4C; B = 8'hF7; #100;
A = 8'h4C; B = 8'hF8; #100;
A = 8'h4C; B = 8'hF9; #100;
A = 8'h4C; B = 8'hFA; #100;
A = 8'h4C; B = 8'hFB; #100;
A = 8'h4C; B = 8'hFC; #100;
A = 8'h4C; B = 8'hFD; #100;
A = 8'h4C; B = 8'hFE; #100;
A = 8'h4C; B = 8'hFF; #100;
A = 8'h4D; B = 8'h0; #100;
A = 8'h4D; B = 8'h1; #100;
A = 8'h4D; B = 8'h2; #100;
A = 8'h4D; B = 8'h3; #100;
A = 8'h4D; B = 8'h4; #100;
A = 8'h4D; B = 8'h5; #100;
A = 8'h4D; B = 8'h6; #100;
A = 8'h4D; B = 8'h7; #100;
A = 8'h4D; B = 8'h8; #100;
A = 8'h4D; B = 8'h9; #100;
A = 8'h4D; B = 8'hA; #100;
A = 8'h4D; B = 8'hB; #100;
A = 8'h4D; B = 8'hC; #100;
A = 8'h4D; B = 8'hD; #100;
A = 8'h4D; B = 8'hE; #100;
A = 8'h4D; B = 8'hF; #100;
A = 8'h4D; B = 8'h10; #100;
A = 8'h4D; B = 8'h11; #100;
A = 8'h4D; B = 8'h12; #100;
A = 8'h4D; B = 8'h13; #100;
A = 8'h4D; B = 8'h14; #100;
A = 8'h4D; B = 8'h15; #100;
A = 8'h4D; B = 8'h16; #100;
A = 8'h4D; B = 8'h17; #100;
A = 8'h4D; B = 8'h18; #100;
A = 8'h4D; B = 8'h19; #100;
A = 8'h4D; B = 8'h1A; #100;
A = 8'h4D; B = 8'h1B; #100;
A = 8'h4D; B = 8'h1C; #100;
A = 8'h4D; B = 8'h1D; #100;
A = 8'h4D; B = 8'h1E; #100;
A = 8'h4D; B = 8'h1F; #100;
A = 8'h4D; B = 8'h20; #100;
A = 8'h4D; B = 8'h21; #100;
A = 8'h4D; B = 8'h22; #100;
A = 8'h4D; B = 8'h23; #100;
A = 8'h4D; B = 8'h24; #100;
A = 8'h4D; B = 8'h25; #100;
A = 8'h4D; B = 8'h26; #100;
A = 8'h4D; B = 8'h27; #100;
A = 8'h4D; B = 8'h28; #100;
A = 8'h4D; B = 8'h29; #100;
A = 8'h4D; B = 8'h2A; #100;
A = 8'h4D; B = 8'h2B; #100;
A = 8'h4D; B = 8'h2C; #100;
A = 8'h4D; B = 8'h2D; #100;
A = 8'h4D; B = 8'h2E; #100;
A = 8'h4D; B = 8'h2F; #100;
A = 8'h4D; B = 8'h30; #100;
A = 8'h4D; B = 8'h31; #100;
A = 8'h4D; B = 8'h32; #100;
A = 8'h4D; B = 8'h33; #100;
A = 8'h4D; B = 8'h34; #100;
A = 8'h4D; B = 8'h35; #100;
A = 8'h4D; B = 8'h36; #100;
A = 8'h4D; B = 8'h37; #100;
A = 8'h4D; B = 8'h38; #100;
A = 8'h4D; B = 8'h39; #100;
A = 8'h4D; B = 8'h3A; #100;
A = 8'h4D; B = 8'h3B; #100;
A = 8'h4D; B = 8'h3C; #100;
A = 8'h4D; B = 8'h3D; #100;
A = 8'h4D; B = 8'h3E; #100;
A = 8'h4D; B = 8'h3F; #100;
A = 8'h4D; B = 8'h40; #100;
A = 8'h4D; B = 8'h41; #100;
A = 8'h4D; B = 8'h42; #100;
A = 8'h4D; B = 8'h43; #100;
A = 8'h4D; B = 8'h44; #100;
A = 8'h4D; B = 8'h45; #100;
A = 8'h4D; B = 8'h46; #100;
A = 8'h4D; B = 8'h47; #100;
A = 8'h4D; B = 8'h48; #100;
A = 8'h4D; B = 8'h49; #100;
A = 8'h4D; B = 8'h4A; #100;
A = 8'h4D; B = 8'h4B; #100;
A = 8'h4D; B = 8'h4C; #100;
A = 8'h4D; B = 8'h4D; #100;
A = 8'h4D; B = 8'h4E; #100;
A = 8'h4D; B = 8'h4F; #100;
A = 8'h4D; B = 8'h50; #100;
A = 8'h4D; B = 8'h51; #100;
A = 8'h4D; B = 8'h52; #100;
A = 8'h4D; B = 8'h53; #100;
A = 8'h4D; B = 8'h54; #100;
A = 8'h4D; B = 8'h55; #100;
A = 8'h4D; B = 8'h56; #100;
A = 8'h4D; B = 8'h57; #100;
A = 8'h4D; B = 8'h58; #100;
A = 8'h4D; B = 8'h59; #100;
A = 8'h4D; B = 8'h5A; #100;
A = 8'h4D; B = 8'h5B; #100;
A = 8'h4D; B = 8'h5C; #100;
A = 8'h4D; B = 8'h5D; #100;
A = 8'h4D; B = 8'h5E; #100;
A = 8'h4D; B = 8'h5F; #100;
A = 8'h4D; B = 8'h60; #100;
A = 8'h4D; B = 8'h61; #100;
A = 8'h4D; B = 8'h62; #100;
A = 8'h4D; B = 8'h63; #100;
A = 8'h4D; B = 8'h64; #100;
A = 8'h4D; B = 8'h65; #100;
A = 8'h4D; B = 8'h66; #100;
A = 8'h4D; B = 8'h67; #100;
A = 8'h4D; B = 8'h68; #100;
A = 8'h4D; B = 8'h69; #100;
A = 8'h4D; B = 8'h6A; #100;
A = 8'h4D; B = 8'h6B; #100;
A = 8'h4D; B = 8'h6C; #100;
A = 8'h4D; B = 8'h6D; #100;
A = 8'h4D; B = 8'h6E; #100;
A = 8'h4D; B = 8'h6F; #100;
A = 8'h4D; B = 8'h70; #100;
A = 8'h4D; B = 8'h71; #100;
A = 8'h4D; B = 8'h72; #100;
A = 8'h4D; B = 8'h73; #100;
A = 8'h4D; B = 8'h74; #100;
A = 8'h4D; B = 8'h75; #100;
A = 8'h4D; B = 8'h76; #100;
A = 8'h4D; B = 8'h77; #100;
A = 8'h4D; B = 8'h78; #100;
A = 8'h4D; B = 8'h79; #100;
A = 8'h4D; B = 8'h7A; #100;
A = 8'h4D; B = 8'h7B; #100;
A = 8'h4D; B = 8'h7C; #100;
A = 8'h4D; B = 8'h7D; #100;
A = 8'h4D; B = 8'h7E; #100;
A = 8'h4D; B = 8'h7F; #100;
A = 8'h4D; B = 8'h80; #100;
A = 8'h4D; B = 8'h81; #100;
A = 8'h4D; B = 8'h82; #100;
A = 8'h4D; B = 8'h83; #100;
A = 8'h4D; B = 8'h84; #100;
A = 8'h4D; B = 8'h85; #100;
A = 8'h4D; B = 8'h86; #100;
A = 8'h4D; B = 8'h87; #100;
A = 8'h4D; B = 8'h88; #100;
A = 8'h4D; B = 8'h89; #100;
A = 8'h4D; B = 8'h8A; #100;
A = 8'h4D; B = 8'h8B; #100;
A = 8'h4D; B = 8'h8C; #100;
A = 8'h4D; B = 8'h8D; #100;
A = 8'h4D; B = 8'h8E; #100;
A = 8'h4D; B = 8'h8F; #100;
A = 8'h4D; B = 8'h90; #100;
A = 8'h4D; B = 8'h91; #100;
A = 8'h4D; B = 8'h92; #100;
A = 8'h4D; B = 8'h93; #100;
A = 8'h4D; B = 8'h94; #100;
A = 8'h4D; B = 8'h95; #100;
A = 8'h4D; B = 8'h96; #100;
A = 8'h4D; B = 8'h97; #100;
A = 8'h4D; B = 8'h98; #100;
A = 8'h4D; B = 8'h99; #100;
A = 8'h4D; B = 8'h9A; #100;
A = 8'h4D; B = 8'h9B; #100;
A = 8'h4D; B = 8'h9C; #100;
A = 8'h4D; B = 8'h9D; #100;
A = 8'h4D; B = 8'h9E; #100;
A = 8'h4D; B = 8'h9F; #100;
A = 8'h4D; B = 8'hA0; #100;
A = 8'h4D; B = 8'hA1; #100;
A = 8'h4D; B = 8'hA2; #100;
A = 8'h4D; B = 8'hA3; #100;
A = 8'h4D; B = 8'hA4; #100;
A = 8'h4D; B = 8'hA5; #100;
A = 8'h4D; B = 8'hA6; #100;
A = 8'h4D; B = 8'hA7; #100;
A = 8'h4D; B = 8'hA8; #100;
A = 8'h4D; B = 8'hA9; #100;
A = 8'h4D; B = 8'hAA; #100;
A = 8'h4D; B = 8'hAB; #100;
A = 8'h4D; B = 8'hAC; #100;
A = 8'h4D; B = 8'hAD; #100;
A = 8'h4D; B = 8'hAE; #100;
A = 8'h4D; B = 8'hAF; #100;
A = 8'h4D; B = 8'hB0; #100;
A = 8'h4D; B = 8'hB1; #100;
A = 8'h4D; B = 8'hB2; #100;
A = 8'h4D; B = 8'hB3; #100;
A = 8'h4D; B = 8'hB4; #100;
A = 8'h4D; B = 8'hB5; #100;
A = 8'h4D; B = 8'hB6; #100;
A = 8'h4D; B = 8'hB7; #100;
A = 8'h4D; B = 8'hB8; #100;
A = 8'h4D; B = 8'hB9; #100;
A = 8'h4D; B = 8'hBA; #100;
A = 8'h4D; B = 8'hBB; #100;
A = 8'h4D; B = 8'hBC; #100;
A = 8'h4D; B = 8'hBD; #100;
A = 8'h4D; B = 8'hBE; #100;
A = 8'h4D; B = 8'hBF; #100;
A = 8'h4D; B = 8'hC0; #100;
A = 8'h4D; B = 8'hC1; #100;
A = 8'h4D; B = 8'hC2; #100;
A = 8'h4D; B = 8'hC3; #100;
A = 8'h4D; B = 8'hC4; #100;
A = 8'h4D; B = 8'hC5; #100;
A = 8'h4D; B = 8'hC6; #100;
A = 8'h4D; B = 8'hC7; #100;
A = 8'h4D; B = 8'hC8; #100;
A = 8'h4D; B = 8'hC9; #100;
A = 8'h4D; B = 8'hCA; #100;
A = 8'h4D; B = 8'hCB; #100;
A = 8'h4D; B = 8'hCC; #100;
A = 8'h4D; B = 8'hCD; #100;
A = 8'h4D; B = 8'hCE; #100;
A = 8'h4D; B = 8'hCF; #100;
A = 8'h4D; B = 8'hD0; #100;
A = 8'h4D; B = 8'hD1; #100;
A = 8'h4D; B = 8'hD2; #100;
A = 8'h4D; B = 8'hD3; #100;
A = 8'h4D; B = 8'hD4; #100;
A = 8'h4D; B = 8'hD5; #100;
A = 8'h4D; B = 8'hD6; #100;
A = 8'h4D; B = 8'hD7; #100;
A = 8'h4D; B = 8'hD8; #100;
A = 8'h4D; B = 8'hD9; #100;
A = 8'h4D; B = 8'hDA; #100;
A = 8'h4D; B = 8'hDB; #100;
A = 8'h4D; B = 8'hDC; #100;
A = 8'h4D; B = 8'hDD; #100;
A = 8'h4D; B = 8'hDE; #100;
A = 8'h4D; B = 8'hDF; #100;
A = 8'h4D; B = 8'hE0; #100;
A = 8'h4D; B = 8'hE1; #100;
A = 8'h4D; B = 8'hE2; #100;
A = 8'h4D; B = 8'hE3; #100;
A = 8'h4D; B = 8'hE4; #100;
A = 8'h4D; B = 8'hE5; #100;
A = 8'h4D; B = 8'hE6; #100;
A = 8'h4D; B = 8'hE7; #100;
A = 8'h4D; B = 8'hE8; #100;
A = 8'h4D; B = 8'hE9; #100;
A = 8'h4D; B = 8'hEA; #100;
A = 8'h4D; B = 8'hEB; #100;
A = 8'h4D; B = 8'hEC; #100;
A = 8'h4D; B = 8'hED; #100;
A = 8'h4D; B = 8'hEE; #100;
A = 8'h4D; B = 8'hEF; #100;
A = 8'h4D; B = 8'hF0; #100;
A = 8'h4D; B = 8'hF1; #100;
A = 8'h4D; B = 8'hF2; #100;
A = 8'h4D; B = 8'hF3; #100;
A = 8'h4D; B = 8'hF4; #100;
A = 8'h4D; B = 8'hF5; #100;
A = 8'h4D; B = 8'hF6; #100;
A = 8'h4D; B = 8'hF7; #100;
A = 8'h4D; B = 8'hF8; #100;
A = 8'h4D; B = 8'hF9; #100;
A = 8'h4D; B = 8'hFA; #100;
A = 8'h4D; B = 8'hFB; #100;
A = 8'h4D; B = 8'hFC; #100;
A = 8'h4D; B = 8'hFD; #100;
A = 8'h4D; B = 8'hFE; #100;
A = 8'h4D; B = 8'hFF; #100;
A = 8'h4E; B = 8'h0; #100;
A = 8'h4E; B = 8'h1; #100;
A = 8'h4E; B = 8'h2; #100;
A = 8'h4E; B = 8'h3; #100;
A = 8'h4E; B = 8'h4; #100;
A = 8'h4E; B = 8'h5; #100;
A = 8'h4E; B = 8'h6; #100;
A = 8'h4E; B = 8'h7; #100;
A = 8'h4E; B = 8'h8; #100;
A = 8'h4E; B = 8'h9; #100;
A = 8'h4E; B = 8'hA; #100;
A = 8'h4E; B = 8'hB; #100;
A = 8'h4E; B = 8'hC; #100;
A = 8'h4E; B = 8'hD; #100;
A = 8'h4E; B = 8'hE; #100;
A = 8'h4E; B = 8'hF; #100;
A = 8'h4E; B = 8'h10; #100;
A = 8'h4E; B = 8'h11; #100;
A = 8'h4E; B = 8'h12; #100;
A = 8'h4E; B = 8'h13; #100;
A = 8'h4E; B = 8'h14; #100;
A = 8'h4E; B = 8'h15; #100;
A = 8'h4E; B = 8'h16; #100;
A = 8'h4E; B = 8'h17; #100;
A = 8'h4E; B = 8'h18; #100;
A = 8'h4E; B = 8'h19; #100;
A = 8'h4E; B = 8'h1A; #100;
A = 8'h4E; B = 8'h1B; #100;
A = 8'h4E; B = 8'h1C; #100;
A = 8'h4E; B = 8'h1D; #100;
A = 8'h4E; B = 8'h1E; #100;
A = 8'h4E; B = 8'h1F; #100;
A = 8'h4E; B = 8'h20; #100;
A = 8'h4E; B = 8'h21; #100;
A = 8'h4E; B = 8'h22; #100;
A = 8'h4E; B = 8'h23; #100;
A = 8'h4E; B = 8'h24; #100;
A = 8'h4E; B = 8'h25; #100;
A = 8'h4E; B = 8'h26; #100;
A = 8'h4E; B = 8'h27; #100;
A = 8'h4E; B = 8'h28; #100;
A = 8'h4E; B = 8'h29; #100;
A = 8'h4E; B = 8'h2A; #100;
A = 8'h4E; B = 8'h2B; #100;
A = 8'h4E; B = 8'h2C; #100;
A = 8'h4E; B = 8'h2D; #100;
A = 8'h4E; B = 8'h2E; #100;
A = 8'h4E; B = 8'h2F; #100;
A = 8'h4E; B = 8'h30; #100;
A = 8'h4E; B = 8'h31; #100;
A = 8'h4E; B = 8'h32; #100;
A = 8'h4E; B = 8'h33; #100;
A = 8'h4E; B = 8'h34; #100;
A = 8'h4E; B = 8'h35; #100;
A = 8'h4E; B = 8'h36; #100;
A = 8'h4E; B = 8'h37; #100;
A = 8'h4E; B = 8'h38; #100;
A = 8'h4E; B = 8'h39; #100;
A = 8'h4E; B = 8'h3A; #100;
A = 8'h4E; B = 8'h3B; #100;
A = 8'h4E; B = 8'h3C; #100;
A = 8'h4E; B = 8'h3D; #100;
A = 8'h4E; B = 8'h3E; #100;
A = 8'h4E; B = 8'h3F; #100;
A = 8'h4E; B = 8'h40; #100;
A = 8'h4E; B = 8'h41; #100;
A = 8'h4E; B = 8'h42; #100;
A = 8'h4E; B = 8'h43; #100;
A = 8'h4E; B = 8'h44; #100;
A = 8'h4E; B = 8'h45; #100;
A = 8'h4E; B = 8'h46; #100;
A = 8'h4E; B = 8'h47; #100;
A = 8'h4E; B = 8'h48; #100;
A = 8'h4E; B = 8'h49; #100;
A = 8'h4E; B = 8'h4A; #100;
A = 8'h4E; B = 8'h4B; #100;
A = 8'h4E; B = 8'h4C; #100;
A = 8'h4E; B = 8'h4D; #100;
A = 8'h4E; B = 8'h4E; #100;
A = 8'h4E; B = 8'h4F; #100;
A = 8'h4E; B = 8'h50; #100;
A = 8'h4E; B = 8'h51; #100;
A = 8'h4E; B = 8'h52; #100;
A = 8'h4E; B = 8'h53; #100;
A = 8'h4E; B = 8'h54; #100;
A = 8'h4E; B = 8'h55; #100;
A = 8'h4E; B = 8'h56; #100;
A = 8'h4E; B = 8'h57; #100;
A = 8'h4E; B = 8'h58; #100;
A = 8'h4E; B = 8'h59; #100;
A = 8'h4E; B = 8'h5A; #100;
A = 8'h4E; B = 8'h5B; #100;
A = 8'h4E; B = 8'h5C; #100;
A = 8'h4E; B = 8'h5D; #100;
A = 8'h4E; B = 8'h5E; #100;
A = 8'h4E; B = 8'h5F; #100;
A = 8'h4E; B = 8'h60; #100;
A = 8'h4E; B = 8'h61; #100;
A = 8'h4E; B = 8'h62; #100;
A = 8'h4E; B = 8'h63; #100;
A = 8'h4E; B = 8'h64; #100;
A = 8'h4E; B = 8'h65; #100;
A = 8'h4E; B = 8'h66; #100;
A = 8'h4E; B = 8'h67; #100;
A = 8'h4E; B = 8'h68; #100;
A = 8'h4E; B = 8'h69; #100;
A = 8'h4E; B = 8'h6A; #100;
A = 8'h4E; B = 8'h6B; #100;
A = 8'h4E; B = 8'h6C; #100;
A = 8'h4E; B = 8'h6D; #100;
A = 8'h4E; B = 8'h6E; #100;
A = 8'h4E; B = 8'h6F; #100;
A = 8'h4E; B = 8'h70; #100;
A = 8'h4E; B = 8'h71; #100;
A = 8'h4E; B = 8'h72; #100;
A = 8'h4E; B = 8'h73; #100;
A = 8'h4E; B = 8'h74; #100;
A = 8'h4E; B = 8'h75; #100;
A = 8'h4E; B = 8'h76; #100;
A = 8'h4E; B = 8'h77; #100;
A = 8'h4E; B = 8'h78; #100;
A = 8'h4E; B = 8'h79; #100;
A = 8'h4E; B = 8'h7A; #100;
A = 8'h4E; B = 8'h7B; #100;
A = 8'h4E; B = 8'h7C; #100;
A = 8'h4E; B = 8'h7D; #100;
A = 8'h4E; B = 8'h7E; #100;
A = 8'h4E; B = 8'h7F; #100;
A = 8'h4E; B = 8'h80; #100;
A = 8'h4E; B = 8'h81; #100;
A = 8'h4E; B = 8'h82; #100;
A = 8'h4E; B = 8'h83; #100;
A = 8'h4E; B = 8'h84; #100;
A = 8'h4E; B = 8'h85; #100;
A = 8'h4E; B = 8'h86; #100;
A = 8'h4E; B = 8'h87; #100;
A = 8'h4E; B = 8'h88; #100;
A = 8'h4E; B = 8'h89; #100;
A = 8'h4E; B = 8'h8A; #100;
A = 8'h4E; B = 8'h8B; #100;
A = 8'h4E; B = 8'h8C; #100;
A = 8'h4E; B = 8'h8D; #100;
A = 8'h4E; B = 8'h8E; #100;
A = 8'h4E; B = 8'h8F; #100;
A = 8'h4E; B = 8'h90; #100;
A = 8'h4E; B = 8'h91; #100;
A = 8'h4E; B = 8'h92; #100;
A = 8'h4E; B = 8'h93; #100;
A = 8'h4E; B = 8'h94; #100;
A = 8'h4E; B = 8'h95; #100;
A = 8'h4E; B = 8'h96; #100;
A = 8'h4E; B = 8'h97; #100;
A = 8'h4E; B = 8'h98; #100;
A = 8'h4E; B = 8'h99; #100;
A = 8'h4E; B = 8'h9A; #100;
A = 8'h4E; B = 8'h9B; #100;
A = 8'h4E; B = 8'h9C; #100;
A = 8'h4E; B = 8'h9D; #100;
A = 8'h4E; B = 8'h9E; #100;
A = 8'h4E; B = 8'h9F; #100;
A = 8'h4E; B = 8'hA0; #100;
A = 8'h4E; B = 8'hA1; #100;
A = 8'h4E; B = 8'hA2; #100;
A = 8'h4E; B = 8'hA3; #100;
A = 8'h4E; B = 8'hA4; #100;
A = 8'h4E; B = 8'hA5; #100;
A = 8'h4E; B = 8'hA6; #100;
A = 8'h4E; B = 8'hA7; #100;
A = 8'h4E; B = 8'hA8; #100;
A = 8'h4E; B = 8'hA9; #100;
A = 8'h4E; B = 8'hAA; #100;
A = 8'h4E; B = 8'hAB; #100;
A = 8'h4E; B = 8'hAC; #100;
A = 8'h4E; B = 8'hAD; #100;
A = 8'h4E; B = 8'hAE; #100;
A = 8'h4E; B = 8'hAF; #100;
A = 8'h4E; B = 8'hB0; #100;
A = 8'h4E; B = 8'hB1; #100;
A = 8'h4E; B = 8'hB2; #100;
A = 8'h4E; B = 8'hB3; #100;
A = 8'h4E; B = 8'hB4; #100;
A = 8'h4E; B = 8'hB5; #100;
A = 8'h4E; B = 8'hB6; #100;
A = 8'h4E; B = 8'hB7; #100;
A = 8'h4E; B = 8'hB8; #100;
A = 8'h4E; B = 8'hB9; #100;
A = 8'h4E; B = 8'hBA; #100;
A = 8'h4E; B = 8'hBB; #100;
A = 8'h4E; B = 8'hBC; #100;
A = 8'h4E; B = 8'hBD; #100;
A = 8'h4E; B = 8'hBE; #100;
A = 8'h4E; B = 8'hBF; #100;
A = 8'h4E; B = 8'hC0; #100;
A = 8'h4E; B = 8'hC1; #100;
A = 8'h4E; B = 8'hC2; #100;
A = 8'h4E; B = 8'hC3; #100;
A = 8'h4E; B = 8'hC4; #100;
A = 8'h4E; B = 8'hC5; #100;
A = 8'h4E; B = 8'hC6; #100;
A = 8'h4E; B = 8'hC7; #100;
A = 8'h4E; B = 8'hC8; #100;
A = 8'h4E; B = 8'hC9; #100;
A = 8'h4E; B = 8'hCA; #100;
A = 8'h4E; B = 8'hCB; #100;
A = 8'h4E; B = 8'hCC; #100;
A = 8'h4E; B = 8'hCD; #100;
A = 8'h4E; B = 8'hCE; #100;
A = 8'h4E; B = 8'hCF; #100;
A = 8'h4E; B = 8'hD0; #100;
A = 8'h4E; B = 8'hD1; #100;
A = 8'h4E; B = 8'hD2; #100;
A = 8'h4E; B = 8'hD3; #100;
A = 8'h4E; B = 8'hD4; #100;
A = 8'h4E; B = 8'hD5; #100;
A = 8'h4E; B = 8'hD6; #100;
A = 8'h4E; B = 8'hD7; #100;
A = 8'h4E; B = 8'hD8; #100;
A = 8'h4E; B = 8'hD9; #100;
A = 8'h4E; B = 8'hDA; #100;
A = 8'h4E; B = 8'hDB; #100;
A = 8'h4E; B = 8'hDC; #100;
A = 8'h4E; B = 8'hDD; #100;
A = 8'h4E; B = 8'hDE; #100;
A = 8'h4E; B = 8'hDF; #100;
A = 8'h4E; B = 8'hE0; #100;
A = 8'h4E; B = 8'hE1; #100;
A = 8'h4E; B = 8'hE2; #100;
A = 8'h4E; B = 8'hE3; #100;
A = 8'h4E; B = 8'hE4; #100;
A = 8'h4E; B = 8'hE5; #100;
A = 8'h4E; B = 8'hE6; #100;
A = 8'h4E; B = 8'hE7; #100;
A = 8'h4E; B = 8'hE8; #100;
A = 8'h4E; B = 8'hE9; #100;
A = 8'h4E; B = 8'hEA; #100;
A = 8'h4E; B = 8'hEB; #100;
A = 8'h4E; B = 8'hEC; #100;
A = 8'h4E; B = 8'hED; #100;
A = 8'h4E; B = 8'hEE; #100;
A = 8'h4E; B = 8'hEF; #100;
A = 8'h4E; B = 8'hF0; #100;
A = 8'h4E; B = 8'hF1; #100;
A = 8'h4E; B = 8'hF2; #100;
A = 8'h4E; B = 8'hF3; #100;
A = 8'h4E; B = 8'hF4; #100;
A = 8'h4E; B = 8'hF5; #100;
A = 8'h4E; B = 8'hF6; #100;
A = 8'h4E; B = 8'hF7; #100;
A = 8'h4E; B = 8'hF8; #100;
A = 8'h4E; B = 8'hF9; #100;
A = 8'h4E; B = 8'hFA; #100;
A = 8'h4E; B = 8'hFB; #100;
A = 8'h4E; B = 8'hFC; #100;
A = 8'h4E; B = 8'hFD; #100;
A = 8'h4E; B = 8'hFE; #100;
A = 8'h4E; B = 8'hFF; #100;
A = 8'h4F; B = 8'h0; #100;
A = 8'h4F; B = 8'h1; #100;
A = 8'h4F; B = 8'h2; #100;
A = 8'h4F; B = 8'h3; #100;
A = 8'h4F; B = 8'h4; #100;
A = 8'h4F; B = 8'h5; #100;
A = 8'h4F; B = 8'h6; #100;
A = 8'h4F; B = 8'h7; #100;
A = 8'h4F; B = 8'h8; #100;
A = 8'h4F; B = 8'h9; #100;
A = 8'h4F; B = 8'hA; #100;
A = 8'h4F; B = 8'hB; #100;
A = 8'h4F; B = 8'hC; #100;
A = 8'h4F; B = 8'hD; #100;
A = 8'h4F; B = 8'hE; #100;
A = 8'h4F; B = 8'hF; #100;
A = 8'h4F; B = 8'h10; #100;
A = 8'h4F; B = 8'h11; #100;
A = 8'h4F; B = 8'h12; #100;
A = 8'h4F; B = 8'h13; #100;
A = 8'h4F; B = 8'h14; #100;
A = 8'h4F; B = 8'h15; #100;
A = 8'h4F; B = 8'h16; #100;
A = 8'h4F; B = 8'h17; #100;
A = 8'h4F; B = 8'h18; #100;
A = 8'h4F; B = 8'h19; #100;
A = 8'h4F; B = 8'h1A; #100;
A = 8'h4F; B = 8'h1B; #100;
A = 8'h4F; B = 8'h1C; #100;
A = 8'h4F; B = 8'h1D; #100;
A = 8'h4F; B = 8'h1E; #100;
A = 8'h4F; B = 8'h1F; #100;
A = 8'h4F; B = 8'h20; #100;
A = 8'h4F; B = 8'h21; #100;
A = 8'h4F; B = 8'h22; #100;
A = 8'h4F; B = 8'h23; #100;
A = 8'h4F; B = 8'h24; #100;
A = 8'h4F; B = 8'h25; #100;
A = 8'h4F; B = 8'h26; #100;
A = 8'h4F; B = 8'h27; #100;
A = 8'h4F; B = 8'h28; #100;
A = 8'h4F; B = 8'h29; #100;
A = 8'h4F; B = 8'h2A; #100;
A = 8'h4F; B = 8'h2B; #100;
A = 8'h4F; B = 8'h2C; #100;
A = 8'h4F; B = 8'h2D; #100;
A = 8'h4F; B = 8'h2E; #100;
A = 8'h4F; B = 8'h2F; #100;
A = 8'h4F; B = 8'h30; #100;
A = 8'h4F; B = 8'h31; #100;
A = 8'h4F; B = 8'h32; #100;
A = 8'h4F; B = 8'h33; #100;
A = 8'h4F; B = 8'h34; #100;
A = 8'h4F; B = 8'h35; #100;
A = 8'h4F; B = 8'h36; #100;
A = 8'h4F; B = 8'h37; #100;
A = 8'h4F; B = 8'h38; #100;
A = 8'h4F; B = 8'h39; #100;
A = 8'h4F; B = 8'h3A; #100;
A = 8'h4F; B = 8'h3B; #100;
A = 8'h4F; B = 8'h3C; #100;
A = 8'h4F; B = 8'h3D; #100;
A = 8'h4F; B = 8'h3E; #100;
A = 8'h4F; B = 8'h3F; #100;
A = 8'h4F; B = 8'h40; #100;
A = 8'h4F; B = 8'h41; #100;
A = 8'h4F; B = 8'h42; #100;
A = 8'h4F; B = 8'h43; #100;
A = 8'h4F; B = 8'h44; #100;
A = 8'h4F; B = 8'h45; #100;
A = 8'h4F; B = 8'h46; #100;
A = 8'h4F; B = 8'h47; #100;
A = 8'h4F; B = 8'h48; #100;
A = 8'h4F; B = 8'h49; #100;
A = 8'h4F; B = 8'h4A; #100;
A = 8'h4F; B = 8'h4B; #100;
A = 8'h4F; B = 8'h4C; #100;
A = 8'h4F; B = 8'h4D; #100;
A = 8'h4F; B = 8'h4E; #100;
A = 8'h4F; B = 8'h4F; #100;
A = 8'h4F; B = 8'h50; #100;
A = 8'h4F; B = 8'h51; #100;
A = 8'h4F; B = 8'h52; #100;
A = 8'h4F; B = 8'h53; #100;
A = 8'h4F; B = 8'h54; #100;
A = 8'h4F; B = 8'h55; #100;
A = 8'h4F; B = 8'h56; #100;
A = 8'h4F; B = 8'h57; #100;
A = 8'h4F; B = 8'h58; #100;
A = 8'h4F; B = 8'h59; #100;
A = 8'h4F; B = 8'h5A; #100;
A = 8'h4F; B = 8'h5B; #100;
A = 8'h4F; B = 8'h5C; #100;
A = 8'h4F; B = 8'h5D; #100;
A = 8'h4F; B = 8'h5E; #100;
A = 8'h4F; B = 8'h5F; #100;
A = 8'h4F; B = 8'h60; #100;
A = 8'h4F; B = 8'h61; #100;
A = 8'h4F; B = 8'h62; #100;
A = 8'h4F; B = 8'h63; #100;
A = 8'h4F; B = 8'h64; #100;
A = 8'h4F; B = 8'h65; #100;
A = 8'h4F; B = 8'h66; #100;
A = 8'h4F; B = 8'h67; #100;
A = 8'h4F; B = 8'h68; #100;
A = 8'h4F; B = 8'h69; #100;
A = 8'h4F; B = 8'h6A; #100;
A = 8'h4F; B = 8'h6B; #100;
A = 8'h4F; B = 8'h6C; #100;
A = 8'h4F; B = 8'h6D; #100;
A = 8'h4F; B = 8'h6E; #100;
A = 8'h4F; B = 8'h6F; #100;
A = 8'h4F; B = 8'h70; #100;
A = 8'h4F; B = 8'h71; #100;
A = 8'h4F; B = 8'h72; #100;
A = 8'h4F; B = 8'h73; #100;
A = 8'h4F; B = 8'h74; #100;
A = 8'h4F; B = 8'h75; #100;
A = 8'h4F; B = 8'h76; #100;
A = 8'h4F; B = 8'h77; #100;
A = 8'h4F; B = 8'h78; #100;
A = 8'h4F; B = 8'h79; #100;
A = 8'h4F; B = 8'h7A; #100;
A = 8'h4F; B = 8'h7B; #100;
A = 8'h4F; B = 8'h7C; #100;
A = 8'h4F; B = 8'h7D; #100;
A = 8'h4F; B = 8'h7E; #100;
A = 8'h4F; B = 8'h7F; #100;
A = 8'h4F; B = 8'h80; #100;
A = 8'h4F; B = 8'h81; #100;
A = 8'h4F; B = 8'h82; #100;
A = 8'h4F; B = 8'h83; #100;
A = 8'h4F; B = 8'h84; #100;
A = 8'h4F; B = 8'h85; #100;
A = 8'h4F; B = 8'h86; #100;
A = 8'h4F; B = 8'h87; #100;
A = 8'h4F; B = 8'h88; #100;
A = 8'h4F; B = 8'h89; #100;
A = 8'h4F; B = 8'h8A; #100;
A = 8'h4F; B = 8'h8B; #100;
A = 8'h4F; B = 8'h8C; #100;
A = 8'h4F; B = 8'h8D; #100;
A = 8'h4F; B = 8'h8E; #100;
A = 8'h4F; B = 8'h8F; #100;
A = 8'h4F; B = 8'h90; #100;
A = 8'h4F; B = 8'h91; #100;
A = 8'h4F; B = 8'h92; #100;
A = 8'h4F; B = 8'h93; #100;
A = 8'h4F; B = 8'h94; #100;
A = 8'h4F; B = 8'h95; #100;
A = 8'h4F; B = 8'h96; #100;
A = 8'h4F; B = 8'h97; #100;
A = 8'h4F; B = 8'h98; #100;
A = 8'h4F; B = 8'h99; #100;
A = 8'h4F; B = 8'h9A; #100;
A = 8'h4F; B = 8'h9B; #100;
A = 8'h4F; B = 8'h9C; #100;
A = 8'h4F; B = 8'h9D; #100;
A = 8'h4F; B = 8'h9E; #100;
A = 8'h4F; B = 8'h9F; #100;
A = 8'h4F; B = 8'hA0; #100;
A = 8'h4F; B = 8'hA1; #100;
A = 8'h4F; B = 8'hA2; #100;
A = 8'h4F; B = 8'hA3; #100;
A = 8'h4F; B = 8'hA4; #100;
A = 8'h4F; B = 8'hA5; #100;
A = 8'h4F; B = 8'hA6; #100;
A = 8'h4F; B = 8'hA7; #100;
A = 8'h4F; B = 8'hA8; #100;
A = 8'h4F; B = 8'hA9; #100;
A = 8'h4F; B = 8'hAA; #100;
A = 8'h4F; B = 8'hAB; #100;
A = 8'h4F; B = 8'hAC; #100;
A = 8'h4F; B = 8'hAD; #100;
A = 8'h4F; B = 8'hAE; #100;
A = 8'h4F; B = 8'hAF; #100;
A = 8'h4F; B = 8'hB0; #100;
A = 8'h4F; B = 8'hB1; #100;
A = 8'h4F; B = 8'hB2; #100;
A = 8'h4F; B = 8'hB3; #100;
A = 8'h4F; B = 8'hB4; #100;
A = 8'h4F; B = 8'hB5; #100;
A = 8'h4F; B = 8'hB6; #100;
A = 8'h4F; B = 8'hB7; #100;
A = 8'h4F; B = 8'hB8; #100;
A = 8'h4F; B = 8'hB9; #100;
A = 8'h4F; B = 8'hBA; #100;
A = 8'h4F; B = 8'hBB; #100;
A = 8'h4F; B = 8'hBC; #100;
A = 8'h4F; B = 8'hBD; #100;
A = 8'h4F; B = 8'hBE; #100;
A = 8'h4F; B = 8'hBF; #100;
A = 8'h4F; B = 8'hC0; #100;
A = 8'h4F; B = 8'hC1; #100;
A = 8'h4F; B = 8'hC2; #100;
A = 8'h4F; B = 8'hC3; #100;
A = 8'h4F; B = 8'hC4; #100;
A = 8'h4F; B = 8'hC5; #100;
A = 8'h4F; B = 8'hC6; #100;
A = 8'h4F; B = 8'hC7; #100;
A = 8'h4F; B = 8'hC8; #100;
A = 8'h4F; B = 8'hC9; #100;
A = 8'h4F; B = 8'hCA; #100;
A = 8'h4F; B = 8'hCB; #100;
A = 8'h4F; B = 8'hCC; #100;
A = 8'h4F; B = 8'hCD; #100;
A = 8'h4F; B = 8'hCE; #100;
A = 8'h4F; B = 8'hCF; #100;
A = 8'h4F; B = 8'hD0; #100;
A = 8'h4F; B = 8'hD1; #100;
A = 8'h4F; B = 8'hD2; #100;
A = 8'h4F; B = 8'hD3; #100;
A = 8'h4F; B = 8'hD4; #100;
A = 8'h4F; B = 8'hD5; #100;
A = 8'h4F; B = 8'hD6; #100;
A = 8'h4F; B = 8'hD7; #100;
A = 8'h4F; B = 8'hD8; #100;
A = 8'h4F; B = 8'hD9; #100;
A = 8'h4F; B = 8'hDA; #100;
A = 8'h4F; B = 8'hDB; #100;
A = 8'h4F; B = 8'hDC; #100;
A = 8'h4F; B = 8'hDD; #100;
A = 8'h4F; B = 8'hDE; #100;
A = 8'h4F; B = 8'hDF; #100;
A = 8'h4F; B = 8'hE0; #100;
A = 8'h4F; B = 8'hE1; #100;
A = 8'h4F; B = 8'hE2; #100;
A = 8'h4F; B = 8'hE3; #100;
A = 8'h4F; B = 8'hE4; #100;
A = 8'h4F; B = 8'hE5; #100;
A = 8'h4F; B = 8'hE6; #100;
A = 8'h4F; B = 8'hE7; #100;
A = 8'h4F; B = 8'hE8; #100;
A = 8'h4F; B = 8'hE9; #100;
A = 8'h4F; B = 8'hEA; #100;
A = 8'h4F; B = 8'hEB; #100;
A = 8'h4F; B = 8'hEC; #100;
A = 8'h4F; B = 8'hED; #100;
A = 8'h4F; B = 8'hEE; #100;
A = 8'h4F; B = 8'hEF; #100;
A = 8'h4F; B = 8'hF0; #100;
A = 8'h4F; B = 8'hF1; #100;
A = 8'h4F; B = 8'hF2; #100;
A = 8'h4F; B = 8'hF3; #100;
A = 8'h4F; B = 8'hF4; #100;
A = 8'h4F; B = 8'hF5; #100;
A = 8'h4F; B = 8'hF6; #100;
A = 8'h4F; B = 8'hF7; #100;
A = 8'h4F; B = 8'hF8; #100;
A = 8'h4F; B = 8'hF9; #100;
A = 8'h4F; B = 8'hFA; #100;
A = 8'h4F; B = 8'hFB; #100;
A = 8'h4F; B = 8'hFC; #100;
A = 8'h4F; B = 8'hFD; #100;
A = 8'h4F; B = 8'hFE; #100;
A = 8'h4F; B = 8'hFF; #100;
A = 8'h50; B = 8'h0; #100;
A = 8'h50; B = 8'h1; #100;
A = 8'h50; B = 8'h2; #100;
A = 8'h50; B = 8'h3; #100;
A = 8'h50; B = 8'h4; #100;
A = 8'h50; B = 8'h5; #100;
A = 8'h50; B = 8'h6; #100;
A = 8'h50; B = 8'h7; #100;
A = 8'h50; B = 8'h8; #100;
A = 8'h50; B = 8'h9; #100;
A = 8'h50; B = 8'hA; #100;
A = 8'h50; B = 8'hB; #100;
A = 8'h50; B = 8'hC; #100;
A = 8'h50; B = 8'hD; #100;
A = 8'h50; B = 8'hE; #100;
A = 8'h50; B = 8'hF; #100;
A = 8'h50; B = 8'h10; #100;
A = 8'h50; B = 8'h11; #100;
A = 8'h50; B = 8'h12; #100;
A = 8'h50; B = 8'h13; #100;
A = 8'h50; B = 8'h14; #100;
A = 8'h50; B = 8'h15; #100;
A = 8'h50; B = 8'h16; #100;
A = 8'h50; B = 8'h17; #100;
A = 8'h50; B = 8'h18; #100;
A = 8'h50; B = 8'h19; #100;
A = 8'h50; B = 8'h1A; #100;
A = 8'h50; B = 8'h1B; #100;
A = 8'h50; B = 8'h1C; #100;
A = 8'h50; B = 8'h1D; #100;
A = 8'h50; B = 8'h1E; #100;
A = 8'h50; B = 8'h1F; #100;
A = 8'h50; B = 8'h20; #100;
A = 8'h50; B = 8'h21; #100;
A = 8'h50; B = 8'h22; #100;
A = 8'h50; B = 8'h23; #100;
A = 8'h50; B = 8'h24; #100;
A = 8'h50; B = 8'h25; #100;
A = 8'h50; B = 8'h26; #100;
A = 8'h50; B = 8'h27; #100;
A = 8'h50; B = 8'h28; #100;
A = 8'h50; B = 8'h29; #100;
A = 8'h50; B = 8'h2A; #100;
A = 8'h50; B = 8'h2B; #100;
A = 8'h50; B = 8'h2C; #100;
A = 8'h50; B = 8'h2D; #100;
A = 8'h50; B = 8'h2E; #100;
A = 8'h50; B = 8'h2F; #100;
A = 8'h50; B = 8'h30; #100;
A = 8'h50; B = 8'h31; #100;
A = 8'h50; B = 8'h32; #100;
A = 8'h50; B = 8'h33; #100;
A = 8'h50; B = 8'h34; #100;
A = 8'h50; B = 8'h35; #100;
A = 8'h50; B = 8'h36; #100;
A = 8'h50; B = 8'h37; #100;
A = 8'h50; B = 8'h38; #100;
A = 8'h50; B = 8'h39; #100;
A = 8'h50; B = 8'h3A; #100;
A = 8'h50; B = 8'h3B; #100;
A = 8'h50; B = 8'h3C; #100;
A = 8'h50; B = 8'h3D; #100;
A = 8'h50; B = 8'h3E; #100;
A = 8'h50; B = 8'h3F; #100;
A = 8'h50; B = 8'h40; #100;
A = 8'h50; B = 8'h41; #100;
A = 8'h50; B = 8'h42; #100;
A = 8'h50; B = 8'h43; #100;
A = 8'h50; B = 8'h44; #100;
A = 8'h50; B = 8'h45; #100;
A = 8'h50; B = 8'h46; #100;
A = 8'h50; B = 8'h47; #100;
A = 8'h50; B = 8'h48; #100;
A = 8'h50; B = 8'h49; #100;
A = 8'h50; B = 8'h4A; #100;
A = 8'h50; B = 8'h4B; #100;
A = 8'h50; B = 8'h4C; #100;
A = 8'h50; B = 8'h4D; #100;
A = 8'h50; B = 8'h4E; #100;
A = 8'h50; B = 8'h4F; #100;
A = 8'h50; B = 8'h50; #100;
A = 8'h50; B = 8'h51; #100;
A = 8'h50; B = 8'h52; #100;
A = 8'h50; B = 8'h53; #100;
A = 8'h50; B = 8'h54; #100;
A = 8'h50; B = 8'h55; #100;
A = 8'h50; B = 8'h56; #100;
A = 8'h50; B = 8'h57; #100;
A = 8'h50; B = 8'h58; #100;
A = 8'h50; B = 8'h59; #100;
A = 8'h50; B = 8'h5A; #100;
A = 8'h50; B = 8'h5B; #100;
A = 8'h50; B = 8'h5C; #100;
A = 8'h50; B = 8'h5D; #100;
A = 8'h50; B = 8'h5E; #100;
A = 8'h50; B = 8'h5F; #100;
A = 8'h50; B = 8'h60; #100;
A = 8'h50; B = 8'h61; #100;
A = 8'h50; B = 8'h62; #100;
A = 8'h50; B = 8'h63; #100;
A = 8'h50; B = 8'h64; #100;
A = 8'h50; B = 8'h65; #100;
A = 8'h50; B = 8'h66; #100;
A = 8'h50; B = 8'h67; #100;
A = 8'h50; B = 8'h68; #100;
A = 8'h50; B = 8'h69; #100;
A = 8'h50; B = 8'h6A; #100;
A = 8'h50; B = 8'h6B; #100;
A = 8'h50; B = 8'h6C; #100;
A = 8'h50; B = 8'h6D; #100;
A = 8'h50; B = 8'h6E; #100;
A = 8'h50; B = 8'h6F; #100;
A = 8'h50; B = 8'h70; #100;
A = 8'h50; B = 8'h71; #100;
A = 8'h50; B = 8'h72; #100;
A = 8'h50; B = 8'h73; #100;
A = 8'h50; B = 8'h74; #100;
A = 8'h50; B = 8'h75; #100;
A = 8'h50; B = 8'h76; #100;
A = 8'h50; B = 8'h77; #100;
A = 8'h50; B = 8'h78; #100;
A = 8'h50; B = 8'h79; #100;
A = 8'h50; B = 8'h7A; #100;
A = 8'h50; B = 8'h7B; #100;
A = 8'h50; B = 8'h7C; #100;
A = 8'h50; B = 8'h7D; #100;
A = 8'h50; B = 8'h7E; #100;
A = 8'h50; B = 8'h7F; #100;
A = 8'h50; B = 8'h80; #100;
A = 8'h50; B = 8'h81; #100;
A = 8'h50; B = 8'h82; #100;
A = 8'h50; B = 8'h83; #100;
A = 8'h50; B = 8'h84; #100;
A = 8'h50; B = 8'h85; #100;
A = 8'h50; B = 8'h86; #100;
A = 8'h50; B = 8'h87; #100;
A = 8'h50; B = 8'h88; #100;
A = 8'h50; B = 8'h89; #100;
A = 8'h50; B = 8'h8A; #100;
A = 8'h50; B = 8'h8B; #100;
A = 8'h50; B = 8'h8C; #100;
A = 8'h50; B = 8'h8D; #100;
A = 8'h50; B = 8'h8E; #100;
A = 8'h50; B = 8'h8F; #100;
A = 8'h50; B = 8'h90; #100;
A = 8'h50; B = 8'h91; #100;
A = 8'h50; B = 8'h92; #100;
A = 8'h50; B = 8'h93; #100;
A = 8'h50; B = 8'h94; #100;
A = 8'h50; B = 8'h95; #100;
A = 8'h50; B = 8'h96; #100;
A = 8'h50; B = 8'h97; #100;
A = 8'h50; B = 8'h98; #100;
A = 8'h50; B = 8'h99; #100;
A = 8'h50; B = 8'h9A; #100;
A = 8'h50; B = 8'h9B; #100;
A = 8'h50; B = 8'h9C; #100;
A = 8'h50; B = 8'h9D; #100;
A = 8'h50; B = 8'h9E; #100;
A = 8'h50; B = 8'h9F; #100;
A = 8'h50; B = 8'hA0; #100;
A = 8'h50; B = 8'hA1; #100;
A = 8'h50; B = 8'hA2; #100;
A = 8'h50; B = 8'hA3; #100;
A = 8'h50; B = 8'hA4; #100;
A = 8'h50; B = 8'hA5; #100;
A = 8'h50; B = 8'hA6; #100;
A = 8'h50; B = 8'hA7; #100;
A = 8'h50; B = 8'hA8; #100;
A = 8'h50; B = 8'hA9; #100;
A = 8'h50; B = 8'hAA; #100;
A = 8'h50; B = 8'hAB; #100;
A = 8'h50; B = 8'hAC; #100;
A = 8'h50; B = 8'hAD; #100;
A = 8'h50; B = 8'hAE; #100;
A = 8'h50; B = 8'hAF; #100;
A = 8'h50; B = 8'hB0; #100;
A = 8'h50; B = 8'hB1; #100;
A = 8'h50; B = 8'hB2; #100;
A = 8'h50; B = 8'hB3; #100;
A = 8'h50; B = 8'hB4; #100;
A = 8'h50; B = 8'hB5; #100;
A = 8'h50; B = 8'hB6; #100;
A = 8'h50; B = 8'hB7; #100;
A = 8'h50; B = 8'hB8; #100;
A = 8'h50; B = 8'hB9; #100;
A = 8'h50; B = 8'hBA; #100;
A = 8'h50; B = 8'hBB; #100;
A = 8'h50; B = 8'hBC; #100;
A = 8'h50; B = 8'hBD; #100;
A = 8'h50; B = 8'hBE; #100;
A = 8'h50; B = 8'hBF; #100;
A = 8'h50; B = 8'hC0; #100;
A = 8'h50; B = 8'hC1; #100;
A = 8'h50; B = 8'hC2; #100;
A = 8'h50; B = 8'hC3; #100;
A = 8'h50; B = 8'hC4; #100;
A = 8'h50; B = 8'hC5; #100;
A = 8'h50; B = 8'hC6; #100;
A = 8'h50; B = 8'hC7; #100;
A = 8'h50; B = 8'hC8; #100;
A = 8'h50; B = 8'hC9; #100;
A = 8'h50; B = 8'hCA; #100;
A = 8'h50; B = 8'hCB; #100;
A = 8'h50; B = 8'hCC; #100;
A = 8'h50; B = 8'hCD; #100;
A = 8'h50; B = 8'hCE; #100;
A = 8'h50; B = 8'hCF; #100;
A = 8'h50; B = 8'hD0; #100;
A = 8'h50; B = 8'hD1; #100;
A = 8'h50; B = 8'hD2; #100;
A = 8'h50; B = 8'hD3; #100;
A = 8'h50; B = 8'hD4; #100;
A = 8'h50; B = 8'hD5; #100;
A = 8'h50; B = 8'hD6; #100;
A = 8'h50; B = 8'hD7; #100;
A = 8'h50; B = 8'hD8; #100;
A = 8'h50; B = 8'hD9; #100;
A = 8'h50; B = 8'hDA; #100;
A = 8'h50; B = 8'hDB; #100;
A = 8'h50; B = 8'hDC; #100;
A = 8'h50; B = 8'hDD; #100;
A = 8'h50; B = 8'hDE; #100;
A = 8'h50; B = 8'hDF; #100;
A = 8'h50; B = 8'hE0; #100;
A = 8'h50; B = 8'hE1; #100;
A = 8'h50; B = 8'hE2; #100;
A = 8'h50; B = 8'hE3; #100;
A = 8'h50; B = 8'hE4; #100;
A = 8'h50; B = 8'hE5; #100;
A = 8'h50; B = 8'hE6; #100;
A = 8'h50; B = 8'hE7; #100;
A = 8'h50; B = 8'hE8; #100;
A = 8'h50; B = 8'hE9; #100;
A = 8'h50; B = 8'hEA; #100;
A = 8'h50; B = 8'hEB; #100;
A = 8'h50; B = 8'hEC; #100;
A = 8'h50; B = 8'hED; #100;
A = 8'h50; B = 8'hEE; #100;
A = 8'h50; B = 8'hEF; #100;
A = 8'h50; B = 8'hF0; #100;
A = 8'h50; B = 8'hF1; #100;
A = 8'h50; B = 8'hF2; #100;
A = 8'h50; B = 8'hF3; #100;
A = 8'h50; B = 8'hF4; #100;
A = 8'h50; B = 8'hF5; #100;
A = 8'h50; B = 8'hF6; #100;
A = 8'h50; B = 8'hF7; #100;
A = 8'h50; B = 8'hF8; #100;
A = 8'h50; B = 8'hF9; #100;
A = 8'h50; B = 8'hFA; #100;
A = 8'h50; B = 8'hFB; #100;
A = 8'h50; B = 8'hFC; #100;
A = 8'h50; B = 8'hFD; #100;
A = 8'h50; B = 8'hFE; #100;
A = 8'h50; B = 8'hFF; #100;
A = 8'h51; B = 8'h0; #100;
A = 8'h51; B = 8'h1; #100;
A = 8'h51; B = 8'h2; #100;
A = 8'h51; B = 8'h3; #100;
A = 8'h51; B = 8'h4; #100;
A = 8'h51; B = 8'h5; #100;
A = 8'h51; B = 8'h6; #100;
A = 8'h51; B = 8'h7; #100;
A = 8'h51; B = 8'h8; #100;
A = 8'h51; B = 8'h9; #100;
A = 8'h51; B = 8'hA; #100;
A = 8'h51; B = 8'hB; #100;
A = 8'h51; B = 8'hC; #100;
A = 8'h51; B = 8'hD; #100;
A = 8'h51; B = 8'hE; #100;
A = 8'h51; B = 8'hF; #100;
A = 8'h51; B = 8'h10; #100;
A = 8'h51; B = 8'h11; #100;
A = 8'h51; B = 8'h12; #100;
A = 8'h51; B = 8'h13; #100;
A = 8'h51; B = 8'h14; #100;
A = 8'h51; B = 8'h15; #100;
A = 8'h51; B = 8'h16; #100;
A = 8'h51; B = 8'h17; #100;
A = 8'h51; B = 8'h18; #100;
A = 8'h51; B = 8'h19; #100;
A = 8'h51; B = 8'h1A; #100;
A = 8'h51; B = 8'h1B; #100;
A = 8'h51; B = 8'h1C; #100;
A = 8'h51; B = 8'h1D; #100;
A = 8'h51; B = 8'h1E; #100;
A = 8'h51; B = 8'h1F; #100;
A = 8'h51; B = 8'h20; #100;
A = 8'h51; B = 8'h21; #100;
A = 8'h51; B = 8'h22; #100;
A = 8'h51; B = 8'h23; #100;
A = 8'h51; B = 8'h24; #100;
A = 8'h51; B = 8'h25; #100;
A = 8'h51; B = 8'h26; #100;
A = 8'h51; B = 8'h27; #100;
A = 8'h51; B = 8'h28; #100;
A = 8'h51; B = 8'h29; #100;
A = 8'h51; B = 8'h2A; #100;
A = 8'h51; B = 8'h2B; #100;
A = 8'h51; B = 8'h2C; #100;
A = 8'h51; B = 8'h2D; #100;
A = 8'h51; B = 8'h2E; #100;
A = 8'h51; B = 8'h2F; #100;
A = 8'h51; B = 8'h30; #100;
A = 8'h51; B = 8'h31; #100;
A = 8'h51; B = 8'h32; #100;
A = 8'h51; B = 8'h33; #100;
A = 8'h51; B = 8'h34; #100;
A = 8'h51; B = 8'h35; #100;
A = 8'h51; B = 8'h36; #100;
A = 8'h51; B = 8'h37; #100;
A = 8'h51; B = 8'h38; #100;
A = 8'h51; B = 8'h39; #100;
A = 8'h51; B = 8'h3A; #100;
A = 8'h51; B = 8'h3B; #100;
A = 8'h51; B = 8'h3C; #100;
A = 8'h51; B = 8'h3D; #100;
A = 8'h51; B = 8'h3E; #100;
A = 8'h51; B = 8'h3F; #100;
A = 8'h51; B = 8'h40; #100;
A = 8'h51; B = 8'h41; #100;
A = 8'h51; B = 8'h42; #100;
A = 8'h51; B = 8'h43; #100;
A = 8'h51; B = 8'h44; #100;
A = 8'h51; B = 8'h45; #100;
A = 8'h51; B = 8'h46; #100;
A = 8'h51; B = 8'h47; #100;
A = 8'h51; B = 8'h48; #100;
A = 8'h51; B = 8'h49; #100;
A = 8'h51; B = 8'h4A; #100;
A = 8'h51; B = 8'h4B; #100;
A = 8'h51; B = 8'h4C; #100;
A = 8'h51; B = 8'h4D; #100;
A = 8'h51; B = 8'h4E; #100;
A = 8'h51; B = 8'h4F; #100;
A = 8'h51; B = 8'h50; #100;
A = 8'h51; B = 8'h51; #100;
A = 8'h51; B = 8'h52; #100;
A = 8'h51; B = 8'h53; #100;
A = 8'h51; B = 8'h54; #100;
A = 8'h51; B = 8'h55; #100;
A = 8'h51; B = 8'h56; #100;
A = 8'h51; B = 8'h57; #100;
A = 8'h51; B = 8'h58; #100;
A = 8'h51; B = 8'h59; #100;
A = 8'h51; B = 8'h5A; #100;
A = 8'h51; B = 8'h5B; #100;
A = 8'h51; B = 8'h5C; #100;
A = 8'h51; B = 8'h5D; #100;
A = 8'h51; B = 8'h5E; #100;
A = 8'h51; B = 8'h5F; #100;
A = 8'h51; B = 8'h60; #100;
A = 8'h51; B = 8'h61; #100;
A = 8'h51; B = 8'h62; #100;
A = 8'h51; B = 8'h63; #100;
A = 8'h51; B = 8'h64; #100;
A = 8'h51; B = 8'h65; #100;
A = 8'h51; B = 8'h66; #100;
A = 8'h51; B = 8'h67; #100;
A = 8'h51; B = 8'h68; #100;
A = 8'h51; B = 8'h69; #100;
A = 8'h51; B = 8'h6A; #100;
A = 8'h51; B = 8'h6B; #100;
A = 8'h51; B = 8'h6C; #100;
A = 8'h51; B = 8'h6D; #100;
A = 8'h51; B = 8'h6E; #100;
A = 8'h51; B = 8'h6F; #100;
A = 8'h51; B = 8'h70; #100;
A = 8'h51; B = 8'h71; #100;
A = 8'h51; B = 8'h72; #100;
A = 8'h51; B = 8'h73; #100;
A = 8'h51; B = 8'h74; #100;
A = 8'h51; B = 8'h75; #100;
A = 8'h51; B = 8'h76; #100;
A = 8'h51; B = 8'h77; #100;
A = 8'h51; B = 8'h78; #100;
A = 8'h51; B = 8'h79; #100;
A = 8'h51; B = 8'h7A; #100;
A = 8'h51; B = 8'h7B; #100;
A = 8'h51; B = 8'h7C; #100;
A = 8'h51; B = 8'h7D; #100;
A = 8'h51; B = 8'h7E; #100;
A = 8'h51; B = 8'h7F; #100;
A = 8'h51; B = 8'h80; #100;
A = 8'h51; B = 8'h81; #100;
A = 8'h51; B = 8'h82; #100;
A = 8'h51; B = 8'h83; #100;
A = 8'h51; B = 8'h84; #100;
A = 8'h51; B = 8'h85; #100;
A = 8'h51; B = 8'h86; #100;
A = 8'h51; B = 8'h87; #100;
A = 8'h51; B = 8'h88; #100;
A = 8'h51; B = 8'h89; #100;
A = 8'h51; B = 8'h8A; #100;
A = 8'h51; B = 8'h8B; #100;
A = 8'h51; B = 8'h8C; #100;
A = 8'h51; B = 8'h8D; #100;
A = 8'h51; B = 8'h8E; #100;
A = 8'h51; B = 8'h8F; #100;
A = 8'h51; B = 8'h90; #100;
A = 8'h51; B = 8'h91; #100;
A = 8'h51; B = 8'h92; #100;
A = 8'h51; B = 8'h93; #100;
A = 8'h51; B = 8'h94; #100;
A = 8'h51; B = 8'h95; #100;
A = 8'h51; B = 8'h96; #100;
A = 8'h51; B = 8'h97; #100;
A = 8'h51; B = 8'h98; #100;
A = 8'h51; B = 8'h99; #100;
A = 8'h51; B = 8'h9A; #100;
A = 8'h51; B = 8'h9B; #100;
A = 8'h51; B = 8'h9C; #100;
A = 8'h51; B = 8'h9D; #100;
A = 8'h51; B = 8'h9E; #100;
A = 8'h51; B = 8'h9F; #100;
A = 8'h51; B = 8'hA0; #100;
A = 8'h51; B = 8'hA1; #100;
A = 8'h51; B = 8'hA2; #100;
A = 8'h51; B = 8'hA3; #100;
A = 8'h51; B = 8'hA4; #100;
A = 8'h51; B = 8'hA5; #100;
A = 8'h51; B = 8'hA6; #100;
A = 8'h51; B = 8'hA7; #100;
A = 8'h51; B = 8'hA8; #100;
A = 8'h51; B = 8'hA9; #100;
A = 8'h51; B = 8'hAA; #100;
A = 8'h51; B = 8'hAB; #100;
A = 8'h51; B = 8'hAC; #100;
A = 8'h51; B = 8'hAD; #100;
A = 8'h51; B = 8'hAE; #100;
A = 8'h51; B = 8'hAF; #100;
A = 8'h51; B = 8'hB0; #100;
A = 8'h51; B = 8'hB1; #100;
A = 8'h51; B = 8'hB2; #100;
A = 8'h51; B = 8'hB3; #100;
A = 8'h51; B = 8'hB4; #100;
A = 8'h51; B = 8'hB5; #100;
A = 8'h51; B = 8'hB6; #100;
A = 8'h51; B = 8'hB7; #100;
A = 8'h51; B = 8'hB8; #100;
A = 8'h51; B = 8'hB9; #100;
A = 8'h51; B = 8'hBA; #100;
A = 8'h51; B = 8'hBB; #100;
A = 8'h51; B = 8'hBC; #100;
A = 8'h51; B = 8'hBD; #100;
A = 8'h51; B = 8'hBE; #100;
A = 8'h51; B = 8'hBF; #100;
A = 8'h51; B = 8'hC0; #100;
A = 8'h51; B = 8'hC1; #100;
A = 8'h51; B = 8'hC2; #100;
A = 8'h51; B = 8'hC3; #100;
A = 8'h51; B = 8'hC4; #100;
A = 8'h51; B = 8'hC5; #100;
A = 8'h51; B = 8'hC6; #100;
A = 8'h51; B = 8'hC7; #100;
A = 8'h51; B = 8'hC8; #100;
A = 8'h51; B = 8'hC9; #100;
A = 8'h51; B = 8'hCA; #100;
A = 8'h51; B = 8'hCB; #100;
A = 8'h51; B = 8'hCC; #100;
A = 8'h51; B = 8'hCD; #100;
A = 8'h51; B = 8'hCE; #100;
A = 8'h51; B = 8'hCF; #100;
A = 8'h51; B = 8'hD0; #100;
A = 8'h51; B = 8'hD1; #100;
A = 8'h51; B = 8'hD2; #100;
A = 8'h51; B = 8'hD3; #100;
A = 8'h51; B = 8'hD4; #100;
A = 8'h51; B = 8'hD5; #100;
A = 8'h51; B = 8'hD6; #100;
A = 8'h51; B = 8'hD7; #100;
A = 8'h51; B = 8'hD8; #100;
A = 8'h51; B = 8'hD9; #100;
A = 8'h51; B = 8'hDA; #100;
A = 8'h51; B = 8'hDB; #100;
A = 8'h51; B = 8'hDC; #100;
A = 8'h51; B = 8'hDD; #100;
A = 8'h51; B = 8'hDE; #100;
A = 8'h51; B = 8'hDF; #100;
A = 8'h51; B = 8'hE0; #100;
A = 8'h51; B = 8'hE1; #100;
A = 8'h51; B = 8'hE2; #100;
A = 8'h51; B = 8'hE3; #100;
A = 8'h51; B = 8'hE4; #100;
A = 8'h51; B = 8'hE5; #100;
A = 8'h51; B = 8'hE6; #100;
A = 8'h51; B = 8'hE7; #100;
A = 8'h51; B = 8'hE8; #100;
A = 8'h51; B = 8'hE9; #100;
A = 8'h51; B = 8'hEA; #100;
A = 8'h51; B = 8'hEB; #100;
A = 8'h51; B = 8'hEC; #100;
A = 8'h51; B = 8'hED; #100;
A = 8'h51; B = 8'hEE; #100;
A = 8'h51; B = 8'hEF; #100;
A = 8'h51; B = 8'hF0; #100;
A = 8'h51; B = 8'hF1; #100;
A = 8'h51; B = 8'hF2; #100;
A = 8'h51; B = 8'hF3; #100;
A = 8'h51; B = 8'hF4; #100;
A = 8'h51; B = 8'hF5; #100;
A = 8'h51; B = 8'hF6; #100;
A = 8'h51; B = 8'hF7; #100;
A = 8'h51; B = 8'hF8; #100;
A = 8'h51; B = 8'hF9; #100;
A = 8'h51; B = 8'hFA; #100;
A = 8'h51; B = 8'hFB; #100;
A = 8'h51; B = 8'hFC; #100;
A = 8'h51; B = 8'hFD; #100;
A = 8'h51; B = 8'hFE; #100;
A = 8'h51; B = 8'hFF; #100;
A = 8'h52; B = 8'h0; #100;
A = 8'h52; B = 8'h1; #100;
A = 8'h52; B = 8'h2; #100;
A = 8'h52; B = 8'h3; #100;
A = 8'h52; B = 8'h4; #100;
A = 8'h52; B = 8'h5; #100;
A = 8'h52; B = 8'h6; #100;
A = 8'h52; B = 8'h7; #100;
A = 8'h52; B = 8'h8; #100;
A = 8'h52; B = 8'h9; #100;
A = 8'h52; B = 8'hA; #100;
A = 8'h52; B = 8'hB; #100;
A = 8'h52; B = 8'hC; #100;
A = 8'h52; B = 8'hD; #100;
A = 8'h52; B = 8'hE; #100;
A = 8'h52; B = 8'hF; #100;
A = 8'h52; B = 8'h10; #100;
A = 8'h52; B = 8'h11; #100;
A = 8'h52; B = 8'h12; #100;
A = 8'h52; B = 8'h13; #100;
A = 8'h52; B = 8'h14; #100;
A = 8'h52; B = 8'h15; #100;
A = 8'h52; B = 8'h16; #100;
A = 8'h52; B = 8'h17; #100;
A = 8'h52; B = 8'h18; #100;
A = 8'h52; B = 8'h19; #100;
A = 8'h52; B = 8'h1A; #100;
A = 8'h52; B = 8'h1B; #100;
A = 8'h52; B = 8'h1C; #100;
A = 8'h52; B = 8'h1D; #100;
A = 8'h52; B = 8'h1E; #100;
A = 8'h52; B = 8'h1F; #100;
A = 8'h52; B = 8'h20; #100;
A = 8'h52; B = 8'h21; #100;
A = 8'h52; B = 8'h22; #100;
A = 8'h52; B = 8'h23; #100;
A = 8'h52; B = 8'h24; #100;
A = 8'h52; B = 8'h25; #100;
A = 8'h52; B = 8'h26; #100;
A = 8'h52; B = 8'h27; #100;
A = 8'h52; B = 8'h28; #100;
A = 8'h52; B = 8'h29; #100;
A = 8'h52; B = 8'h2A; #100;
A = 8'h52; B = 8'h2B; #100;
A = 8'h52; B = 8'h2C; #100;
A = 8'h52; B = 8'h2D; #100;
A = 8'h52; B = 8'h2E; #100;
A = 8'h52; B = 8'h2F; #100;
A = 8'h52; B = 8'h30; #100;
A = 8'h52; B = 8'h31; #100;
A = 8'h52; B = 8'h32; #100;
A = 8'h52; B = 8'h33; #100;
A = 8'h52; B = 8'h34; #100;
A = 8'h52; B = 8'h35; #100;
A = 8'h52; B = 8'h36; #100;
A = 8'h52; B = 8'h37; #100;
A = 8'h52; B = 8'h38; #100;
A = 8'h52; B = 8'h39; #100;
A = 8'h52; B = 8'h3A; #100;
A = 8'h52; B = 8'h3B; #100;
A = 8'h52; B = 8'h3C; #100;
A = 8'h52; B = 8'h3D; #100;
A = 8'h52; B = 8'h3E; #100;
A = 8'h52; B = 8'h3F; #100;
A = 8'h52; B = 8'h40; #100;
A = 8'h52; B = 8'h41; #100;
A = 8'h52; B = 8'h42; #100;
A = 8'h52; B = 8'h43; #100;
A = 8'h52; B = 8'h44; #100;
A = 8'h52; B = 8'h45; #100;
A = 8'h52; B = 8'h46; #100;
A = 8'h52; B = 8'h47; #100;
A = 8'h52; B = 8'h48; #100;
A = 8'h52; B = 8'h49; #100;
A = 8'h52; B = 8'h4A; #100;
A = 8'h52; B = 8'h4B; #100;
A = 8'h52; B = 8'h4C; #100;
A = 8'h52; B = 8'h4D; #100;
A = 8'h52; B = 8'h4E; #100;
A = 8'h52; B = 8'h4F; #100;
A = 8'h52; B = 8'h50; #100;
A = 8'h52; B = 8'h51; #100;
A = 8'h52; B = 8'h52; #100;
A = 8'h52; B = 8'h53; #100;
A = 8'h52; B = 8'h54; #100;
A = 8'h52; B = 8'h55; #100;
A = 8'h52; B = 8'h56; #100;
A = 8'h52; B = 8'h57; #100;
A = 8'h52; B = 8'h58; #100;
A = 8'h52; B = 8'h59; #100;
A = 8'h52; B = 8'h5A; #100;
A = 8'h52; B = 8'h5B; #100;
A = 8'h52; B = 8'h5C; #100;
A = 8'h52; B = 8'h5D; #100;
A = 8'h52; B = 8'h5E; #100;
A = 8'h52; B = 8'h5F; #100;
A = 8'h52; B = 8'h60; #100;
A = 8'h52; B = 8'h61; #100;
A = 8'h52; B = 8'h62; #100;
A = 8'h52; B = 8'h63; #100;
A = 8'h52; B = 8'h64; #100;
A = 8'h52; B = 8'h65; #100;
A = 8'h52; B = 8'h66; #100;
A = 8'h52; B = 8'h67; #100;
A = 8'h52; B = 8'h68; #100;
A = 8'h52; B = 8'h69; #100;
A = 8'h52; B = 8'h6A; #100;
A = 8'h52; B = 8'h6B; #100;
A = 8'h52; B = 8'h6C; #100;
A = 8'h52; B = 8'h6D; #100;
A = 8'h52; B = 8'h6E; #100;
A = 8'h52; B = 8'h6F; #100;
A = 8'h52; B = 8'h70; #100;
A = 8'h52; B = 8'h71; #100;
A = 8'h52; B = 8'h72; #100;
A = 8'h52; B = 8'h73; #100;
A = 8'h52; B = 8'h74; #100;
A = 8'h52; B = 8'h75; #100;
A = 8'h52; B = 8'h76; #100;
A = 8'h52; B = 8'h77; #100;
A = 8'h52; B = 8'h78; #100;
A = 8'h52; B = 8'h79; #100;
A = 8'h52; B = 8'h7A; #100;
A = 8'h52; B = 8'h7B; #100;
A = 8'h52; B = 8'h7C; #100;
A = 8'h52; B = 8'h7D; #100;
A = 8'h52; B = 8'h7E; #100;
A = 8'h52; B = 8'h7F; #100;
A = 8'h52; B = 8'h80; #100;
A = 8'h52; B = 8'h81; #100;
A = 8'h52; B = 8'h82; #100;
A = 8'h52; B = 8'h83; #100;
A = 8'h52; B = 8'h84; #100;
A = 8'h52; B = 8'h85; #100;
A = 8'h52; B = 8'h86; #100;
A = 8'h52; B = 8'h87; #100;
A = 8'h52; B = 8'h88; #100;
A = 8'h52; B = 8'h89; #100;
A = 8'h52; B = 8'h8A; #100;
A = 8'h52; B = 8'h8B; #100;
A = 8'h52; B = 8'h8C; #100;
A = 8'h52; B = 8'h8D; #100;
A = 8'h52; B = 8'h8E; #100;
A = 8'h52; B = 8'h8F; #100;
A = 8'h52; B = 8'h90; #100;
A = 8'h52; B = 8'h91; #100;
A = 8'h52; B = 8'h92; #100;
A = 8'h52; B = 8'h93; #100;
A = 8'h52; B = 8'h94; #100;
A = 8'h52; B = 8'h95; #100;
A = 8'h52; B = 8'h96; #100;
A = 8'h52; B = 8'h97; #100;
A = 8'h52; B = 8'h98; #100;
A = 8'h52; B = 8'h99; #100;
A = 8'h52; B = 8'h9A; #100;
A = 8'h52; B = 8'h9B; #100;
A = 8'h52; B = 8'h9C; #100;
A = 8'h52; B = 8'h9D; #100;
A = 8'h52; B = 8'h9E; #100;
A = 8'h52; B = 8'h9F; #100;
A = 8'h52; B = 8'hA0; #100;
A = 8'h52; B = 8'hA1; #100;
A = 8'h52; B = 8'hA2; #100;
A = 8'h52; B = 8'hA3; #100;
A = 8'h52; B = 8'hA4; #100;
A = 8'h52; B = 8'hA5; #100;
A = 8'h52; B = 8'hA6; #100;
A = 8'h52; B = 8'hA7; #100;
A = 8'h52; B = 8'hA8; #100;
A = 8'h52; B = 8'hA9; #100;
A = 8'h52; B = 8'hAA; #100;
A = 8'h52; B = 8'hAB; #100;
A = 8'h52; B = 8'hAC; #100;
A = 8'h52; B = 8'hAD; #100;
A = 8'h52; B = 8'hAE; #100;
A = 8'h52; B = 8'hAF; #100;
A = 8'h52; B = 8'hB0; #100;
A = 8'h52; B = 8'hB1; #100;
A = 8'h52; B = 8'hB2; #100;
A = 8'h52; B = 8'hB3; #100;
A = 8'h52; B = 8'hB4; #100;
A = 8'h52; B = 8'hB5; #100;
A = 8'h52; B = 8'hB6; #100;
A = 8'h52; B = 8'hB7; #100;
A = 8'h52; B = 8'hB8; #100;
A = 8'h52; B = 8'hB9; #100;
A = 8'h52; B = 8'hBA; #100;
A = 8'h52; B = 8'hBB; #100;
A = 8'h52; B = 8'hBC; #100;
A = 8'h52; B = 8'hBD; #100;
A = 8'h52; B = 8'hBE; #100;
A = 8'h52; B = 8'hBF; #100;
A = 8'h52; B = 8'hC0; #100;
A = 8'h52; B = 8'hC1; #100;
A = 8'h52; B = 8'hC2; #100;
A = 8'h52; B = 8'hC3; #100;
A = 8'h52; B = 8'hC4; #100;
A = 8'h52; B = 8'hC5; #100;
A = 8'h52; B = 8'hC6; #100;
A = 8'h52; B = 8'hC7; #100;
A = 8'h52; B = 8'hC8; #100;
A = 8'h52; B = 8'hC9; #100;
A = 8'h52; B = 8'hCA; #100;
A = 8'h52; B = 8'hCB; #100;
A = 8'h52; B = 8'hCC; #100;
A = 8'h52; B = 8'hCD; #100;
A = 8'h52; B = 8'hCE; #100;
A = 8'h52; B = 8'hCF; #100;
A = 8'h52; B = 8'hD0; #100;
A = 8'h52; B = 8'hD1; #100;
A = 8'h52; B = 8'hD2; #100;
A = 8'h52; B = 8'hD3; #100;
A = 8'h52; B = 8'hD4; #100;
A = 8'h52; B = 8'hD5; #100;
A = 8'h52; B = 8'hD6; #100;
A = 8'h52; B = 8'hD7; #100;
A = 8'h52; B = 8'hD8; #100;
A = 8'h52; B = 8'hD9; #100;
A = 8'h52; B = 8'hDA; #100;
A = 8'h52; B = 8'hDB; #100;
A = 8'h52; B = 8'hDC; #100;
A = 8'h52; B = 8'hDD; #100;
A = 8'h52; B = 8'hDE; #100;
A = 8'h52; B = 8'hDF; #100;
A = 8'h52; B = 8'hE0; #100;
A = 8'h52; B = 8'hE1; #100;
A = 8'h52; B = 8'hE2; #100;
A = 8'h52; B = 8'hE3; #100;
A = 8'h52; B = 8'hE4; #100;
A = 8'h52; B = 8'hE5; #100;
A = 8'h52; B = 8'hE6; #100;
A = 8'h52; B = 8'hE7; #100;
A = 8'h52; B = 8'hE8; #100;
A = 8'h52; B = 8'hE9; #100;
A = 8'h52; B = 8'hEA; #100;
A = 8'h52; B = 8'hEB; #100;
A = 8'h52; B = 8'hEC; #100;
A = 8'h52; B = 8'hED; #100;
A = 8'h52; B = 8'hEE; #100;
A = 8'h52; B = 8'hEF; #100;
A = 8'h52; B = 8'hF0; #100;
A = 8'h52; B = 8'hF1; #100;
A = 8'h52; B = 8'hF2; #100;
A = 8'h52; B = 8'hF3; #100;
A = 8'h52; B = 8'hF4; #100;
A = 8'h52; B = 8'hF5; #100;
A = 8'h52; B = 8'hF6; #100;
A = 8'h52; B = 8'hF7; #100;
A = 8'h52; B = 8'hF8; #100;
A = 8'h52; B = 8'hF9; #100;
A = 8'h52; B = 8'hFA; #100;
A = 8'h52; B = 8'hFB; #100;
A = 8'h52; B = 8'hFC; #100;
A = 8'h52; B = 8'hFD; #100;
A = 8'h52; B = 8'hFE; #100;
A = 8'h52; B = 8'hFF; #100;
A = 8'h53; B = 8'h0; #100;
A = 8'h53; B = 8'h1; #100;
A = 8'h53; B = 8'h2; #100;
A = 8'h53; B = 8'h3; #100;
A = 8'h53; B = 8'h4; #100;
A = 8'h53; B = 8'h5; #100;
A = 8'h53; B = 8'h6; #100;
A = 8'h53; B = 8'h7; #100;
A = 8'h53; B = 8'h8; #100;
A = 8'h53; B = 8'h9; #100;
A = 8'h53; B = 8'hA; #100;
A = 8'h53; B = 8'hB; #100;
A = 8'h53; B = 8'hC; #100;
A = 8'h53; B = 8'hD; #100;
A = 8'h53; B = 8'hE; #100;
A = 8'h53; B = 8'hF; #100;
A = 8'h53; B = 8'h10; #100;
A = 8'h53; B = 8'h11; #100;
A = 8'h53; B = 8'h12; #100;
A = 8'h53; B = 8'h13; #100;
A = 8'h53; B = 8'h14; #100;
A = 8'h53; B = 8'h15; #100;
A = 8'h53; B = 8'h16; #100;
A = 8'h53; B = 8'h17; #100;
A = 8'h53; B = 8'h18; #100;
A = 8'h53; B = 8'h19; #100;
A = 8'h53; B = 8'h1A; #100;
A = 8'h53; B = 8'h1B; #100;
A = 8'h53; B = 8'h1C; #100;
A = 8'h53; B = 8'h1D; #100;
A = 8'h53; B = 8'h1E; #100;
A = 8'h53; B = 8'h1F; #100;
A = 8'h53; B = 8'h20; #100;
A = 8'h53; B = 8'h21; #100;
A = 8'h53; B = 8'h22; #100;
A = 8'h53; B = 8'h23; #100;
A = 8'h53; B = 8'h24; #100;
A = 8'h53; B = 8'h25; #100;
A = 8'h53; B = 8'h26; #100;
A = 8'h53; B = 8'h27; #100;
A = 8'h53; B = 8'h28; #100;
A = 8'h53; B = 8'h29; #100;
A = 8'h53; B = 8'h2A; #100;
A = 8'h53; B = 8'h2B; #100;
A = 8'h53; B = 8'h2C; #100;
A = 8'h53; B = 8'h2D; #100;
A = 8'h53; B = 8'h2E; #100;
A = 8'h53; B = 8'h2F; #100;
A = 8'h53; B = 8'h30; #100;
A = 8'h53; B = 8'h31; #100;
A = 8'h53; B = 8'h32; #100;
A = 8'h53; B = 8'h33; #100;
A = 8'h53; B = 8'h34; #100;
A = 8'h53; B = 8'h35; #100;
A = 8'h53; B = 8'h36; #100;
A = 8'h53; B = 8'h37; #100;
A = 8'h53; B = 8'h38; #100;
A = 8'h53; B = 8'h39; #100;
A = 8'h53; B = 8'h3A; #100;
A = 8'h53; B = 8'h3B; #100;
A = 8'h53; B = 8'h3C; #100;
A = 8'h53; B = 8'h3D; #100;
A = 8'h53; B = 8'h3E; #100;
A = 8'h53; B = 8'h3F; #100;
A = 8'h53; B = 8'h40; #100;
A = 8'h53; B = 8'h41; #100;
A = 8'h53; B = 8'h42; #100;
A = 8'h53; B = 8'h43; #100;
A = 8'h53; B = 8'h44; #100;
A = 8'h53; B = 8'h45; #100;
A = 8'h53; B = 8'h46; #100;
A = 8'h53; B = 8'h47; #100;
A = 8'h53; B = 8'h48; #100;
A = 8'h53; B = 8'h49; #100;
A = 8'h53; B = 8'h4A; #100;
A = 8'h53; B = 8'h4B; #100;
A = 8'h53; B = 8'h4C; #100;
A = 8'h53; B = 8'h4D; #100;
A = 8'h53; B = 8'h4E; #100;
A = 8'h53; B = 8'h4F; #100;
A = 8'h53; B = 8'h50; #100;
A = 8'h53; B = 8'h51; #100;
A = 8'h53; B = 8'h52; #100;
A = 8'h53; B = 8'h53; #100;
A = 8'h53; B = 8'h54; #100;
A = 8'h53; B = 8'h55; #100;
A = 8'h53; B = 8'h56; #100;
A = 8'h53; B = 8'h57; #100;
A = 8'h53; B = 8'h58; #100;
A = 8'h53; B = 8'h59; #100;
A = 8'h53; B = 8'h5A; #100;
A = 8'h53; B = 8'h5B; #100;
A = 8'h53; B = 8'h5C; #100;
A = 8'h53; B = 8'h5D; #100;
A = 8'h53; B = 8'h5E; #100;
A = 8'h53; B = 8'h5F; #100;
A = 8'h53; B = 8'h60; #100;
A = 8'h53; B = 8'h61; #100;
A = 8'h53; B = 8'h62; #100;
A = 8'h53; B = 8'h63; #100;
A = 8'h53; B = 8'h64; #100;
A = 8'h53; B = 8'h65; #100;
A = 8'h53; B = 8'h66; #100;
A = 8'h53; B = 8'h67; #100;
A = 8'h53; B = 8'h68; #100;
A = 8'h53; B = 8'h69; #100;
A = 8'h53; B = 8'h6A; #100;
A = 8'h53; B = 8'h6B; #100;
A = 8'h53; B = 8'h6C; #100;
A = 8'h53; B = 8'h6D; #100;
A = 8'h53; B = 8'h6E; #100;
A = 8'h53; B = 8'h6F; #100;
A = 8'h53; B = 8'h70; #100;
A = 8'h53; B = 8'h71; #100;
A = 8'h53; B = 8'h72; #100;
A = 8'h53; B = 8'h73; #100;
A = 8'h53; B = 8'h74; #100;
A = 8'h53; B = 8'h75; #100;
A = 8'h53; B = 8'h76; #100;
A = 8'h53; B = 8'h77; #100;
A = 8'h53; B = 8'h78; #100;
A = 8'h53; B = 8'h79; #100;
A = 8'h53; B = 8'h7A; #100;
A = 8'h53; B = 8'h7B; #100;
A = 8'h53; B = 8'h7C; #100;
A = 8'h53; B = 8'h7D; #100;
A = 8'h53; B = 8'h7E; #100;
A = 8'h53; B = 8'h7F; #100;
A = 8'h53; B = 8'h80; #100;
A = 8'h53; B = 8'h81; #100;
A = 8'h53; B = 8'h82; #100;
A = 8'h53; B = 8'h83; #100;
A = 8'h53; B = 8'h84; #100;
A = 8'h53; B = 8'h85; #100;
A = 8'h53; B = 8'h86; #100;
A = 8'h53; B = 8'h87; #100;
A = 8'h53; B = 8'h88; #100;
A = 8'h53; B = 8'h89; #100;
A = 8'h53; B = 8'h8A; #100;
A = 8'h53; B = 8'h8B; #100;
A = 8'h53; B = 8'h8C; #100;
A = 8'h53; B = 8'h8D; #100;
A = 8'h53; B = 8'h8E; #100;
A = 8'h53; B = 8'h8F; #100;
A = 8'h53; B = 8'h90; #100;
A = 8'h53; B = 8'h91; #100;
A = 8'h53; B = 8'h92; #100;
A = 8'h53; B = 8'h93; #100;
A = 8'h53; B = 8'h94; #100;
A = 8'h53; B = 8'h95; #100;
A = 8'h53; B = 8'h96; #100;
A = 8'h53; B = 8'h97; #100;
A = 8'h53; B = 8'h98; #100;
A = 8'h53; B = 8'h99; #100;
A = 8'h53; B = 8'h9A; #100;
A = 8'h53; B = 8'h9B; #100;
A = 8'h53; B = 8'h9C; #100;
A = 8'h53; B = 8'h9D; #100;
A = 8'h53; B = 8'h9E; #100;
A = 8'h53; B = 8'h9F; #100;
A = 8'h53; B = 8'hA0; #100;
A = 8'h53; B = 8'hA1; #100;
A = 8'h53; B = 8'hA2; #100;
A = 8'h53; B = 8'hA3; #100;
A = 8'h53; B = 8'hA4; #100;
A = 8'h53; B = 8'hA5; #100;
A = 8'h53; B = 8'hA6; #100;
A = 8'h53; B = 8'hA7; #100;
A = 8'h53; B = 8'hA8; #100;
A = 8'h53; B = 8'hA9; #100;
A = 8'h53; B = 8'hAA; #100;
A = 8'h53; B = 8'hAB; #100;
A = 8'h53; B = 8'hAC; #100;
A = 8'h53; B = 8'hAD; #100;
A = 8'h53; B = 8'hAE; #100;
A = 8'h53; B = 8'hAF; #100;
A = 8'h53; B = 8'hB0; #100;
A = 8'h53; B = 8'hB1; #100;
A = 8'h53; B = 8'hB2; #100;
A = 8'h53; B = 8'hB3; #100;
A = 8'h53; B = 8'hB4; #100;
A = 8'h53; B = 8'hB5; #100;
A = 8'h53; B = 8'hB6; #100;
A = 8'h53; B = 8'hB7; #100;
A = 8'h53; B = 8'hB8; #100;
A = 8'h53; B = 8'hB9; #100;
A = 8'h53; B = 8'hBA; #100;
A = 8'h53; B = 8'hBB; #100;
A = 8'h53; B = 8'hBC; #100;
A = 8'h53; B = 8'hBD; #100;
A = 8'h53; B = 8'hBE; #100;
A = 8'h53; B = 8'hBF; #100;
A = 8'h53; B = 8'hC0; #100;
A = 8'h53; B = 8'hC1; #100;
A = 8'h53; B = 8'hC2; #100;
A = 8'h53; B = 8'hC3; #100;
A = 8'h53; B = 8'hC4; #100;
A = 8'h53; B = 8'hC5; #100;
A = 8'h53; B = 8'hC6; #100;
A = 8'h53; B = 8'hC7; #100;
A = 8'h53; B = 8'hC8; #100;
A = 8'h53; B = 8'hC9; #100;
A = 8'h53; B = 8'hCA; #100;
A = 8'h53; B = 8'hCB; #100;
A = 8'h53; B = 8'hCC; #100;
A = 8'h53; B = 8'hCD; #100;
A = 8'h53; B = 8'hCE; #100;
A = 8'h53; B = 8'hCF; #100;
A = 8'h53; B = 8'hD0; #100;
A = 8'h53; B = 8'hD1; #100;
A = 8'h53; B = 8'hD2; #100;
A = 8'h53; B = 8'hD3; #100;
A = 8'h53; B = 8'hD4; #100;
A = 8'h53; B = 8'hD5; #100;
A = 8'h53; B = 8'hD6; #100;
A = 8'h53; B = 8'hD7; #100;
A = 8'h53; B = 8'hD8; #100;
A = 8'h53; B = 8'hD9; #100;
A = 8'h53; B = 8'hDA; #100;
A = 8'h53; B = 8'hDB; #100;
A = 8'h53; B = 8'hDC; #100;
A = 8'h53; B = 8'hDD; #100;
A = 8'h53; B = 8'hDE; #100;
A = 8'h53; B = 8'hDF; #100;
A = 8'h53; B = 8'hE0; #100;
A = 8'h53; B = 8'hE1; #100;
A = 8'h53; B = 8'hE2; #100;
A = 8'h53; B = 8'hE3; #100;
A = 8'h53; B = 8'hE4; #100;
A = 8'h53; B = 8'hE5; #100;
A = 8'h53; B = 8'hE6; #100;
A = 8'h53; B = 8'hE7; #100;
A = 8'h53; B = 8'hE8; #100;
A = 8'h53; B = 8'hE9; #100;
A = 8'h53; B = 8'hEA; #100;
A = 8'h53; B = 8'hEB; #100;
A = 8'h53; B = 8'hEC; #100;
A = 8'h53; B = 8'hED; #100;
A = 8'h53; B = 8'hEE; #100;
A = 8'h53; B = 8'hEF; #100;
A = 8'h53; B = 8'hF0; #100;
A = 8'h53; B = 8'hF1; #100;
A = 8'h53; B = 8'hF2; #100;
A = 8'h53; B = 8'hF3; #100;
A = 8'h53; B = 8'hF4; #100;
A = 8'h53; B = 8'hF5; #100;
A = 8'h53; B = 8'hF6; #100;
A = 8'h53; B = 8'hF7; #100;
A = 8'h53; B = 8'hF8; #100;
A = 8'h53; B = 8'hF9; #100;
A = 8'h53; B = 8'hFA; #100;
A = 8'h53; B = 8'hFB; #100;
A = 8'h53; B = 8'hFC; #100;
A = 8'h53; B = 8'hFD; #100;
A = 8'h53; B = 8'hFE; #100;
A = 8'h53; B = 8'hFF; #100;
A = 8'h54; B = 8'h0; #100;
A = 8'h54; B = 8'h1; #100;
A = 8'h54; B = 8'h2; #100;
A = 8'h54; B = 8'h3; #100;
A = 8'h54; B = 8'h4; #100;
A = 8'h54; B = 8'h5; #100;
A = 8'h54; B = 8'h6; #100;
A = 8'h54; B = 8'h7; #100;
A = 8'h54; B = 8'h8; #100;
A = 8'h54; B = 8'h9; #100;
A = 8'h54; B = 8'hA; #100;
A = 8'h54; B = 8'hB; #100;
A = 8'h54; B = 8'hC; #100;
A = 8'h54; B = 8'hD; #100;
A = 8'h54; B = 8'hE; #100;
A = 8'h54; B = 8'hF; #100;
A = 8'h54; B = 8'h10; #100;
A = 8'h54; B = 8'h11; #100;
A = 8'h54; B = 8'h12; #100;
A = 8'h54; B = 8'h13; #100;
A = 8'h54; B = 8'h14; #100;
A = 8'h54; B = 8'h15; #100;
A = 8'h54; B = 8'h16; #100;
A = 8'h54; B = 8'h17; #100;
A = 8'h54; B = 8'h18; #100;
A = 8'h54; B = 8'h19; #100;
A = 8'h54; B = 8'h1A; #100;
A = 8'h54; B = 8'h1B; #100;
A = 8'h54; B = 8'h1C; #100;
A = 8'h54; B = 8'h1D; #100;
A = 8'h54; B = 8'h1E; #100;
A = 8'h54; B = 8'h1F; #100;
A = 8'h54; B = 8'h20; #100;
A = 8'h54; B = 8'h21; #100;
A = 8'h54; B = 8'h22; #100;
A = 8'h54; B = 8'h23; #100;
A = 8'h54; B = 8'h24; #100;
A = 8'h54; B = 8'h25; #100;
A = 8'h54; B = 8'h26; #100;
A = 8'h54; B = 8'h27; #100;
A = 8'h54; B = 8'h28; #100;
A = 8'h54; B = 8'h29; #100;
A = 8'h54; B = 8'h2A; #100;
A = 8'h54; B = 8'h2B; #100;
A = 8'h54; B = 8'h2C; #100;
A = 8'h54; B = 8'h2D; #100;
A = 8'h54; B = 8'h2E; #100;
A = 8'h54; B = 8'h2F; #100;
A = 8'h54; B = 8'h30; #100;
A = 8'h54; B = 8'h31; #100;
A = 8'h54; B = 8'h32; #100;
A = 8'h54; B = 8'h33; #100;
A = 8'h54; B = 8'h34; #100;
A = 8'h54; B = 8'h35; #100;
A = 8'h54; B = 8'h36; #100;
A = 8'h54; B = 8'h37; #100;
A = 8'h54; B = 8'h38; #100;
A = 8'h54; B = 8'h39; #100;
A = 8'h54; B = 8'h3A; #100;
A = 8'h54; B = 8'h3B; #100;
A = 8'h54; B = 8'h3C; #100;
A = 8'h54; B = 8'h3D; #100;
A = 8'h54; B = 8'h3E; #100;
A = 8'h54; B = 8'h3F; #100;
A = 8'h54; B = 8'h40; #100;
A = 8'h54; B = 8'h41; #100;
A = 8'h54; B = 8'h42; #100;
A = 8'h54; B = 8'h43; #100;
A = 8'h54; B = 8'h44; #100;
A = 8'h54; B = 8'h45; #100;
A = 8'h54; B = 8'h46; #100;
A = 8'h54; B = 8'h47; #100;
A = 8'h54; B = 8'h48; #100;
A = 8'h54; B = 8'h49; #100;
A = 8'h54; B = 8'h4A; #100;
A = 8'h54; B = 8'h4B; #100;
A = 8'h54; B = 8'h4C; #100;
A = 8'h54; B = 8'h4D; #100;
A = 8'h54; B = 8'h4E; #100;
A = 8'h54; B = 8'h4F; #100;
A = 8'h54; B = 8'h50; #100;
A = 8'h54; B = 8'h51; #100;
A = 8'h54; B = 8'h52; #100;
A = 8'h54; B = 8'h53; #100;
A = 8'h54; B = 8'h54; #100;
A = 8'h54; B = 8'h55; #100;
A = 8'h54; B = 8'h56; #100;
A = 8'h54; B = 8'h57; #100;
A = 8'h54; B = 8'h58; #100;
A = 8'h54; B = 8'h59; #100;
A = 8'h54; B = 8'h5A; #100;
A = 8'h54; B = 8'h5B; #100;
A = 8'h54; B = 8'h5C; #100;
A = 8'h54; B = 8'h5D; #100;
A = 8'h54; B = 8'h5E; #100;
A = 8'h54; B = 8'h5F; #100;
A = 8'h54; B = 8'h60; #100;
A = 8'h54; B = 8'h61; #100;
A = 8'h54; B = 8'h62; #100;
A = 8'h54; B = 8'h63; #100;
A = 8'h54; B = 8'h64; #100;
A = 8'h54; B = 8'h65; #100;
A = 8'h54; B = 8'h66; #100;
A = 8'h54; B = 8'h67; #100;
A = 8'h54; B = 8'h68; #100;
A = 8'h54; B = 8'h69; #100;
A = 8'h54; B = 8'h6A; #100;
A = 8'h54; B = 8'h6B; #100;
A = 8'h54; B = 8'h6C; #100;
A = 8'h54; B = 8'h6D; #100;
A = 8'h54; B = 8'h6E; #100;
A = 8'h54; B = 8'h6F; #100;
A = 8'h54; B = 8'h70; #100;
A = 8'h54; B = 8'h71; #100;
A = 8'h54; B = 8'h72; #100;
A = 8'h54; B = 8'h73; #100;
A = 8'h54; B = 8'h74; #100;
A = 8'h54; B = 8'h75; #100;
A = 8'h54; B = 8'h76; #100;
A = 8'h54; B = 8'h77; #100;
A = 8'h54; B = 8'h78; #100;
A = 8'h54; B = 8'h79; #100;
A = 8'h54; B = 8'h7A; #100;
A = 8'h54; B = 8'h7B; #100;
A = 8'h54; B = 8'h7C; #100;
A = 8'h54; B = 8'h7D; #100;
A = 8'h54; B = 8'h7E; #100;
A = 8'h54; B = 8'h7F; #100;
A = 8'h54; B = 8'h80; #100;
A = 8'h54; B = 8'h81; #100;
A = 8'h54; B = 8'h82; #100;
A = 8'h54; B = 8'h83; #100;
A = 8'h54; B = 8'h84; #100;
A = 8'h54; B = 8'h85; #100;
A = 8'h54; B = 8'h86; #100;
A = 8'h54; B = 8'h87; #100;
A = 8'h54; B = 8'h88; #100;
A = 8'h54; B = 8'h89; #100;
A = 8'h54; B = 8'h8A; #100;
A = 8'h54; B = 8'h8B; #100;
A = 8'h54; B = 8'h8C; #100;
A = 8'h54; B = 8'h8D; #100;
A = 8'h54; B = 8'h8E; #100;
A = 8'h54; B = 8'h8F; #100;
A = 8'h54; B = 8'h90; #100;
A = 8'h54; B = 8'h91; #100;
A = 8'h54; B = 8'h92; #100;
A = 8'h54; B = 8'h93; #100;
A = 8'h54; B = 8'h94; #100;
A = 8'h54; B = 8'h95; #100;
A = 8'h54; B = 8'h96; #100;
A = 8'h54; B = 8'h97; #100;
A = 8'h54; B = 8'h98; #100;
A = 8'h54; B = 8'h99; #100;
A = 8'h54; B = 8'h9A; #100;
A = 8'h54; B = 8'h9B; #100;
A = 8'h54; B = 8'h9C; #100;
A = 8'h54; B = 8'h9D; #100;
A = 8'h54; B = 8'h9E; #100;
A = 8'h54; B = 8'h9F; #100;
A = 8'h54; B = 8'hA0; #100;
A = 8'h54; B = 8'hA1; #100;
A = 8'h54; B = 8'hA2; #100;
A = 8'h54; B = 8'hA3; #100;
A = 8'h54; B = 8'hA4; #100;
A = 8'h54; B = 8'hA5; #100;
A = 8'h54; B = 8'hA6; #100;
A = 8'h54; B = 8'hA7; #100;
A = 8'h54; B = 8'hA8; #100;
A = 8'h54; B = 8'hA9; #100;
A = 8'h54; B = 8'hAA; #100;
A = 8'h54; B = 8'hAB; #100;
A = 8'h54; B = 8'hAC; #100;
A = 8'h54; B = 8'hAD; #100;
A = 8'h54; B = 8'hAE; #100;
A = 8'h54; B = 8'hAF; #100;
A = 8'h54; B = 8'hB0; #100;
A = 8'h54; B = 8'hB1; #100;
A = 8'h54; B = 8'hB2; #100;
A = 8'h54; B = 8'hB3; #100;
A = 8'h54; B = 8'hB4; #100;
A = 8'h54; B = 8'hB5; #100;
A = 8'h54; B = 8'hB6; #100;
A = 8'h54; B = 8'hB7; #100;
A = 8'h54; B = 8'hB8; #100;
A = 8'h54; B = 8'hB9; #100;
A = 8'h54; B = 8'hBA; #100;
A = 8'h54; B = 8'hBB; #100;
A = 8'h54; B = 8'hBC; #100;
A = 8'h54; B = 8'hBD; #100;
A = 8'h54; B = 8'hBE; #100;
A = 8'h54; B = 8'hBF; #100;
A = 8'h54; B = 8'hC0; #100;
A = 8'h54; B = 8'hC1; #100;
A = 8'h54; B = 8'hC2; #100;
A = 8'h54; B = 8'hC3; #100;
A = 8'h54; B = 8'hC4; #100;
A = 8'h54; B = 8'hC5; #100;
A = 8'h54; B = 8'hC6; #100;
A = 8'h54; B = 8'hC7; #100;
A = 8'h54; B = 8'hC8; #100;
A = 8'h54; B = 8'hC9; #100;
A = 8'h54; B = 8'hCA; #100;
A = 8'h54; B = 8'hCB; #100;
A = 8'h54; B = 8'hCC; #100;
A = 8'h54; B = 8'hCD; #100;
A = 8'h54; B = 8'hCE; #100;
A = 8'h54; B = 8'hCF; #100;
A = 8'h54; B = 8'hD0; #100;
A = 8'h54; B = 8'hD1; #100;
A = 8'h54; B = 8'hD2; #100;
A = 8'h54; B = 8'hD3; #100;
A = 8'h54; B = 8'hD4; #100;
A = 8'h54; B = 8'hD5; #100;
A = 8'h54; B = 8'hD6; #100;
A = 8'h54; B = 8'hD7; #100;
A = 8'h54; B = 8'hD8; #100;
A = 8'h54; B = 8'hD9; #100;
A = 8'h54; B = 8'hDA; #100;
A = 8'h54; B = 8'hDB; #100;
A = 8'h54; B = 8'hDC; #100;
A = 8'h54; B = 8'hDD; #100;
A = 8'h54; B = 8'hDE; #100;
A = 8'h54; B = 8'hDF; #100;
A = 8'h54; B = 8'hE0; #100;
A = 8'h54; B = 8'hE1; #100;
A = 8'h54; B = 8'hE2; #100;
A = 8'h54; B = 8'hE3; #100;
A = 8'h54; B = 8'hE4; #100;
A = 8'h54; B = 8'hE5; #100;
A = 8'h54; B = 8'hE6; #100;
A = 8'h54; B = 8'hE7; #100;
A = 8'h54; B = 8'hE8; #100;
A = 8'h54; B = 8'hE9; #100;
A = 8'h54; B = 8'hEA; #100;
A = 8'h54; B = 8'hEB; #100;
A = 8'h54; B = 8'hEC; #100;
A = 8'h54; B = 8'hED; #100;
A = 8'h54; B = 8'hEE; #100;
A = 8'h54; B = 8'hEF; #100;
A = 8'h54; B = 8'hF0; #100;
A = 8'h54; B = 8'hF1; #100;
A = 8'h54; B = 8'hF2; #100;
A = 8'h54; B = 8'hF3; #100;
A = 8'h54; B = 8'hF4; #100;
A = 8'h54; B = 8'hF5; #100;
A = 8'h54; B = 8'hF6; #100;
A = 8'h54; B = 8'hF7; #100;
A = 8'h54; B = 8'hF8; #100;
A = 8'h54; B = 8'hF9; #100;
A = 8'h54; B = 8'hFA; #100;
A = 8'h54; B = 8'hFB; #100;
A = 8'h54; B = 8'hFC; #100;
A = 8'h54; B = 8'hFD; #100;
A = 8'h54; B = 8'hFE; #100;
A = 8'h54; B = 8'hFF; #100;
A = 8'h55; B = 8'h0; #100;
A = 8'h55; B = 8'h1; #100;
A = 8'h55; B = 8'h2; #100;
A = 8'h55; B = 8'h3; #100;
A = 8'h55; B = 8'h4; #100;
A = 8'h55; B = 8'h5; #100;
A = 8'h55; B = 8'h6; #100;
A = 8'h55; B = 8'h7; #100;
A = 8'h55; B = 8'h8; #100;
A = 8'h55; B = 8'h9; #100;
A = 8'h55; B = 8'hA; #100;
A = 8'h55; B = 8'hB; #100;
A = 8'h55; B = 8'hC; #100;
A = 8'h55; B = 8'hD; #100;
A = 8'h55; B = 8'hE; #100;
A = 8'h55; B = 8'hF; #100;
A = 8'h55; B = 8'h10; #100;
A = 8'h55; B = 8'h11; #100;
A = 8'h55; B = 8'h12; #100;
A = 8'h55; B = 8'h13; #100;
A = 8'h55; B = 8'h14; #100;
A = 8'h55; B = 8'h15; #100;
A = 8'h55; B = 8'h16; #100;
A = 8'h55; B = 8'h17; #100;
A = 8'h55; B = 8'h18; #100;
A = 8'h55; B = 8'h19; #100;
A = 8'h55; B = 8'h1A; #100;
A = 8'h55; B = 8'h1B; #100;
A = 8'h55; B = 8'h1C; #100;
A = 8'h55; B = 8'h1D; #100;
A = 8'h55; B = 8'h1E; #100;
A = 8'h55; B = 8'h1F; #100;
A = 8'h55; B = 8'h20; #100;
A = 8'h55; B = 8'h21; #100;
A = 8'h55; B = 8'h22; #100;
A = 8'h55; B = 8'h23; #100;
A = 8'h55; B = 8'h24; #100;
A = 8'h55; B = 8'h25; #100;
A = 8'h55; B = 8'h26; #100;
A = 8'h55; B = 8'h27; #100;
A = 8'h55; B = 8'h28; #100;
A = 8'h55; B = 8'h29; #100;
A = 8'h55; B = 8'h2A; #100;
A = 8'h55; B = 8'h2B; #100;
A = 8'h55; B = 8'h2C; #100;
A = 8'h55; B = 8'h2D; #100;
A = 8'h55; B = 8'h2E; #100;
A = 8'h55; B = 8'h2F; #100;
A = 8'h55; B = 8'h30; #100;
A = 8'h55; B = 8'h31; #100;
A = 8'h55; B = 8'h32; #100;
A = 8'h55; B = 8'h33; #100;
A = 8'h55; B = 8'h34; #100;
A = 8'h55; B = 8'h35; #100;
A = 8'h55; B = 8'h36; #100;
A = 8'h55; B = 8'h37; #100;
A = 8'h55; B = 8'h38; #100;
A = 8'h55; B = 8'h39; #100;
A = 8'h55; B = 8'h3A; #100;
A = 8'h55; B = 8'h3B; #100;
A = 8'h55; B = 8'h3C; #100;
A = 8'h55; B = 8'h3D; #100;
A = 8'h55; B = 8'h3E; #100;
A = 8'h55; B = 8'h3F; #100;
A = 8'h55; B = 8'h40; #100;
A = 8'h55; B = 8'h41; #100;
A = 8'h55; B = 8'h42; #100;
A = 8'h55; B = 8'h43; #100;
A = 8'h55; B = 8'h44; #100;
A = 8'h55; B = 8'h45; #100;
A = 8'h55; B = 8'h46; #100;
A = 8'h55; B = 8'h47; #100;
A = 8'h55; B = 8'h48; #100;
A = 8'h55; B = 8'h49; #100;
A = 8'h55; B = 8'h4A; #100;
A = 8'h55; B = 8'h4B; #100;
A = 8'h55; B = 8'h4C; #100;
A = 8'h55; B = 8'h4D; #100;
A = 8'h55; B = 8'h4E; #100;
A = 8'h55; B = 8'h4F; #100;
A = 8'h55; B = 8'h50; #100;
A = 8'h55; B = 8'h51; #100;
A = 8'h55; B = 8'h52; #100;
A = 8'h55; B = 8'h53; #100;
A = 8'h55; B = 8'h54; #100;
A = 8'h55; B = 8'h55; #100;
A = 8'h55; B = 8'h56; #100;
A = 8'h55; B = 8'h57; #100;
A = 8'h55; B = 8'h58; #100;
A = 8'h55; B = 8'h59; #100;
A = 8'h55; B = 8'h5A; #100;
A = 8'h55; B = 8'h5B; #100;
A = 8'h55; B = 8'h5C; #100;
A = 8'h55; B = 8'h5D; #100;
A = 8'h55; B = 8'h5E; #100;
A = 8'h55; B = 8'h5F; #100;
A = 8'h55; B = 8'h60; #100;
A = 8'h55; B = 8'h61; #100;
A = 8'h55; B = 8'h62; #100;
A = 8'h55; B = 8'h63; #100;
A = 8'h55; B = 8'h64; #100;
A = 8'h55; B = 8'h65; #100;
A = 8'h55; B = 8'h66; #100;
A = 8'h55; B = 8'h67; #100;
A = 8'h55; B = 8'h68; #100;
A = 8'h55; B = 8'h69; #100;
A = 8'h55; B = 8'h6A; #100;
A = 8'h55; B = 8'h6B; #100;
A = 8'h55; B = 8'h6C; #100;
A = 8'h55; B = 8'h6D; #100;
A = 8'h55; B = 8'h6E; #100;
A = 8'h55; B = 8'h6F; #100;
A = 8'h55; B = 8'h70; #100;
A = 8'h55; B = 8'h71; #100;
A = 8'h55; B = 8'h72; #100;
A = 8'h55; B = 8'h73; #100;
A = 8'h55; B = 8'h74; #100;
A = 8'h55; B = 8'h75; #100;
A = 8'h55; B = 8'h76; #100;
A = 8'h55; B = 8'h77; #100;
A = 8'h55; B = 8'h78; #100;
A = 8'h55; B = 8'h79; #100;
A = 8'h55; B = 8'h7A; #100;
A = 8'h55; B = 8'h7B; #100;
A = 8'h55; B = 8'h7C; #100;
A = 8'h55; B = 8'h7D; #100;
A = 8'h55; B = 8'h7E; #100;
A = 8'h55; B = 8'h7F; #100;
A = 8'h55; B = 8'h80; #100;
A = 8'h55; B = 8'h81; #100;
A = 8'h55; B = 8'h82; #100;
A = 8'h55; B = 8'h83; #100;
A = 8'h55; B = 8'h84; #100;
A = 8'h55; B = 8'h85; #100;
A = 8'h55; B = 8'h86; #100;
A = 8'h55; B = 8'h87; #100;
A = 8'h55; B = 8'h88; #100;
A = 8'h55; B = 8'h89; #100;
A = 8'h55; B = 8'h8A; #100;
A = 8'h55; B = 8'h8B; #100;
A = 8'h55; B = 8'h8C; #100;
A = 8'h55; B = 8'h8D; #100;
A = 8'h55; B = 8'h8E; #100;
A = 8'h55; B = 8'h8F; #100;
A = 8'h55; B = 8'h90; #100;
A = 8'h55; B = 8'h91; #100;
A = 8'h55; B = 8'h92; #100;
A = 8'h55; B = 8'h93; #100;
A = 8'h55; B = 8'h94; #100;
A = 8'h55; B = 8'h95; #100;
A = 8'h55; B = 8'h96; #100;
A = 8'h55; B = 8'h97; #100;
A = 8'h55; B = 8'h98; #100;
A = 8'h55; B = 8'h99; #100;
A = 8'h55; B = 8'h9A; #100;
A = 8'h55; B = 8'h9B; #100;
A = 8'h55; B = 8'h9C; #100;
A = 8'h55; B = 8'h9D; #100;
A = 8'h55; B = 8'h9E; #100;
A = 8'h55; B = 8'h9F; #100;
A = 8'h55; B = 8'hA0; #100;
A = 8'h55; B = 8'hA1; #100;
A = 8'h55; B = 8'hA2; #100;
A = 8'h55; B = 8'hA3; #100;
A = 8'h55; B = 8'hA4; #100;
A = 8'h55; B = 8'hA5; #100;
A = 8'h55; B = 8'hA6; #100;
A = 8'h55; B = 8'hA7; #100;
A = 8'h55; B = 8'hA8; #100;
A = 8'h55; B = 8'hA9; #100;
A = 8'h55; B = 8'hAA; #100;
A = 8'h55; B = 8'hAB; #100;
A = 8'h55; B = 8'hAC; #100;
A = 8'h55; B = 8'hAD; #100;
A = 8'h55; B = 8'hAE; #100;
A = 8'h55; B = 8'hAF; #100;
A = 8'h55; B = 8'hB0; #100;
A = 8'h55; B = 8'hB1; #100;
A = 8'h55; B = 8'hB2; #100;
A = 8'h55; B = 8'hB3; #100;
A = 8'h55; B = 8'hB4; #100;
A = 8'h55; B = 8'hB5; #100;
A = 8'h55; B = 8'hB6; #100;
A = 8'h55; B = 8'hB7; #100;
A = 8'h55; B = 8'hB8; #100;
A = 8'h55; B = 8'hB9; #100;
A = 8'h55; B = 8'hBA; #100;
A = 8'h55; B = 8'hBB; #100;
A = 8'h55; B = 8'hBC; #100;
A = 8'h55; B = 8'hBD; #100;
A = 8'h55; B = 8'hBE; #100;
A = 8'h55; B = 8'hBF; #100;
A = 8'h55; B = 8'hC0; #100;
A = 8'h55; B = 8'hC1; #100;
A = 8'h55; B = 8'hC2; #100;
A = 8'h55; B = 8'hC3; #100;
A = 8'h55; B = 8'hC4; #100;
A = 8'h55; B = 8'hC5; #100;
A = 8'h55; B = 8'hC6; #100;
A = 8'h55; B = 8'hC7; #100;
A = 8'h55; B = 8'hC8; #100;
A = 8'h55; B = 8'hC9; #100;
A = 8'h55; B = 8'hCA; #100;
A = 8'h55; B = 8'hCB; #100;
A = 8'h55; B = 8'hCC; #100;
A = 8'h55; B = 8'hCD; #100;
A = 8'h55; B = 8'hCE; #100;
A = 8'h55; B = 8'hCF; #100;
A = 8'h55; B = 8'hD0; #100;
A = 8'h55; B = 8'hD1; #100;
A = 8'h55; B = 8'hD2; #100;
A = 8'h55; B = 8'hD3; #100;
A = 8'h55; B = 8'hD4; #100;
A = 8'h55; B = 8'hD5; #100;
A = 8'h55; B = 8'hD6; #100;
A = 8'h55; B = 8'hD7; #100;
A = 8'h55; B = 8'hD8; #100;
A = 8'h55; B = 8'hD9; #100;
A = 8'h55; B = 8'hDA; #100;
A = 8'h55; B = 8'hDB; #100;
A = 8'h55; B = 8'hDC; #100;
A = 8'h55; B = 8'hDD; #100;
A = 8'h55; B = 8'hDE; #100;
A = 8'h55; B = 8'hDF; #100;
A = 8'h55; B = 8'hE0; #100;
A = 8'h55; B = 8'hE1; #100;
A = 8'h55; B = 8'hE2; #100;
A = 8'h55; B = 8'hE3; #100;
A = 8'h55; B = 8'hE4; #100;
A = 8'h55; B = 8'hE5; #100;
A = 8'h55; B = 8'hE6; #100;
A = 8'h55; B = 8'hE7; #100;
A = 8'h55; B = 8'hE8; #100;
A = 8'h55; B = 8'hE9; #100;
A = 8'h55; B = 8'hEA; #100;
A = 8'h55; B = 8'hEB; #100;
A = 8'h55; B = 8'hEC; #100;
A = 8'h55; B = 8'hED; #100;
A = 8'h55; B = 8'hEE; #100;
A = 8'h55; B = 8'hEF; #100;
A = 8'h55; B = 8'hF0; #100;
A = 8'h55; B = 8'hF1; #100;
A = 8'h55; B = 8'hF2; #100;
A = 8'h55; B = 8'hF3; #100;
A = 8'h55; B = 8'hF4; #100;
A = 8'h55; B = 8'hF5; #100;
A = 8'h55; B = 8'hF6; #100;
A = 8'h55; B = 8'hF7; #100;
A = 8'h55; B = 8'hF8; #100;
A = 8'h55; B = 8'hF9; #100;
A = 8'h55; B = 8'hFA; #100;
A = 8'h55; B = 8'hFB; #100;
A = 8'h55; B = 8'hFC; #100;
A = 8'h55; B = 8'hFD; #100;
A = 8'h55; B = 8'hFE; #100;
A = 8'h55; B = 8'hFF; #100;
A = 8'h56; B = 8'h0; #100;
A = 8'h56; B = 8'h1; #100;
A = 8'h56; B = 8'h2; #100;
A = 8'h56; B = 8'h3; #100;
A = 8'h56; B = 8'h4; #100;
A = 8'h56; B = 8'h5; #100;
A = 8'h56; B = 8'h6; #100;
A = 8'h56; B = 8'h7; #100;
A = 8'h56; B = 8'h8; #100;
A = 8'h56; B = 8'h9; #100;
A = 8'h56; B = 8'hA; #100;
A = 8'h56; B = 8'hB; #100;
A = 8'h56; B = 8'hC; #100;
A = 8'h56; B = 8'hD; #100;
A = 8'h56; B = 8'hE; #100;
A = 8'h56; B = 8'hF; #100;
A = 8'h56; B = 8'h10; #100;
A = 8'h56; B = 8'h11; #100;
A = 8'h56; B = 8'h12; #100;
A = 8'h56; B = 8'h13; #100;
A = 8'h56; B = 8'h14; #100;
A = 8'h56; B = 8'h15; #100;
A = 8'h56; B = 8'h16; #100;
A = 8'h56; B = 8'h17; #100;
A = 8'h56; B = 8'h18; #100;
A = 8'h56; B = 8'h19; #100;
A = 8'h56; B = 8'h1A; #100;
A = 8'h56; B = 8'h1B; #100;
A = 8'h56; B = 8'h1C; #100;
A = 8'h56; B = 8'h1D; #100;
A = 8'h56; B = 8'h1E; #100;
A = 8'h56; B = 8'h1F; #100;
A = 8'h56; B = 8'h20; #100;
A = 8'h56; B = 8'h21; #100;
A = 8'h56; B = 8'h22; #100;
A = 8'h56; B = 8'h23; #100;
A = 8'h56; B = 8'h24; #100;
A = 8'h56; B = 8'h25; #100;
A = 8'h56; B = 8'h26; #100;
A = 8'h56; B = 8'h27; #100;
A = 8'h56; B = 8'h28; #100;
A = 8'h56; B = 8'h29; #100;
A = 8'h56; B = 8'h2A; #100;
A = 8'h56; B = 8'h2B; #100;
A = 8'h56; B = 8'h2C; #100;
A = 8'h56; B = 8'h2D; #100;
A = 8'h56; B = 8'h2E; #100;
A = 8'h56; B = 8'h2F; #100;
A = 8'h56; B = 8'h30; #100;
A = 8'h56; B = 8'h31; #100;
A = 8'h56; B = 8'h32; #100;
A = 8'h56; B = 8'h33; #100;
A = 8'h56; B = 8'h34; #100;
A = 8'h56; B = 8'h35; #100;
A = 8'h56; B = 8'h36; #100;
A = 8'h56; B = 8'h37; #100;
A = 8'h56; B = 8'h38; #100;
A = 8'h56; B = 8'h39; #100;
A = 8'h56; B = 8'h3A; #100;
A = 8'h56; B = 8'h3B; #100;
A = 8'h56; B = 8'h3C; #100;
A = 8'h56; B = 8'h3D; #100;
A = 8'h56; B = 8'h3E; #100;
A = 8'h56; B = 8'h3F; #100;
A = 8'h56; B = 8'h40; #100;
A = 8'h56; B = 8'h41; #100;
A = 8'h56; B = 8'h42; #100;
A = 8'h56; B = 8'h43; #100;
A = 8'h56; B = 8'h44; #100;
A = 8'h56; B = 8'h45; #100;
A = 8'h56; B = 8'h46; #100;
A = 8'h56; B = 8'h47; #100;
A = 8'h56; B = 8'h48; #100;
A = 8'h56; B = 8'h49; #100;
A = 8'h56; B = 8'h4A; #100;
A = 8'h56; B = 8'h4B; #100;
A = 8'h56; B = 8'h4C; #100;
A = 8'h56; B = 8'h4D; #100;
A = 8'h56; B = 8'h4E; #100;
A = 8'h56; B = 8'h4F; #100;
A = 8'h56; B = 8'h50; #100;
A = 8'h56; B = 8'h51; #100;
A = 8'h56; B = 8'h52; #100;
A = 8'h56; B = 8'h53; #100;
A = 8'h56; B = 8'h54; #100;
A = 8'h56; B = 8'h55; #100;
A = 8'h56; B = 8'h56; #100;
A = 8'h56; B = 8'h57; #100;
A = 8'h56; B = 8'h58; #100;
A = 8'h56; B = 8'h59; #100;
A = 8'h56; B = 8'h5A; #100;
A = 8'h56; B = 8'h5B; #100;
A = 8'h56; B = 8'h5C; #100;
A = 8'h56; B = 8'h5D; #100;
A = 8'h56; B = 8'h5E; #100;
A = 8'h56; B = 8'h5F; #100;
A = 8'h56; B = 8'h60; #100;
A = 8'h56; B = 8'h61; #100;
A = 8'h56; B = 8'h62; #100;
A = 8'h56; B = 8'h63; #100;
A = 8'h56; B = 8'h64; #100;
A = 8'h56; B = 8'h65; #100;
A = 8'h56; B = 8'h66; #100;
A = 8'h56; B = 8'h67; #100;
A = 8'h56; B = 8'h68; #100;
A = 8'h56; B = 8'h69; #100;
A = 8'h56; B = 8'h6A; #100;
A = 8'h56; B = 8'h6B; #100;
A = 8'h56; B = 8'h6C; #100;
A = 8'h56; B = 8'h6D; #100;
A = 8'h56; B = 8'h6E; #100;
A = 8'h56; B = 8'h6F; #100;
A = 8'h56; B = 8'h70; #100;
A = 8'h56; B = 8'h71; #100;
A = 8'h56; B = 8'h72; #100;
A = 8'h56; B = 8'h73; #100;
A = 8'h56; B = 8'h74; #100;
A = 8'h56; B = 8'h75; #100;
A = 8'h56; B = 8'h76; #100;
A = 8'h56; B = 8'h77; #100;
A = 8'h56; B = 8'h78; #100;
A = 8'h56; B = 8'h79; #100;
A = 8'h56; B = 8'h7A; #100;
A = 8'h56; B = 8'h7B; #100;
A = 8'h56; B = 8'h7C; #100;
A = 8'h56; B = 8'h7D; #100;
A = 8'h56; B = 8'h7E; #100;
A = 8'h56; B = 8'h7F; #100;
A = 8'h56; B = 8'h80; #100;
A = 8'h56; B = 8'h81; #100;
A = 8'h56; B = 8'h82; #100;
A = 8'h56; B = 8'h83; #100;
A = 8'h56; B = 8'h84; #100;
A = 8'h56; B = 8'h85; #100;
A = 8'h56; B = 8'h86; #100;
A = 8'h56; B = 8'h87; #100;
A = 8'h56; B = 8'h88; #100;
A = 8'h56; B = 8'h89; #100;
A = 8'h56; B = 8'h8A; #100;
A = 8'h56; B = 8'h8B; #100;
A = 8'h56; B = 8'h8C; #100;
A = 8'h56; B = 8'h8D; #100;
A = 8'h56; B = 8'h8E; #100;
A = 8'h56; B = 8'h8F; #100;
A = 8'h56; B = 8'h90; #100;
A = 8'h56; B = 8'h91; #100;
A = 8'h56; B = 8'h92; #100;
A = 8'h56; B = 8'h93; #100;
A = 8'h56; B = 8'h94; #100;
A = 8'h56; B = 8'h95; #100;
A = 8'h56; B = 8'h96; #100;
A = 8'h56; B = 8'h97; #100;
A = 8'h56; B = 8'h98; #100;
A = 8'h56; B = 8'h99; #100;
A = 8'h56; B = 8'h9A; #100;
A = 8'h56; B = 8'h9B; #100;
A = 8'h56; B = 8'h9C; #100;
A = 8'h56; B = 8'h9D; #100;
A = 8'h56; B = 8'h9E; #100;
A = 8'h56; B = 8'h9F; #100;
A = 8'h56; B = 8'hA0; #100;
A = 8'h56; B = 8'hA1; #100;
A = 8'h56; B = 8'hA2; #100;
A = 8'h56; B = 8'hA3; #100;
A = 8'h56; B = 8'hA4; #100;
A = 8'h56; B = 8'hA5; #100;
A = 8'h56; B = 8'hA6; #100;
A = 8'h56; B = 8'hA7; #100;
A = 8'h56; B = 8'hA8; #100;
A = 8'h56; B = 8'hA9; #100;
A = 8'h56; B = 8'hAA; #100;
A = 8'h56; B = 8'hAB; #100;
A = 8'h56; B = 8'hAC; #100;
A = 8'h56; B = 8'hAD; #100;
A = 8'h56; B = 8'hAE; #100;
A = 8'h56; B = 8'hAF; #100;
A = 8'h56; B = 8'hB0; #100;
A = 8'h56; B = 8'hB1; #100;
A = 8'h56; B = 8'hB2; #100;
A = 8'h56; B = 8'hB3; #100;
A = 8'h56; B = 8'hB4; #100;
A = 8'h56; B = 8'hB5; #100;
A = 8'h56; B = 8'hB6; #100;
A = 8'h56; B = 8'hB7; #100;
A = 8'h56; B = 8'hB8; #100;
A = 8'h56; B = 8'hB9; #100;
A = 8'h56; B = 8'hBA; #100;
A = 8'h56; B = 8'hBB; #100;
A = 8'h56; B = 8'hBC; #100;
A = 8'h56; B = 8'hBD; #100;
A = 8'h56; B = 8'hBE; #100;
A = 8'h56; B = 8'hBF; #100;
A = 8'h56; B = 8'hC0; #100;
A = 8'h56; B = 8'hC1; #100;
A = 8'h56; B = 8'hC2; #100;
A = 8'h56; B = 8'hC3; #100;
A = 8'h56; B = 8'hC4; #100;
A = 8'h56; B = 8'hC5; #100;
A = 8'h56; B = 8'hC6; #100;
A = 8'h56; B = 8'hC7; #100;
A = 8'h56; B = 8'hC8; #100;
A = 8'h56; B = 8'hC9; #100;
A = 8'h56; B = 8'hCA; #100;
A = 8'h56; B = 8'hCB; #100;
A = 8'h56; B = 8'hCC; #100;
A = 8'h56; B = 8'hCD; #100;
A = 8'h56; B = 8'hCE; #100;
A = 8'h56; B = 8'hCF; #100;
A = 8'h56; B = 8'hD0; #100;
A = 8'h56; B = 8'hD1; #100;
A = 8'h56; B = 8'hD2; #100;
A = 8'h56; B = 8'hD3; #100;
A = 8'h56; B = 8'hD4; #100;
A = 8'h56; B = 8'hD5; #100;
A = 8'h56; B = 8'hD6; #100;
A = 8'h56; B = 8'hD7; #100;
A = 8'h56; B = 8'hD8; #100;
A = 8'h56; B = 8'hD9; #100;
A = 8'h56; B = 8'hDA; #100;
A = 8'h56; B = 8'hDB; #100;
A = 8'h56; B = 8'hDC; #100;
A = 8'h56; B = 8'hDD; #100;
A = 8'h56; B = 8'hDE; #100;
A = 8'h56; B = 8'hDF; #100;
A = 8'h56; B = 8'hE0; #100;
A = 8'h56; B = 8'hE1; #100;
A = 8'h56; B = 8'hE2; #100;
A = 8'h56; B = 8'hE3; #100;
A = 8'h56; B = 8'hE4; #100;
A = 8'h56; B = 8'hE5; #100;
A = 8'h56; B = 8'hE6; #100;
A = 8'h56; B = 8'hE7; #100;
A = 8'h56; B = 8'hE8; #100;
A = 8'h56; B = 8'hE9; #100;
A = 8'h56; B = 8'hEA; #100;
A = 8'h56; B = 8'hEB; #100;
A = 8'h56; B = 8'hEC; #100;
A = 8'h56; B = 8'hED; #100;
A = 8'h56; B = 8'hEE; #100;
A = 8'h56; B = 8'hEF; #100;
A = 8'h56; B = 8'hF0; #100;
A = 8'h56; B = 8'hF1; #100;
A = 8'h56; B = 8'hF2; #100;
A = 8'h56; B = 8'hF3; #100;
A = 8'h56; B = 8'hF4; #100;
A = 8'h56; B = 8'hF5; #100;
A = 8'h56; B = 8'hF6; #100;
A = 8'h56; B = 8'hF7; #100;
A = 8'h56; B = 8'hF8; #100;
A = 8'h56; B = 8'hF9; #100;
A = 8'h56; B = 8'hFA; #100;
A = 8'h56; B = 8'hFB; #100;
A = 8'h56; B = 8'hFC; #100;
A = 8'h56; B = 8'hFD; #100;
A = 8'h56; B = 8'hFE; #100;
A = 8'h56; B = 8'hFF; #100;
A = 8'h57; B = 8'h0; #100;
A = 8'h57; B = 8'h1; #100;
A = 8'h57; B = 8'h2; #100;
A = 8'h57; B = 8'h3; #100;
A = 8'h57; B = 8'h4; #100;
A = 8'h57; B = 8'h5; #100;
A = 8'h57; B = 8'h6; #100;
A = 8'h57; B = 8'h7; #100;
A = 8'h57; B = 8'h8; #100;
A = 8'h57; B = 8'h9; #100;
A = 8'h57; B = 8'hA; #100;
A = 8'h57; B = 8'hB; #100;
A = 8'h57; B = 8'hC; #100;
A = 8'h57; B = 8'hD; #100;
A = 8'h57; B = 8'hE; #100;
A = 8'h57; B = 8'hF; #100;
A = 8'h57; B = 8'h10; #100;
A = 8'h57; B = 8'h11; #100;
A = 8'h57; B = 8'h12; #100;
A = 8'h57; B = 8'h13; #100;
A = 8'h57; B = 8'h14; #100;
A = 8'h57; B = 8'h15; #100;
A = 8'h57; B = 8'h16; #100;
A = 8'h57; B = 8'h17; #100;
A = 8'h57; B = 8'h18; #100;
A = 8'h57; B = 8'h19; #100;
A = 8'h57; B = 8'h1A; #100;
A = 8'h57; B = 8'h1B; #100;
A = 8'h57; B = 8'h1C; #100;
A = 8'h57; B = 8'h1D; #100;
A = 8'h57; B = 8'h1E; #100;
A = 8'h57; B = 8'h1F; #100;
A = 8'h57; B = 8'h20; #100;
A = 8'h57; B = 8'h21; #100;
A = 8'h57; B = 8'h22; #100;
A = 8'h57; B = 8'h23; #100;
A = 8'h57; B = 8'h24; #100;
A = 8'h57; B = 8'h25; #100;
A = 8'h57; B = 8'h26; #100;
A = 8'h57; B = 8'h27; #100;
A = 8'h57; B = 8'h28; #100;
A = 8'h57; B = 8'h29; #100;
A = 8'h57; B = 8'h2A; #100;
A = 8'h57; B = 8'h2B; #100;
A = 8'h57; B = 8'h2C; #100;
A = 8'h57; B = 8'h2D; #100;
A = 8'h57; B = 8'h2E; #100;
A = 8'h57; B = 8'h2F; #100;
A = 8'h57; B = 8'h30; #100;
A = 8'h57; B = 8'h31; #100;
A = 8'h57; B = 8'h32; #100;
A = 8'h57; B = 8'h33; #100;
A = 8'h57; B = 8'h34; #100;
A = 8'h57; B = 8'h35; #100;
A = 8'h57; B = 8'h36; #100;
A = 8'h57; B = 8'h37; #100;
A = 8'h57; B = 8'h38; #100;
A = 8'h57; B = 8'h39; #100;
A = 8'h57; B = 8'h3A; #100;
A = 8'h57; B = 8'h3B; #100;
A = 8'h57; B = 8'h3C; #100;
A = 8'h57; B = 8'h3D; #100;
A = 8'h57; B = 8'h3E; #100;
A = 8'h57; B = 8'h3F; #100;
A = 8'h57; B = 8'h40; #100;
A = 8'h57; B = 8'h41; #100;
A = 8'h57; B = 8'h42; #100;
A = 8'h57; B = 8'h43; #100;
A = 8'h57; B = 8'h44; #100;
A = 8'h57; B = 8'h45; #100;
A = 8'h57; B = 8'h46; #100;
A = 8'h57; B = 8'h47; #100;
A = 8'h57; B = 8'h48; #100;
A = 8'h57; B = 8'h49; #100;
A = 8'h57; B = 8'h4A; #100;
A = 8'h57; B = 8'h4B; #100;
A = 8'h57; B = 8'h4C; #100;
A = 8'h57; B = 8'h4D; #100;
A = 8'h57; B = 8'h4E; #100;
A = 8'h57; B = 8'h4F; #100;
A = 8'h57; B = 8'h50; #100;
A = 8'h57; B = 8'h51; #100;
A = 8'h57; B = 8'h52; #100;
A = 8'h57; B = 8'h53; #100;
A = 8'h57; B = 8'h54; #100;
A = 8'h57; B = 8'h55; #100;
A = 8'h57; B = 8'h56; #100;
A = 8'h57; B = 8'h57; #100;
A = 8'h57; B = 8'h58; #100;
A = 8'h57; B = 8'h59; #100;
A = 8'h57; B = 8'h5A; #100;
A = 8'h57; B = 8'h5B; #100;
A = 8'h57; B = 8'h5C; #100;
A = 8'h57; B = 8'h5D; #100;
A = 8'h57; B = 8'h5E; #100;
A = 8'h57; B = 8'h5F; #100;
A = 8'h57; B = 8'h60; #100;
A = 8'h57; B = 8'h61; #100;
A = 8'h57; B = 8'h62; #100;
A = 8'h57; B = 8'h63; #100;
A = 8'h57; B = 8'h64; #100;
A = 8'h57; B = 8'h65; #100;
A = 8'h57; B = 8'h66; #100;
A = 8'h57; B = 8'h67; #100;
A = 8'h57; B = 8'h68; #100;
A = 8'h57; B = 8'h69; #100;
A = 8'h57; B = 8'h6A; #100;
A = 8'h57; B = 8'h6B; #100;
A = 8'h57; B = 8'h6C; #100;
A = 8'h57; B = 8'h6D; #100;
A = 8'h57; B = 8'h6E; #100;
A = 8'h57; B = 8'h6F; #100;
A = 8'h57; B = 8'h70; #100;
A = 8'h57; B = 8'h71; #100;
A = 8'h57; B = 8'h72; #100;
A = 8'h57; B = 8'h73; #100;
A = 8'h57; B = 8'h74; #100;
A = 8'h57; B = 8'h75; #100;
A = 8'h57; B = 8'h76; #100;
A = 8'h57; B = 8'h77; #100;
A = 8'h57; B = 8'h78; #100;
A = 8'h57; B = 8'h79; #100;
A = 8'h57; B = 8'h7A; #100;
A = 8'h57; B = 8'h7B; #100;
A = 8'h57; B = 8'h7C; #100;
A = 8'h57; B = 8'h7D; #100;
A = 8'h57; B = 8'h7E; #100;
A = 8'h57; B = 8'h7F; #100;
A = 8'h57; B = 8'h80; #100;
A = 8'h57; B = 8'h81; #100;
A = 8'h57; B = 8'h82; #100;
A = 8'h57; B = 8'h83; #100;
A = 8'h57; B = 8'h84; #100;
A = 8'h57; B = 8'h85; #100;
A = 8'h57; B = 8'h86; #100;
A = 8'h57; B = 8'h87; #100;
A = 8'h57; B = 8'h88; #100;
A = 8'h57; B = 8'h89; #100;
A = 8'h57; B = 8'h8A; #100;
A = 8'h57; B = 8'h8B; #100;
A = 8'h57; B = 8'h8C; #100;
A = 8'h57; B = 8'h8D; #100;
A = 8'h57; B = 8'h8E; #100;
A = 8'h57; B = 8'h8F; #100;
A = 8'h57; B = 8'h90; #100;
A = 8'h57; B = 8'h91; #100;
A = 8'h57; B = 8'h92; #100;
A = 8'h57; B = 8'h93; #100;
A = 8'h57; B = 8'h94; #100;
A = 8'h57; B = 8'h95; #100;
A = 8'h57; B = 8'h96; #100;
A = 8'h57; B = 8'h97; #100;
A = 8'h57; B = 8'h98; #100;
A = 8'h57; B = 8'h99; #100;
A = 8'h57; B = 8'h9A; #100;
A = 8'h57; B = 8'h9B; #100;
A = 8'h57; B = 8'h9C; #100;
A = 8'h57; B = 8'h9D; #100;
A = 8'h57; B = 8'h9E; #100;
A = 8'h57; B = 8'h9F; #100;
A = 8'h57; B = 8'hA0; #100;
A = 8'h57; B = 8'hA1; #100;
A = 8'h57; B = 8'hA2; #100;
A = 8'h57; B = 8'hA3; #100;
A = 8'h57; B = 8'hA4; #100;
A = 8'h57; B = 8'hA5; #100;
A = 8'h57; B = 8'hA6; #100;
A = 8'h57; B = 8'hA7; #100;
A = 8'h57; B = 8'hA8; #100;
A = 8'h57; B = 8'hA9; #100;
A = 8'h57; B = 8'hAA; #100;
A = 8'h57; B = 8'hAB; #100;
A = 8'h57; B = 8'hAC; #100;
A = 8'h57; B = 8'hAD; #100;
A = 8'h57; B = 8'hAE; #100;
A = 8'h57; B = 8'hAF; #100;
A = 8'h57; B = 8'hB0; #100;
A = 8'h57; B = 8'hB1; #100;
A = 8'h57; B = 8'hB2; #100;
A = 8'h57; B = 8'hB3; #100;
A = 8'h57; B = 8'hB4; #100;
A = 8'h57; B = 8'hB5; #100;
A = 8'h57; B = 8'hB6; #100;
A = 8'h57; B = 8'hB7; #100;
A = 8'h57; B = 8'hB8; #100;
A = 8'h57; B = 8'hB9; #100;
A = 8'h57; B = 8'hBA; #100;
A = 8'h57; B = 8'hBB; #100;
A = 8'h57; B = 8'hBC; #100;
A = 8'h57; B = 8'hBD; #100;
A = 8'h57; B = 8'hBE; #100;
A = 8'h57; B = 8'hBF; #100;
A = 8'h57; B = 8'hC0; #100;
A = 8'h57; B = 8'hC1; #100;
A = 8'h57; B = 8'hC2; #100;
A = 8'h57; B = 8'hC3; #100;
A = 8'h57; B = 8'hC4; #100;
A = 8'h57; B = 8'hC5; #100;
A = 8'h57; B = 8'hC6; #100;
A = 8'h57; B = 8'hC7; #100;
A = 8'h57; B = 8'hC8; #100;
A = 8'h57; B = 8'hC9; #100;
A = 8'h57; B = 8'hCA; #100;
A = 8'h57; B = 8'hCB; #100;
A = 8'h57; B = 8'hCC; #100;
A = 8'h57; B = 8'hCD; #100;
A = 8'h57; B = 8'hCE; #100;
A = 8'h57; B = 8'hCF; #100;
A = 8'h57; B = 8'hD0; #100;
A = 8'h57; B = 8'hD1; #100;
A = 8'h57; B = 8'hD2; #100;
A = 8'h57; B = 8'hD3; #100;
A = 8'h57; B = 8'hD4; #100;
A = 8'h57; B = 8'hD5; #100;
A = 8'h57; B = 8'hD6; #100;
A = 8'h57; B = 8'hD7; #100;
A = 8'h57; B = 8'hD8; #100;
A = 8'h57; B = 8'hD9; #100;
A = 8'h57; B = 8'hDA; #100;
A = 8'h57; B = 8'hDB; #100;
A = 8'h57; B = 8'hDC; #100;
A = 8'h57; B = 8'hDD; #100;
A = 8'h57; B = 8'hDE; #100;
A = 8'h57; B = 8'hDF; #100;
A = 8'h57; B = 8'hE0; #100;
A = 8'h57; B = 8'hE1; #100;
A = 8'h57; B = 8'hE2; #100;
A = 8'h57; B = 8'hE3; #100;
A = 8'h57; B = 8'hE4; #100;
A = 8'h57; B = 8'hE5; #100;
A = 8'h57; B = 8'hE6; #100;
A = 8'h57; B = 8'hE7; #100;
A = 8'h57; B = 8'hE8; #100;
A = 8'h57; B = 8'hE9; #100;
A = 8'h57; B = 8'hEA; #100;
A = 8'h57; B = 8'hEB; #100;
A = 8'h57; B = 8'hEC; #100;
A = 8'h57; B = 8'hED; #100;
A = 8'h57; B = 8'hEE; #100;
A = 8'h57; B = 8'hEF; #100;
A = 8'h57; B = 8'hF0; #100;
A = 8'h57; B = 8'hF1; #100;
A = 8'h57; B = 8'hF2; #100;
A = 8'h57; B = 8'hF3; #100;
A = 8'h57; B = 8'hF4; #100;
A = 8'h57; B = 8'hF5; #100;
A = 8'h57; B = 8'hF6; #100;
A = 8'h57; B = 8'hF7; #100;
A = 8'h57; B = 8'hF8; #100;
A = 8'h57; B = 8'hF9; #100;
A = 8'h57; B = 8'hFA; #100;
A = 8'h57; B = 8'hFB; #100;
A = 8'h57; B = 8'hFC; #100;
A = 8'h57; B = 8'hFD; #100;
A = 8'h57; B = 8'hFE; #100;
A = 8'h57; B = 8'hFF; #100;
A = 8'h58; B = 8'h0; #100;
A = 8'h58; B = 8'h1; #100;
A = 8'h58; B = 8'h2; #100;
A = 8'h58; B = 8'h3; #100;
A = 8'h58; B = 8'h4; #100;
A = 8'h58; B = 8'h5; #100;
A = 8'h58; B = 8'h6; #100;
A = 8'h58; B = 8'h7; #100;
A = 8'h58; B = 8'h8; #100;
A = 8'h58; B = 8'h9; #100;
A = 8'h58; B = 8'hA; #100;
A = 8'h58; B = 8'hB; #100;
A = 8'h58; B = 8'hC; #100;
A = 8'h58; B = 8'hD; #100;
A = 8'h58; B = 8'hE; #100;
A = 8'h58; B = 8'hF; #100;
A = 8'h58; B = 8'h10; #100;
A = 8'h58; B = 8'h11; #100;
A = 8'h58; B = 8'h12; #100;
A = 8'h58; B = 8'h13; #100;
A = 8'h58; B = 8'h14; #100;
A = 8'h58; B = 8'h15; #100;
A = 8'h58; B = 8'h16; #100;
A = 8'h58; B = 8'h17; #100;
A = 8'h58; B = 8'h18; #100;
A = 8'h58; B = 8'h19; #100;
A = 8'h58; B = 8'h1A; #100;
A = 8'h58; B = 8'h1B; #100;
A = 8'h58; B = 8'h1C; #100;
A = 8'h58; B = 8'h1D; #100;
A = 8'h58; B = 8'h1E; #100;
A = 8'h58; B = 8'h1F; #100;
A = 8'h58; B = 8'h20; #100;
A = 8'h58; B = 8'h21; #100;
A = 8'h58; B = 8'h22; #100;
A = 8'h58; B = 8'h23; #100;
A = 8'h58; B = 8'h24; #100;
A = 8'h58; B = 8'h25; #100;
A = 8'h58; B = 8'h26; #100;
A = 8'h58; B = 8'h27; #100;
A = 8'h58; B = 8'h28; #100;
A = 8'h58; B = 8'h29; #100;
A = 8'h58; B = 8'h2A; #100;
A = 8'h58; B = 8'h2B; #100;
A = 8'h58; B = 8'h2C; #100;
A = 8'h58; B = 8'h2D; #100;
A = 8'h58; B = 8'h2E; #100;
A = 8'h58; B = 8'h2F; #100;
A = 8'h58; B = 8'h30; #100;
A = 8'h58; B = 8'h31; #100;
A = 8'h58; B = 8'h32; #100;
A = 8'h58; B = 8'h33; #100;
A = 8'h58; B = 8'h34; #100;
A = 8'h58; B = 8'h35; #100;
A = 8'h58; B = 8'h36; #100;
A = 8'h58; B = 8'h37; #100;
A = 8'h58; B = 8'h38; #100;
A = 8'h58; B = 8'h39; #100;
A = 8'h58; B = 8'h3A; #100;
A = 8'h58; B = 8'h3B; #100;
A = 8'h58; B = 8'h3C; #100;
A = 8'h58; B = 8'h3D; #100;
A = 8'h58; B = 8'h3E; #100;
A = 8'h58; B = 8'h3F; #100;
A = 8'h58; B = 8'h40; #100;
A = 8'h58; B = 8'h41; #100;
A = 8'h58; B = 8'h42; #100;
A = 8'h58; B = 8'h43; #100;
A = 8'h58; B = 8'h44; #100;
A = 8'h58; B = 8'h45; #100;
A = 8'h58; B = 8'h46; #100;
A = 8'h58; B = 8'h47; #100;
A = 8'h58; B = 8'h48; #100;
A = 8'h58; B = 8'h49; #100;
A = 8'h58; B = 8'h4A; #100;
A = 8'h58; B = 8'h4B; #100;
A = 8'h58; B = 8'h4C; #100;
A = 8'h58; B = 8'h4D; #100;
A = 8'h58; B = 8'h4E; #100;
A = 8'h58; B = 8'h4F; #100;
A = 8'h58; B = 8'h50; #100;
A = 8'h58; B = 8'h51; #100;
A = 8'h58; B = 8'h52; #100;
A = 8'h58; B = 8'h53; #100;
A = 8'h58; B = 8'h54; #100;
A = 8'h58; B = 8'h55; #100;
A = 8'h58; B = 8'h56; #100;
A = 8'h58; B = 8'h57; #100;
A = 8'h58; B = 8'h58; #100;
A = 8'h58; B = 8'h59; #100;
A = 8'h58; B = 8'h5A; #100;
A = 8'h58; B = 8'h5B; #100;
A = 8'h58; B = 8'h5C; #100;
A = 8'h58; B = 8'h5D; #100;
A = 8'h58; B = 8'h5E; #100;
A = 8'h58; B = 8'h5F; #100;
A = 8'h58; B = 8'h60; #100;
A = 8'h58; B = 8'h61; #100;
A = 8'h58; B = 8'h62; #100;
A = 8'h58; B = 8'h63; #100;
A = 8'h58; B = 8'h64; #100;
A = 8'h58; B = 8'h65; #100;
A = 8'h58; B = 8'h66; #100;
A = 8'h58; B = 8'h67; #100;
A = 8'h58; B = 8'h68; #100;
A = 8'h58; B = 8'h69; #100;
A = 8'h58; B = 8'h6A; #100;
A = 8'h58; B = 8'h6B; #100;
A = 8'h58; B = 8'h6C; #100;
A = 8'h58; B = 8'h6D; #100;
A = 8'h58; B = 8'h6E; #100;
A = 8'h58; B = 8'h6F; #100;
A = 8'h58; B = 8'h70; #100;
A = 8'h58; B = 8'h71; #100;
A = 8'h58; B = 8'h72; #100;
A = 8'h58; B = 8'h73; #100;
A = 8'h58; B = 8'h74; #100;
A = 8'h58; B = 8'h75; #100;
A = 8'h58; B = 8'h76; #100;
A = 8'h58; B = 8'h77; #100;
A = 8'h58; B = 8'h78; #100;
A = 8'h58; B = 8'h79; #100;
A = 8'h58; B = 8'h7A; #100;
A = 8'h58; B = 8'h7B; #100;
A = 8'h58; B = 8'h7C; #100;
A = 8'h58; B = 8'h7D; #100;
A = 8'h58; B = 8'h7E; #100;
A = 8'h58; B = 8'h7F; #100;
A = 8'h58; B = 8'h80; #100;
A = 8'h58; B = 8'h81; #100;
A = 8'h58; B = 8'h82; #100;
A = 8'h58; B = 8'h83; #100;
A = 8'h58; B = 8'h84; #100;
A = 8'h58; B = 8'h85; #100;
A = 8'h58; B = 8'h86; #100;
A = 8'h58; B = 8'h87; #100;
A = 8'h58; B = 8'h88; #100;
A = 8'h58; B = 8'h89; #100;
A = 8'h58; B = 8'h8A; #100;
A = 8'h58; B = 8'h8B; #100;
A = 8'h58; B = 8'h8C; #100;
A = 8'h58; B = 8'h8D; #100;
A = 8'h58; B = 8'h8E; #100;
A = 8'h58; B = 8'h8F; #100;
A = 8'h58; B = 8'h90; #100;
A = 8'h58; B = 8'h91; #100;
A = 8'h58; B = 8'h92; #100;
A = 8'h58; B = 8'h93; #100;
A = 8'h58; B = 8'h94; #100;
A = 8'h58; B = 8'h95; #100;
A = 8'h58; B = 8'h96; #100;
A = 8'h58; B = 8'h97; #100;
A = 8'h58; B = 8'h98; #100;
A = 8'h58; B = 8'h99; #100;
A = 8'h58; B = 8'h9A; #100;
A = 8'h58; B = 8'h9B; #100;
A = 8'h58; B = 8'h9C; #100;
A = 8'h58; B = 8'h9D; #100;
A = 8'h58; B = 8'h9E; #100;
A = 8'h58; B = 8'h9F; #100;
A = 8'h58; B = 8'hA0; #100;
A = 8'h58; B = 8'hA1; #100;
A = 8'h58; B = 8'hA2; #100;
A = 8'h58; B = 8'hA3; #100;
A = 8'h58; B = 8'hA4; #100;
A = 8'h58; B = 8'hA5; #100;
A = 8'h58; B = 8'hA6; #100;
A = 8'h58; B = 8'hA7; #100;
A = 8'h58; B = 8'hA8; #100;
A = 8'h58; B = 8'hA9; #100;
A = 8'h58; B = 8'hAA; #100;
A = 8'h58; B = 8'hAB; #100;
A = 8'h58; B = 8'hAC; #100;
A = 8'h58; B = 8'hAD; #100;
A = 8'h58; B = 8'hAE; #100;
A = 8'h58; B = 8'hAF; #100;
A = 8'h58; B = 8'hB0; #100;
A = 8'h58; B = 8'hB1; #100;
A = 8'h58; B = 8'hB2; #100;
A = 8'h58; B = 8'hB3; #100;
A = 8'h58; B = 8'hB4; #100;
A = 8'h58; B = 8'hB5; #100;
A = 8'h58; B = 8'hB6; #100;
A = 8'h58; B = 8'hB7; #100;
A = 8'h58; B = 8'hB8; #100;
A = 8'h58; B = 8'hB9; #100;
A = 8'h58; B = 8'hBA; #100;
A = 8'h58; B = 8'hBB; #100;
A = 8'h58; B = 8'hBC; #100;
A = 8'h58; B = 8'hBD; #100;
A = 8'h58; B = 8'hBE; #100;
A = 8'h58; B = 8'hBF; #100;
A = 8'h58; B = 8'hC0; #100;
A = 8'h58; B = 8'hC1; #100;
A = 8'h58; B = 8'hC2; #100;
A = 8'h58; B = 8'hC3; #100;
A = 8'h58; B = 8'hC4; #100;
A = 8'h58; B = 8'hC5; #100;
A = 8'h58; B = 8'hC6; #100;
A = 8'h58; B = 8'hC7; #100;
A = 8'h58; B = 8'hC8; #100;
A = 8'h58; B = 8'hC9; #100;
A = 8'h58; B = 8'hCA; #100;
A = 8'h58; B = 8'hCB; #100;
A = 8'h58; B = 8'hCC; #100;
A = 8'h58; B = 8'hCD; #100;
A = 8'h58; B = 8'hCE; #100;
A = 8'h58; B = 8'hCF; #100;
A = 8'h58; B = 8'hD0; #100;
A = 8'h58; B = 8'hD1; #100;
A = 8'h58; B = 8'hD2; #100;
A = 8'h58; B = 8'hD3; #100;
A = 8'h58; B = 8'hD4; #100;
A = 8'h58; B = 8'hD5; #100;
A = 8'h58; B = 8'hD6; #100;
A = 8'h58; B = 8'hD7; #100;
A = 8'h58; B = 8'hD8; #100;
A = 8'h58; B = 8'hD9; #100;
A = 8'h58; B = 8'hDA; #100;
A = 8'h58; B = 8'hDB; #100;
A = 8'h58; B = 8'hDC; #100;
A = 8'h58; B = 8'hDD; #100;
A = 8'h58; B = 8'hDE; #100;
A = 8'h58; B = 8'hDF; #100;
A = 8'h58; B = 8'hE0; #100;
A = 8'h58; B = 8'hE1; #100;
A = 8'h58; B = 8'hE2; #100;
A = 8'h58; B = 8'hE3; #100;
A = 8'h58; B = 8'hE4; #100;
A = 8'h58; B = 8'hE5; #100;
A = 8'h58; B = 8'hE6; #100;
A = 8'h58; B = 8'hE7; #100;
A = 8'h58; B = 8'hE8; #100;
A = 8'h58; B = 8'hE9; #100;
A = 8'h58; B = 8'hEA; #100;
A = 8'h58; B = 8'hEB; #100;
A = 8'h58; B = 8'hEC; #100;
A = 8'h58; B = 8'hED; #100;
A = 8'h58; B = 8'hEE; #100;
A = 8'h58; B = 8'hEF; #100;
A = 8'h58; B = 8'hF0; #100;
A = 8'h58; B = 8'hF1; #100;
A = 8'h58; B = 8'hF2; #100;
A = 8'h58; B = 8'hF3; #100;
A = 8'h58; B = 8'hF4; #100;
A = 8'h58; B = 8'hF5; #100;
A = 8'h58; B = 8'hF6; #100;
A = 8'h58; B = 8'hF7; #100;
A = 8'h58; B = 8'hF8; #100;
A = 8'h58; B = 8'hF9; #100;
A = 8'h58; B = 8'hFA; #100;
A = 8'h58; B = 8'hFB; #100;
A = 8'h58; B = 8'hFC; #100;
A = 8'h58; B = 8'hFD; #100;
A = 8'h58; B = 8'hFE; #100;
A = 8'h58; B = 8'hFF; #100;
A = 8'h59; B = 8'h0; #100;
A = 8'h59; B = 8'h1; #100;
A = 8'h59; B = 8'h2; #100;
A = 8'h59; B = 8'h3; #100;
A = 8'h59; B = 8'h4; #100;
A = 8'h59; B = 8'h5; #100;
A = 8'h59; B = 8'h6; #100;
A = 8'h59; B = 8'h7; #100;
A = 8'h59; B = 8'h8; #100;
A = 8'h59; B = 8'h9; #100;
A = 8'h59; B = 8'hA; #100;
A = 8'h59; B = 8'hB; #100;
A = 8'h59; B = 8'hC; #100;
A = 8'h59; B = 8'hD; #100;
A = 8'h59; B = 8'hE; #100;
A = 8'h59; B = 8'hF; #100;
A = 8'h59; B = 8'h10; #100;
A = 8'h59; B = 8'h11; #100;
A = 8'h59; B = 8'h12; #100;
A = 8'h59; B = 8'h13; #100;
A = 8'h59; B = 8'h14; #100;
A = 8'h59; B = 8'h15; #100;
A = 8'h59; B = 8'h16; #100;
A = 8'h59; B = 8'h17; #100;
A = 8'h59; B = 8'h18; #100;
A = 8'h59; B = 8'h19; #100;
A = 8'h59; B = 8'h1A; #100;
A = 8'h59; B = 8'h1B; #100;
A = 8'h59; B = 8'h1C; #100;
A = 8'h59; B = 8'h1D; #100;
A = 8'h59; B = 8'h1E; #100;
A = 8'h59; B = 8'h1F; #100;
A = 8'h59; B = 8'h20; #100;
A = 8'h59; B = 8'h21; #100;
A = 8'h59; B = 8'h22; #100;
A = 8'h59; B = 8'h23; #100;
A = 8'h59; B = 8'h24; #100;
A = 8'h59; B = 8'h25; #100;
A = 8'h59; B = 8'h26; #100;
A = 8'h59; B = 8'h27; #100;
A = 8'h59; B = 8'h28; #100;
A = 8'h59; B = 8'h29; #100;
A = 8'h59; B = 8'h2A; #100;
A = 8'h59; B = 8'h2B; #100;
A = 8'h59; B = 8'h2C; #100;
A = 8'h59; B = 8'h2D; #100;
A = 8'h59; B = 8'h2E; #100;
A = 8'h59; B = 8'h2F; #100;
A = 8'h59; B = 8'h30; #100;
A = 8'h59; B = 8'h31; #100;
A = 8'h59; B = 8'h32; #100;
A = 8'h59; B = 8'h33; #100;
A = 8'h59; B = 8'h34; #100;
A = 8'h59; B = 8'h35; #100;
A = 8'h59; B = 8'h36; #100;
A = 8'h59; B = 8'h37; #100;
A = 8'h59; B = 8'h38; #100;
A = 8'h59; B = 8'h39; #100;
A = 8'h59; B = 8'h3A; #100;
A = 8'h59; B = 8'h3B; #100;
A = 8'h59; B = 8'h3C; #100;
A = 8'h59; B = 8'h3D; #100;
A = 8'h59; B = 8'h3E; #100;
A = 8'h59; B = 8'h3F; #100;
A = 8'h59; B = 8'h40; #100;
A = 8'h59; B = 8'h41; #100;
A = 8'h59; B = 8'h42; #100;
A = 8'h59; B = 8'h43; #100;
A = 8'h59; B = 8'h44; #100;
A = 8'h59; B = 8'h45; #100;
A = 8'h59; B = 8'h46; #100;
A = 8'h59; B = 8'h47; #100;
A = 8'h59; B = 8'h48; #100;
A = 8'h59; B = 8'h49; #100;
A = 8'h59; B = 8'h4A; #100;
A = 8'h59; B = 8'h4B; #100;
A = 8'h59; B = 8'h4C; #100;
A = 8'h59; B = 8'h4D; #100;
A = 8'h59; B = 8'h4E; #100;
A = 8'h59; B = 8'h4F; #100;
A = 8'h59; B = 8'h50; #100;
A = 8'h59; B = 8'h51; #100;
A = 8'h59; B = 8'h52; #100;
A = 8'h59; B = 8'h53; #100;
A = 8'h59; B = 8'h54; #100;
A = 8'h59; B = 8'h55; #100;
A = 8'h59; B = 8'h56; #100;
A = 8'h59; B = 8'h57; #100;
A = 8'h59; B = 8'h58; #100;
A = 8'h59; B = 8'h59; #100;
A = 8'h59; B = 8'h5A; #100;
A = 8'h59; B = 8'h5B; #100;
A = 8'h59; B = 8'h5C; #100;
A = 8'h59; B = 8'h5D; #100;
A = 8'h59; B = 8'h5E; #100;
A = 8'h59; B = 8'h5F; #100;
A = 8'h59; B = 8'h60; #100;
A = 8'h59; B = 8'h61; #100;
A = 8'h59; B = 8'h62; #100;
A = 8'h59; B = 8'h63; #100;
A = 8'h59; B = 8'h64; #100;
A = 8'h59; B = 8'h65; #100;
A = 8'h59; B = 8'h66; #100;
A = 8'h59; B = 8'h67; #100;
A = 8'h59; B = 8'h68; #100;
A = 8'h59; B = 8'h69; #100;
A = 8'h59; B = 8'h6A; #100;
A = 8'h59; B = 8'h6B; #100;
A = 8'h59; B = 8'h6C; #100;
A = 8'h59; B = 8'h6D; #100;
A = 8'h59; B = 8'h6E; #100;
A = 8'h59; B = 8'h6F; #100;
A = 8'h59; B = 8'h70; #100;
A = 8'h59; B = 8'h71; #100;
A = 8'h59; B = 8'h72; #100;
A = 8'h59; B = 8'h73; #100;
A = 8'h59; B = 8'h74; #100;
A = 8'h59; B = 8'h75; #100;
A = 8'h59; B = 8'h76; #100;
A = 8'h59; B = 8'h77; #100;
A = 8'h59; B = 8'h78; #100;
A = 8'h59; B = 8'h79; #100;
A = 8'h59; B = 8'h7A; #100;
A = 8'h59; B = 8'h7B; #100;
A = 8'h59; B = 8'h7C; #100;
A = 8'h59; B = 8'h7D; #100;
A = 8'h59; B = 8'h7E; #100;
A = 8'h59; B = 8'h7F; #100;
A = 8'h59; B = 8'h80; #100;
A = 8'h59; B = 8'h81; #100;
A = 8'h59; B = 8'h82; #100;
A = 8'h59; B = 8'h83; #100;
A = 8'h59; B = 8'h84; #100;
A = 8'h59; B = 8'h85; #100;
A = 8'h59; B = 8'h86; #100;
A = 8'h59; B = 8'h87; #100;
A = 8'h59; B = 8'h88; #100;
A = 8'h59; B = 8'h89; #100;
A = 8'h59; B = 8'h8A; #100;
A = 8'h59; B = 8'h8B; #100;
A = 8'h59; B = 8'h8C; #100;
A = 8'h59; B = 8'h8D; #100;
A = 8'h59; B = 8'h8E; #100;
A = 8'h59; B = 8'h8F; #100;
A = 8'h59; B = 8'h90; #100;
A = 8'h59; B = 8'h91; #100;
A = 8'h59; B = 8'h92; #100;
A = 8'h59; B = 8'h93; #100;
A = 8'h59; B = 8'h94; #100;
A = 8'h59; B = 8'h95; #100;
A = 8'h59; B = 8'h96; #100;
A = 8'h59; B = 8'h97; #100;
A = 8'h59; B = 8'h98; #100;
A = 8'h59; B = 8'h99; #100;
A = 8'h59; B = 8'h9A; #100;
A = 8'h59; B = 8'h9B; #100;
A = 8'h59; B = 8'h9C; #100;
A = 8'h59; B = 8'h9D; #100;
A = 8'h59; B = 8'h9E; #100;
A = 8'h59; B = 8'h9F; #100;
A = 8'h59; B = 8'hA0; #100;
A = 8'h59; B = 8'hA1; #100;
A = 8'h59; B = 8'hA2; #100;
A = 8'h59; B = 8'hA3; #100;
A = 8'h59; B = 8'hA4; #100;
A = 8'h59; B = 8'hA5; #100;
A = 8'h59; B = 8'hA6; #100;
A = 8'h59; B = 8'hA7; #100;
A = 8'h59; B = 8'hA8; #100;
A = 8'h59; B = 8'hA9; #100;
A = 8'h59; B = 8'hAA; #100;
A = 8'h59; B = 8'hAB; #100;
A = 8'h59; B = 8'hAC; #100;
A = 8'h59; B = 8'hAD; #100;
A = 8'h59; B = 8'hAE; #100;
A = 8'h59; B = 8'hAF; #100;
A = 8'h59; B = 8'hB0; #100;
A = 8'h59; B = 8'hB1; #100;
A = 8'h59; B = 8'hB2; #100;
A = 8'h59; B = 8'hB3; #100;
A = 8'h59; B = 8'hB4; #100;
A = 8'h59; B = 8'hB5; #100;
A = 8'h59; B = 8'hB6; #100;
A = 8'h59; B = 8'hB7; #100;
A = 8'h59; B = 8'hB8; #100;
A = 8'h59; B = 8'hB9; #100;
A = 8'h59; B = 8'hBA; #100;
A = 8'h59; B = 8'hBB; #100;
A = 8'h59; B = 8'hBC; #100;
A = 8'h59; B = 8'hBD; #100;
A = 8'h59; B = 8'hBE; #100;
A = 8'h59; B = 8'hBF; #100;
A = 8'h59; B = 8'hC0; #100;
A = 8'h59; B = 8'hC1; #100;
A = 8'h59; B = 8'hC2; #100;
A = 8'h59; B = 8'hC3; #100;
A = 8'h59; B = 8'hC4; #100;
A = 8'h59; B = 8'hC5; #100;
A = 8'h59; B = 8'hC6; #100;
A = 8'h59; B = 8'hC7; #100;
A = 8'h59; B = 8'hC8; #100;
A = 8'h59; B = 8'hC9; #100;
A = 8'h59; B = 8'hCA; #100;
A = 8'h59; B = 8'hCB; #100;
A = 8'h59; B = 8'hCC; #100;
A = 8'h59; B = 8'hCD; #100;
A = 8'h59; B = 8'hCE; #100;
A = 8'h59; B = 8'hCF; #100;
A = 8'h59; B = 8'hD0; #100;
A = 8'h59; B = 8'hD1; #100;
A = 8'h59; B = 8'hD2; #100;
A = 8'h59; B = 8'hD3; #100;
A = 8'h59; B = 8'hD4; #100;
A = 8'h59; B = 8'hD5; #100;
A = 8'h59; B = 8'hD6; #100;
A = 8'h59; B = 8'hD7; #100;
A = 8'h59; B = 8'hD8; #100;
A = 8'h59; B = 8'hD9; #100;
A = 8'h59; B = 8'hDA; #100;
A = 8'h59; B = 8'hDB; #100;
A = 8'h59; B = 8'hDC; #100;
A = 8'h59; B = 8'hDD; #100;
A = 8'h59; B = 8'hDE; #100;
A = 8'h59; B = 8'hDF; #100;
A = 8'h59; B = 8'hE0; #100;
A = 8'h59; B = 8'hE1; #100;
A = 8'h59; B = 8'hE2; #100;
A = 8'h59; B = 8'hE3; #100;
A = 8'h59; B = 8'hE4; #100;
A = 8'h59; B = 8'hE5; #100;
A = 8'h59; B = 8'hE6; #100;
A = 8'h59; B = 8'hE7; #100;
A = 8'h59; B = 8'hE8; #100;
A = 8'h59; B = 8'hE9; #100;
A = 8'h59; B = 8'hEA; #100;
A = 8'h59; B = 8'hEB; #100;
A = 8'h59; B = 8'hEC; #100;
A = 8'h59; B = 8'hED; #100;
A = 8'h59; B = 8'hEE; #100;
A = 8'h59; B = 8'hEF; #100;
A = 8'h59; B = 8'hF0; #100;
A = 8'h59; B = 8'hF1; #100;
A = 8'h59; B = 8'hF2; #100;
A = 8'h59; B = 8'hF3; #100;
A = 8'h59; B = 8'hF4; #100;
A = 8'h59; B = 8'hF5; #100;
A = 8'h59; B = 8'hF6; #100;
A = 8'h59; B = 8'hF7; #100;
A = 8'h59; B = 8'hF8; #100;
A = 8'h59; B = 8'hF9; #100;
A = 8'h59; B = 8'hFA; #100;
A = 8'h59; B = 8'hFB; #100;
A = 8'h59; B = 8'hFC; #100;
A = 8'h59; B = 8'hFD; #100;
A = 8'h59; B = 8'hFE; #100;
A = 8'h59; B = 8'hFF; #100;
A = 8'h5A; B = 8'h0; #100;
A = 8'h5A; B = 8'h1; #100;
A = 8'h5A; B = 8'h2; #100;
A = 8'h5A; B = 8'h3; #100;
A = 8'h5A; B = 8'h4; #100;
A = 8'h5A; B = 8'h5; #100;
A = 8'h5A; B = 8'h6; #100;
A = 8'h5A; B = 8'h7; #100;
A = 8'h5A; B = 8'h8; #100;
A = 8'h5A; B = 8'h9; #100;
A = 8'h5A; B = 8'hA; #100;
A = 8'h5A; B = 8'hB; #100;
A = 8'h5A; B = 8'hC; #100;
A = 8'h5A; B = 8'hD; #100;
A = 8'h5A; B = 8'hE; #100;
A = 8'h5A; B = 8'hF; #100;
A = 8'h5A; B = 8'h10; #100;
A = 8'h5A; B = 8'h11; #100;
A = 8'h5A; B = 8'h12; #100;
A = 8'h5A; B = 8'h13; #100;
A = 8'h5A; B = 8'h14; #100;
A = 8'h5A; B = 8'h15; #100;
A = 8'h5A; B = 8'h16; #100;
A = 8'h5A; B = 8'h17; #100;
A = 8'h5A; B = 8'h18; #100;
A = 8'h5A; B = 8'h19; #100;
A = 8'h5A; B = 8'h1A; #100;
A = 8'h5A; B = 8'h1B; #100;
A = 8'h5A; B = 8'h1C; #100;
A = 8'h5A; B = 8'h1D; #100;
A = 8'h5A; B = 8'h1E; #100;
A = 8'h5A; B = 8'h1F; #100;
A = 8'h5A; B = 8'h20; #100;
A = 8'h5A; B = 8'h21; #100;
A = 8'h5A; B = 8'h22; #100;
A = 8'h5A; B = 8'h23; #100;
A = 8'h5A; B = 8'h24; #100;
A = 8'h5A; B = 8'h25; #100;
A = 8'h5A; B = 8'h26; #100;
A = 8'h5A; B = 8'h27; #100;
A = 8'h5A; B = 8'h28; #100;
A = 8'h5A; B = 8'h29; #100;
A = 8'h5A; B = 8'h2A; #100;
A = 8'h5A; B = 8'h2B; #100;
A = 8'h5A; B = 8'h2C; #100;
A = 8'h5A; B = 8'h2D; #100;
A = 8'h5A; B = 8'h2E; #100;
A = 8'h5A; B = 8'h2F; #100;
A = 8'h5A; B = 8'h30; #100;
A = 8'h5A; B = 8'h31; #100;
A = 8'h5A; B = 8'h32; #100;
A = 8'h5A; B = 8'h33; #100;
A = 8'h5A; B = 8'h34; #100;
A = 8'h5A; B = 8'h35; #100;
A = 8'h5A; B = 8'h36; #100;
A = 8'h5A; B = 8'h37; #100;
A = 8'h5A; B = 8'h38; #100;
A = 8'h5A; B = 8'h39; #100;
A = 8'h5A; B = 8'h3A; #100;
A = 8'h5A; B = 8'h3B; #100;
A = 8'h5A; B = 8'h3C; #100;
A = 8'h5A; B = 8'h3D; #100;
A = 8'h5A; B = 8'h3E; #100;
A = 8'h5A; B = 8'h3F; #100;
A = 8'h5A; B = 8'h40; #100;
A = 8'h5A; B = 8'h41; #100;
A = 8'h5A; B = 8'h42; #100;
A = 8'h5A; B = 8'h43; #100;
A = 8'h5A; B = 8'h44; #100;
A = 8'h5A; B = 8'h45; #100;
A = 8'h5A; B = 8'h46; #100;
A = 8'h5A; B = 8'h47; #100;
A = 8'h5A; B = 8'h48; #100;
A = 8'h5A; B = 8'h49; #100;
A = 8'h5A; B = 8'h4A; #100;
A = 8'h5A; B = 8'h4B; #100;
A = 8'h5A; B = 8'h4C; #100;
A = 8'h5A; B = 8'h4D; #100;
A = 8'h5A; B = 8'h4E; #100;
A = 8'h5A; B = 8'h4F; #100;
A = 8'h5A; B = 8'h50; #100;
A = 8'h5A; B = 8'h51; #100;
A = 8'h5A; B = 8'h52; #100;
A = 8'h5A; B = 8'h53; #100;
A = 8'h5A; B = 8'h54; #100;
A = 8'h5A; B = 8'h55; #100;
A = 8'h5A; B = 8'h56; #100;
A = 8'h5A; B = 8'h57; #100;
A = 8'h5A; B = 8'h58; #100;
A = 8'h5A; B = 8'h59; #100;
A = 8'h5A; B = 8'h5A; #100;
A = 8'h5A; B = 8'h5B; #100;
A = 8'h5A; B = 8'h5C; #100;
A = 8'h5A; B = 8'h5D; #100;
A = 8'h5A; B = 8'h5E; #100;
A = 8'h5A; B = 8'h5F; #100;
A = 8'h5A; B = 8'h60; #100;
A = 8'h5A; B = 8'h61; #100;
A = 8'h5A; B = 8'h62; #100;
A = 8'h5A; B = 8'h63; #100;
A = 8'h5A; B = 8'h64; #100;
A = 8'h5A; B = 8'h65; #100;
A = 8'h5A; B = 8'h66; #100;
A = 8'h5A; B = 8'h67; #100;
A = 8'h5A; B = 8'h68; #100;
A = 8'h5A; B = 8'h69; #100;
A = 8'h5A; B = 8'h6A; #100;
A = 8'h5A; B = 8'h6B; #100;
A = 8'h5A; B = 8'h6C; #100;
A = 8'h5A; B = 8'h6D; #100;
A = 8'h5A; B = 8'h6E; #100;
A = 8'h5A; B = 8'h6F; #100;
A = 8'h5A; B = 8'h70; #100;
A = 8'h5A; B = 8'h71; #100;
A = 8'h5A; B = 8'h72; #100;
A = 8'h5A; B = 8'h73; #100;
A = 8'h5A; B = 8'h74; #100;
A = 8'h5A; B = 8'h75; #100;
A = 8'h5A; B = 8'h76; #100;
A = 8'h5A; B = 8'h77; #100;
A = 8'h5A; B = 8'h78; #100;
A = 8'h5A; B = 8'h79; #100;
A = 8'h5A; B = 8'h7A; #100;
A = 8'h5A; B = 8'h7B; #100;
A = 8'h5A; B = 8'h7C; #100;
A = 8'h5A; B = 8'h7D; #100;
A = 8'h5A; B = 8'h7E; #100;
A = 8'h5A; B = 8'h7F; #100;
A = 8'h5A; B = 8'h80; #100;
A = 8'h5A; B = 8'h81; #100;
A = 8'h5A; B = 8'h82; #100;
A = 8'h5A; B = 8'h83; #100;
A = 8'h5A; B = 8'h84; #100;
A = 8'h5A; B = 8'h85; #100;
A = 8'h5A; B = 8'h86; #100;
A = 8'h5A; B = 8'h87; #100;
A = 8'h5A; B = 8'h88; #100;
A = 8'h5A; B = 8'h89; #100;
A = 8'h5A; B = 8'h8A; #100;
A = 8'h5A; B = 8'h8B; #100;
A = 8'h5A; B = 8'h8C; #100;
A = 8'h5A; B = 8'h8D; #100;
A = 8'h5A; B = 8'h8E; #100;
A = 8'h5A; B = 8'h8F; #100;
A = 8'h5A; B = 8'h90; #100;
A = 8'h5A; B = 8'h91; #100;
A = 8'h5A; B = 8'h92; #100;
A = 8'h5A; B = 8'h93; #100;
A = 8'h5A; B = 8'h94; #100;
A = 8'h5A; B = 8'h95; #100;
A = 8'h5A; B = 8'h96; #100;
A = 8'h5A; B = 8'h97; #100;
A = 8'h5A; B = 8'h98; #100;
A = 8'h5A; B = 8'h99; #100;
A = 8'h5A; B = 8'h9A; #100;
A = 8'h5A; B = 8'h9B; #100;
A = 8'h5A; B = 8'h9C; #100;
A = 8'h5A; B = 8'h9D; #100;
A = 8'h5A; B = 8'h9E; #100;
A = 8'h5A; B = 8'h9F; #100;
A = 8'h5A; B = 8'hA0; #100;
A = 8'h5A; B = 8'hA1; #100;
A = 8'h5A; B = 8'hA2; #100;
A = 8'h5A; B = 8'hA3; #100;
A = 8'h5A; B = 8'hA4; #100;
A = 8'h5A; B = 8'hA5; #100;
A = 8'h5A; B = 8'hA6; #100;
A = 8'h5A; B = 8'hA7; #100;
A = 8'h5A; B = 8'hA8; #100;
A = 8'h5A; B = 8'hA9; #100;
A = 8'h5A; B = 8'hAA; #100;
A = 8'h5A; B = 8'hAB; #100;
A = 8'h5A; B = 8'hAC; #100;
A = 8'h5A; B = 8'hAD; #100;
A = 8'h5A; B = 8'hAE; #100;
A = 8'h5A; B = 8'hAF; #100;
A = 8'h5A; B = 8'hB0; #100;
A = 8'h5A; B = 8'hB1; #100;
A = 8'h5A; B = 8'hB2; #100;
A = 8'h5A; B = 8'hB3; #100;
A = 8'h5A; B = 8'hB4; #100;
A = 8'h5A; B = 8'hB5; #100;
A = 8'h5A; B = 8'hB6; #100;
A = 8'h5A; B = 8'hB7; #100;
A = 8'h5A; B = 8'hB8; #100;
A = 8'h5A; B = 8'hB9; #100;
A = 8'h5A; B = 8'hBA; #100;
A = 8'h5A; B = 8'hBB; #100;
A = 8'h5A; B = 8'hBC; #100;
A = 8'h5A; B = 8'hBD; #100;
A = 8'h5A; B = 8'hBE; #100;
A = 8'h5A; B = 8'hBF; #100;
A = 8'h5A; B = 8'hC0; #100;
A = 8'h5A; B = 8'hC1; #100;
A = 8'h5A; B = 8'hC2; #100;
A = 8'h5A; B = 8'hC3; #100;
A = 8'h5A; B = 8'hC4; #100;
A = 8'h5A; B = 8'hC5; #100;
A = 8'h5A; B = 8'hC6; #100;
A = 8'h5A; B = 8'hC7; #100;
A = 8'h5A; B = 8'hC8; #100;
A = 8'h5A; B = 8'hC9; #100;
A = 8'h5A; B = 8'hCA; #100;
A = 8'h5A; B = 8'hCB; #100;
A = 8'h5A; B = 8'hCC; #100;
A = 8'h5A; B = 8'hCD; #100;
A = 8'h5A; B = 8'hCE; #100;
A = 8'h5A; B = 8'hCF; #100;
A = 8'h5A; B = 8'hD0; #100;
A = 8'h5A; B = 8'hD1; #100;
A = 8'h5A; B = 8'hD2; #100;
A = 8'h5A; B = 8'hD3; #100;
A = 8'h5A; B = 8'hD4; #100;
A = 8'h5A; B = 8'hD5; #100;
A = 8'h5A; B = 8'hD6; #100;
A = 8'h5A; B = 8'hD7; #100;
A = 8'h5A; B = 8'hD8; #100;
A = 8'h5A; B = 8'hD9; #100;
A = 8'h5A; B = 8'hDA; #100;
A = 8'h5A; B = 8'hDB; #100;
A = 8'h5A; B = 8'hDC; #100;
A = 8'h5A; B = 8'hDD; #100;
A = 8'h5A; B = 8'hDE; #100;
A = 8'h5A; B = 8'hDF; #100;
A = 8'h5A; B = 8'hE0; #100;
A = 8'h5A; B = 8'hE1; #100;
A = 8'h5A; B = 8'hE2; #100;
A = 8'h5A; B = 8'hE3; #100;
A = 8'h5A; B = 8'hE4; #100;
A = 8'h5A; B = 8'hE5; #100;
A = 8'h5A; B = 8'hE6; #100;
A = 8'h5A; B = 8'hE7; #100;
A = 8'h5A; B = 8'hE8; #100;
A = 8'h5A; B = 8'hE9; #100;
A = 8'h5A; B = 8'hEA; #100;
A = 8'h5A; B = 8'hEB; #100;
A = 8'h5A; B = 8'hEC; #100;
A = 8'h5A; B = 8'hED; #100;
A = 8'h5A; B = 8'hEE; #100;
A = 8'h5A; B = 8'hEF; #100;
A = 8'h5A; B = 8'hF0; #100;
A = 8'h5A; B = 8'hF1; #100;
A = 8'h5A; B = 8'hF2; #100;
A = 8'h5A; B = 8'hF3; #100;
A = 8'h5A; B = 8'hF4; #100;
A = 8'h5A; B = 8'hF5; #100;
A = 8'h5A; B = 8'hF6; #100;
A = 8'h5A; B = 8'hF7; #100;
A = 8'h5A; B = 8'hF8; #100;
A = 8'h5A; B = 8'hF9; #100;
A = 8'h5A; B = 8'hFA; #100;
A = 8'h5A; B = 8'hFB; #100;
A = 8'h5A; B = 8'hFC; #100;
A = 8'h5A; B = 8'hFD; #100;
A = 8'h5A; B = 8'hFE; #100;
A = 8'h5A; B = 8'hFF; #100;
A = 8'h5B; B = 8'h0; #100;
A = 8'h5B; B = 8'h1; #100;
A = 8'h5B; B = 8'h2; #100;
A = 8'h5B; B = 8'h3; #100;
A = 8'h5B; B = 8'h4; #100;
A = 8'h5B; B = 8'h5; #100;
A = 8'h5B; B = 8'h6; #100;
A = 8'h5B; B = 8'h7; #100;
A = 8'h5B; B = 8'h8; #100;
A = 8'h5B; B = 8'h9; #100;
A = 8'h5B; B = 8'hA; #100;
A = 8'h5B; B = 8'hB; #100;
A = 8'h5B; B = 8'hC; #100;
A = 8'h5B; B = 8'hD; #100;
A = 8'h5B; B = 8'hE; #100;
A = 8'h5B; B = 8'hF; #100;
A = 8'h5B; B = 8'h10; #100;
A = 8'h5B; B = 8'h11; #100;
A = 8'h5B; B = 8'h12; #100;
A = 8'h5B; B = 8'h13; #100;
A = 8'h5B; B = 8'h14; #100;
A = 8'h5B; B = 8'h15; #100;
A = 8'h5B; B = 8'h16; #100;
A = 8'h5B; B = 8'h17; #100;
A = 8'h5B; B = 8'h18; #100;
A = 8'h5B; B = 8'h19; #100;
A = 8'h5B; B = 8'h1A; #100;
A = 8'h5B; B = 8'h1B; #100;
A = 8'h5B; B = 8'h1C; #100;
A = 8'h5B; B = 8'h1D; #100;
A = 8'h5B; B = 8'h1E; #100;
A = 8'h5B; B = 8'h1F; #100;
A = 8'h5B; B = 8'h20; #100;
A = 8'h5B; B = 8'h21; #100;
A = 8'h5B; B = 8'h22; #100;
A = 8'h5B; B = 8'h23; #100;
A = 8'h5B; B = 8'h24; #100;
A = 8'h5B; B = 8'h25; #100;
A = 8'h5B; B = 8'h26; #100;
A = 8'h5B; B = 8'h27; #100;
A = 8'h5B; B = 8'h28; #100;
A = 8'h5B; B = 8'h29; #100;
A = 8'h5B; B = 8'h2A; #100;
A = 8'h5B; B = 8'h2B; #100;
A = 8'h5B; B = 8'h2C; #100;
A = 8'h5B; B = 8'h2D; #100;
A = 8'h5B; B = 8'h2E; #100;
A = 8'h5B; B = 8'h2F; #100;
A = 8'h5B; B = 8'h30; #100;
A = 8'h5B; B = 8'h31; #100;
A = 8'h5B; B = 8'h32; #100;
A = 8'h5B; B = 8'h33; #100;
A = 8'h5B; B = 8'h34; #100;
A = 8'h5B; B = 8'h35; #100;
A = 8'h5B; B = 8'h36; #100;
A = 8'h5B; B = 8'h37; #100;
A = 8'h5B; B = 8'h38; #100;
A = 8'h5B; B = 8'h39; #100;
A = 8'h5B; B = 8'h3A; #100;
A = 8'h5B; B = 8'h3B; #100;
A = 8'h5B; B = 8'h3C; #100;
A = 8'h5B; B = 8'h3D; #100;
A = 8'h5B; B = 8'h3E; #100;
A = 8'h5B; B = 8'h3F; #100;
A = 8'h5B; B = 8'h40; #100;
A = 8'h5B; B = 8'h41; #100;
A = 8'h5B; B = 8'h42; #100;
A = 8'h5B; B = 8'h43; #100;
A = 8'h5B; B = 8'h44; #100;
A = 8'h5B; B = 8'h45; #100;
A = 8'h5B; B = 8'h46; #100;
A = 8'h5B; B = 8'h47; #100;
A = 8'h5B; B = 8'h48; #100;
A = 8'h5B; B = 8'h49; #100;
A = 8'h5B; B = 8'h4A; #100;
A = 8'h5B; B = 8'h4B; #100;
A = 8'h5B; B = 8'h4C; #100;
A = 8'h5B; B = 8'h4D; #100;
A = 8'h5B; B = 8'h4E; #100;
A = 8'h5B; B = 8'h4F; #100;
A = 8'h5B; B = 8'h50; #100;
A = 8'h5B; B = 8'h51; #100;
A = 8'h5B; B = 8'h52; #100;
A = 8'h5B; B = 8'h53; #100;
A = 8'h5B; B = 8'h54; #100;
A = 8'h5B; B = 8'h55; #100;
A = 8'h5B; B = 8'h56; #100;
A = 8'h5B; B = 8'h57; #100;
A = 8'h5B; B = 8'h58; #100;
A = 8'h5B; B = 8'h59; #100;
A = 8'h5B; B = 8'h5A; #100;
A = 8'h5B; B = 8'h5B; #100;
A = 8'h5B; B = 8'h5C; #100;
A = 8'h5B; B = 8'h5D; #100;
A = 8'h5B; B = 8'h5E; #100;
A = 8'h5B; B = 8'h5F; #100;
A = 8'h5B; B = 8'h60; #100;
A = 8'h5B; B = 8'h61; #100;
A = 8'h5B; B = 8'h62; #100;
A = 8'h5B; B = 8'h63; #100;
A = 8'h5B; B = 8'h64; #100;
A = 8'h5B; B = 8'h65; #100;
A = 8'h5B; B = 8'h66; #100;
A = 8'h5B; B = 8'h67; #100;
A = 8'h5B; B = 8'h68; #100;
A = 8'h5B; B = 8'h69; #100;
A = 8'h5B; B = 8'h6A; #100;
A = 8'h5B; B = 8'h6B; #100;
A = 8'h5B; B = 8'h6C; #100;
A = 8'h5B; B = 8'h6D; #100;
A = 8'h5B; B = 8'h6E; #100;
A = 8'h5B; B = 8'h6F; #100;
A = 8'h5B; B = 8'h70; #100;
A = 8'h5B; B = 8'h71; #100;
A = 8'h5B; B = 8'h72; #100;
A = 8'h5B; B = 8'h73; #100;
A = 8'h5B; B = 8'h74; #100;
A = 8'h5B; B = 8'h75; #100;
A = 8'h5B; B = 8'h76; #100;
A = 8'h5B; B = 8'h77; #100;
A = 8'h5B; B = 8'h78; #100;
A = 8'h5B; B = 8'h79; #100;
A = 8'h5B; B = 8'h7A; #100;
A = 8'h5B; B = 8'h7B; #100;
A = 8'h5B; B = 8'h7C; #100;
A = 8'h5B; B = 8'h7D; #100;
A = 8'h5B; B = 8'h7E; #100;
A = 8'h5B; B = 8'h7F; #100;
A = 8'h5B; B = 8'h80; #100;
A = 8'h5B; B = 8'h81; #100;
A = 8'h5B; B = 8'h82; #100;
A = 8'h5B; B = 8'h83; #100;
A = 8'h5B; B = 8'h84; #100;
A = 8'h5B; B = 8'h85; #100;
A = 8'h5B; B = 8'h86; #100;
A = 8'h5B; B = 8'h87; #100;
A = 8'h5B; B = 8'h88; #100;
A = 8'h5B; B = 8'h89; #100;
A = 8'h5B; B = 8'h8A; #100;
A = 8'h5B; B = 8'h8B; #100;
A = 8'h5B; B = 8'h8C; #100;
A = 8'h5B; B = 8'h8D; #100;
A = 8'h5B; B = 8'h8E; #100;
A = 8'h5B; B = 8'h8F; #100;
A = 8'h5B; B = 8'h90; #100;
A = 8'h5B; B = 8'h91; #100;
A = 8'h5B; B = 8'h92; #100;
A = 8'h5B; B = 8'h93; #100;
A = 8'h5B; B = 8'h94; #100;
A = 8'h5B; B = 8'h95; #100;
A = 8'h5B; B = 8'h96; #100;
A = 8'h5B; B = 8'h97; #100;
A = 8'h5B; B = 8'h98; #100;
A = 8'h5B; B = 8'h99; #100;
A = 8'h5B; B = 8'h9A; #100;
A = 8'h5B; B = 8'h9B; #100;
A = 8'h5B; B = 8'h9C; #100;
A = 8'h5B; B = 8'h9D; #100;
A = 8'h5B; B = 8'h9E; #100;
A = 8'h5B; B = 8'h9F; #100;
A = 8'h5B; B = 8'hA0; #100;
A = 8'h5B; B = 8'hA1; #100;
A = 8'h5B; B = 8'hA2; #100;
A = 8'h5B; B = 8'hA3; #100;
A = 8'h5B; B = 8'hA4; #100;
A = 8'h5B; B = 8'hA5; #100;
A = 8'h5B; B = 8'hA6; #100;
A = 8'h5B; B = 8'hA7; #100;
A = 8'h5B; B = 8'hA8; #100;
A = 8'h5B; B = 8'hA9; #100;
A = 8'h5B; B = 8'hAA; #100;
A = 8'h5B; B = 8'hAB; #100;
A = 8'h5B; B = 8'hAC; #100;
A = 8'h5B; B = 8'hAD; #100;
A = 8'h5B; B = 8'hAE; #100;
A = 8'h5B; B = 8'hAF; #100;
A = 8'h5B; B = 8'hB0; #100;
A = 8'h5B; B = 8'hB1; #100;
A = 8'h5B; B = 8'hB2; #100;
A = 8'h5B; B = 8'hB3; #100;
A = 8'h5B; B = 8'hB4; #100;
A = 8'h5B; B = 8'hB5; #100;
A = 8'h5B; B = 8'hB6; #100;
A = 8'h5B; B = 8'hB7; #100;
A = 8'h5B; B = 8'hB8; #100;
A = 8'h5B; B = 8'hB9; #100;
A = 8'h5B; B = 8'hBA; #100;
A = 8'h5B; B = 8'hBB; #100;
A = 8'h5B; B = 8'hBC; #100;
A = 8'h5B; B = 8'hBD; #100;
A = 8'h5B; B = 8'hBE; #100;
A = 8'h5B; B = 8'hBF; #100;
A = 8'h5B; B = 8'hC0; #100;
A = 8'h5B; B = 8'hC1; #100;
A = 8'h5B; B = 8'hC2; #100;
A = 8'h5B; B = 8'hC3; #100;
A = 8'h5B; B = 8'hC4; #100;
A = 8'h5B; B = 8'hC5; #100;
A = 8'h5B; B = 8'hC6; #100;
A = 8'h5B; B = 8'hC7; #100;
A = 8'h5B; B = 8'hC8; #100;
A = 8'h5B; B = 8'hC9; #100;
A = 8'h5B; B = 8'hCA; #100;
A = 8'h5B; B = 8'hCB; #100;
A = 8'h5B; B = 8'hCC; #100;
A = 8'h5B; B = 8'hCD; #100;
A = 8'h5B; B = 8'hCE; #100;
A = 8'h5B; B = 8'hCF; #100;
A = 8'h5B; B = 8'hD0; #100;
A = 8'h5B; B = 8'hD1; #100;
A = 8'h5B; B = 8'hD2; #100;
A = 8'h5B; B = 8'hD3; #100;
A = 8'h5B; B = 8'hD4; #100;
A = 8'h5B; B = 8'hD5; #100;
A = 8'h5B; B = 8'hD6; #100;
A = 8'h5B; B = 8'hD7; #100;
A = 8'h5B; B = 8'hD8; #100;
A = 8'h5B; B = 8'hD9; #100;
A = 8'h5B; B = 8'hDA; #100;
A = 8'h5B; B = 8'hDB; #100;
A = 8'h5B; B = 8'hDC; #100;
A = 8'h5B; B = 8'hDD; #100;
A = 8'h5B; B = 8'hDE; #100;
A = 8'h5B; B = 8'hDF; #100;
A = 8'h5B; B = 8'hE0; #100;
A = 8'h5B; B = 8'hE1; #100;
A = 8'h5B; B = 8'hE2; #100;
A = 8'h5B; B = 8'hE3; #100;
A = 8'h5B; B = 8'hE4; #100;
A = 8'h5B; B = 8'hE5; #100;
A = 8'h5B; B = 8'hE6; #100;
A = 8'h5B; B = 8'hE7; #100;
A = 8'h5B; B = 8'hE8; #100;
A = 8'h5B; B = 8'hE9; #100;
A = 8'h5B; B = 8'hEA; #100;
A = 8'h5B; B = 8'hEB; #100;
A = 8'h5B; B = 8'hEC; #100;
A = 8'h5B; B = 8'hED; #100;
A = 8'h5B; B = 8'hEE; #100;
A = 8'h5B; B = 8'hEF; #100;
A = 8'h5B; B = 8'hF0; #100;
A = 8'h5B; B = 8'hF1; #100;
A = 8'h5B; B = 8'hF2; #100;
A = 8'h5B; B = 8'hF3; #100;
A = 8'h5B; B = 8'hF4; #100;
A = 8'h5B; B = 8'hF5; #100;
A = 8'h5B; B = 8'hF6; #100;
A = 8'h5B; B = 8'hF7; #100;
A = 8'h5B; B = 8'hF8; #100;
A = 8'h5B; B = 8'hF9; #100;
A = 8'h5B; B = 8'hFA; #100;
A = 8'h5B; B = 8'hFB; #100;
A = 8'h5B; B = 8'hFC; #100;
A = 8'h5B; B = 8'hFD; #100;
A = 8'h5B; B = 8'hFE; #100;
A = 8'h5B; B = 8'hFF; #100;
A = 8'h5C; B = 8'h0; #100;
A = 8'h5C; B = 8'h1; #100;
A = 8'h5C; B = 8'h2; #100;
A = 8'h5C; B = 8'h3; #100;
A = 8'h5C; B = 8'h4; #100;
A = 8'h5C; B = 8'h5; #100;
A = 8'h5C; B = 8'h6; #100;
A = 8'h5C; B = 8'h7; #100;
A = 8'h5C; B = 8'h8; #100;
A = 8'h5C; B = 8'h9; #100;
A = 8'h5C; B = 8'hA; #100;
A = 8'h5C; B = 8'hB; #100;
A = 8'h5C; B = 8'hC; #100;
A = 8'h5C; B = 8'hD; #100;
A = 8'h5C; B = 8'hE; #100;
A = 8'h5C; B = 8'hF; #100;
A = 8'h5C; B = 8'h10; #100;
A = 8'h5C; B = 8'h11; #100;
A = 8'h5C; B = 8'h12; #100;
A = 8'h5C; B = 8'h13; #100;
A = 8'h5C; B = 8'h14; #100;
A = 8'h5C; B = 8'h15; #100;
A = 8'h5C; B = 8'h16; #100;
A = 8'h5C; B = 8'h17; #100;
A = 8'h5C; B = 8'h18; #100;
A = 8'h5C; B = 8'h19; #100;
A = 8'h5C; B = 8'h1A; #100;
A = 8'h5C; B = 8'h1B; #100;
A = 8'h5C; B = 8'h1C; #100;
A = 8'h5C; B = 8'h1D; #100;
A = 8'h5C; B = 8'h1E; #100;
A = 8'h5C; B = 8'h1F; #100;
A = 8'h5C; B = 8'h20; #100;
A = 8'h5C; B = 8'h21; #100;
A = 8'h5C; B = 8'h22; #100;
A = 8'h5C; B = 8'h23; #100;
A = 8'h5C; B = 8'h24; #100;
A = 8'h5C; B = 8'h25; #100;
A = 8'h5C; B = 8'h26; #100;
A = 8'h5C; B = 8'h27; #100;
A = 8'h5C; B = 8'h28; #100;
A = 8'h5C; B = 8'h29; #100;
A = 8'h5C; B = 8'h2A; #100;
A = 8'h5C; B = 8'h2B; #100;
A = 8'h5C; B = 8'h2C; #100;
A = 8'h5C; B = 8'h2D; #100;
A = 8'h5C; B = 8'h2E; #100;
A = 8'h5C; B = 8'h2F; #100;
A = 8'h5C; B = 8'h30; #100;
A = 8'h5C; B = 8'h31; #100;
A = 8'h5C; B = 8'h32; #100;
A = 8'h5C; B = 8'h33; #100;
A = 8'h5C; B = 8'h34; #100;
A = 8'h5C; B = 8'h35; #100;
A = 8'h5C; B = 8'h36; #100;
A = 8'h5C; B = 8'h37; #100;
A = 8'h5C; B = 8'h38; #100;
A = 8'h5C; B = 8'h39; #100;
A = 8'h5C; B = 8'h3A; #100;
A = 8'h5C; B = 8'h3B; #100;
A = 8'h5C; B = 8'h3C; #100;
A = 8'h5C; B = 8'h3D; #100;
A = 8'h5C; B = 8'h3E; #100;
A = 8'h5C; B = 8'h3F; #100;
A = 8'h5C; B = 8'h40; #100;
A = 8'h5C; B = 8'h41; #100;
A = 8'h5C; B = 8'h42; #100;
A = 8'h5C; B = 8'h43; #100;
A = 8'h5C; B = 8'h44; #100;
A = 8'h5C; B = 8'h45; #100;
A = 8'h5C; B = 8'h46; #100;
A = 8'h5C; B = 8'h47; #100;
A = 8'h5C; B = 8'h48; #100;
A = 8'h5C; B = 8'h49; #100;
A = 8'h5C; B = 8'h4A; #100;
A = 8'h5C; B = 8'h4B; #100;
A = 8'h5C; B = 8'h4C; #100;
A = 8'h5C; B = 8'h4D; #100;
A = 8'h5C; B = 8'h4E; #100;
A = 8'h5C; B = 8'h4F; #100;
A = 8'h5C; B = 8'h50; #100;
A = 8'h5C; B = 8'h51; #100;
A = 8'h5C; B = 8'h52; #100;
A = 8'h5C; B = 8'h53; #100;
A = 8'h5C; B = 8'h54; #100;
A = 8'h5C; B = 8'h55; #100;
A = 8'h5C; B = 8'h56; #100;
A = 8'h5C; B = 8'h57; #100;
A = 8'h5C; B = 8'h58; #100;
A = 8'h5C; B = 8'h59; #100;
A = 8'h5C; B = 8'h5A; #100;
A = 8'h5C; B = 8'h5B; #100;
A = 8'h5C; B = 8'h5C; #100;
A = 8'h5C; B = 8'h5D; #100;
A = 8'h5C; B = 8'h5E; #100;
A = 8'h5C; B = 8'h5F; #100;
A = 8'h5C; B = 8'h60; #100;
A = 8'h5C; B = 8'h61; #100;
A = 8'h5C; B = 8'h62; #100;
A = 8'h5C; B = 8'h63; #100;
A = 8'h5C; B = 8'h64; #100;
A = 8'h5C; B = 8'h65; #100;
A = 8'h5C; B = 8'h66; #100;
A = 8'h5C; B = 8'h67; #100;
A = 8'h5C; B = 8'h68; #100;
A = 8'h5C; B = 8'h69; #100;
A = 8'h5C; B = 8'h6A; #100;
A = 8'h5C; B = 8'h6B; #100;
A = 8'h5C; B = 8'h6C; #100;
A = 8'h5C; B = 8'h6D; #100;
A = 8'h5C; B = 8'h6E; #100;
A = 8'h5C; B = 8'h6F; #100;
A = 8'h5C; B = 8'h70; #100;
A = 8'h5C; B = 8'h71; #100;
A = 8'h5C; B = 8'h72; #100;
A = 8'h5C; B = 8'h73; #100;
A = 8'h5C; B = 8'h74; #100;
A = 8'h5C; B = 8'h75; #100;
A = 8'h5C; B = 8'h76; #100;
A = 8'h5C; B = 8'h77; #100;
A = 8'h5C; B = 8'h78; #100;
A = 8'h5C; B = 8'h79; #100;
A = 8'h5C; B = 8'h7A; #100;
A = 8'h5C; B = 8'h7B; #100;
A = 8'h5C; B = 8'h7C; #100;
A = 8'h5C; B = 8'h7D; #100;
A = 8'h5C; B = 8'h7E; #100;
A = 8'h5C; B = 8'h7F; #100;
A = 8'h5C; B = 8'h80; #100;
A = 8'h5C; B = 8'h81; #100;
A = 8'h5C; B = 8'h82; #100;
A = 8'h5C; B = 8'h83; #100;
A = 8'h5C; B = 8'h84; #100;
A = 8'h5C; B = 8'h85; #100;
A = 8'h5C; B = 8'h86; #100;
A = 8'h5C; B = 8'h87; #100;
A = 8'h5C; B = 8'h88; #100;
A = 8'h5C; B = 8'h89; #100;
A = 8'h5C; B = 8'h8A; #100;
A = 8'h5C; B = 8'h8B; #100;
A = 8'h5C; B = 8'h8C; #100;
A = 8'h5C; B = 8'h8D; #100;
A = 8'h5C; B = 8'h8E; #100;
A = 8'h5C; B = 8'h8F; #100;
A = 8'h5C; B = 8'h90; #100;
A = 8'h5C; B = 8'h91; #100;
A = 8'h5C; B = 8'h92; #100;
A = 8'h5C; B = 8'h93; #100;
A = 8'h5C; B = 8'h94; #100;
A = 8'h5C; B = 8'h95; #100;
A = 8'h5C; B = 8'h96; #100;
A = 8'h5C; B = 8'h97; #100;
A = 8'h5C; B = 8'h98; #100;
A = 8'h5C; B = 8'h99; #100;
A = 8'h5C; B = 8'h9A; #100;
A = 8'h5C; B = 8'h9B; #100;
A = 8'h5C; B = 8'h9C; #100;
A = 8'h5C; B = 8'h9D; #100;
A = 8'h5C; B = 8'h9E; #100;
A = 8'h5C; B = 8'h9F; #100;
A = 8'h5C; B = 8'hA0; #100;
A = 8'h5C; B = 8'hA1; #100;
A = 8'h5C; B = 8'hA2; #100;
A = 8'h5C; B = 8'hA3; #100;
A = 8'h5C; B = 8'hA4; #100;
A = 8'h5C; B = 8'hA5; #100;
A = 8'h5C; B = 8'hA6; #100;
A = 8'h5C; B = 8'hA7; #100;
A = 8'h5C; B = 8'hA8; #100;
A = 8'h5C; B = 8'hA9; #100;
A = 8'h5C; B = 8'hAA; #100;
A = 8'h5C; B = 8'hAB; #100;
A = 8'h5C; B = 8'hAC; #100;
A = 8'h5C; B = 8'hAD; #100;
A = 8'h5C; B = 8'hAE; #100;
A = 8'h5C; B = 8'hAF; #100;
A = 8'h5C; B = 8'hB0; #100;
A = 8'h5C; B = 8'hB1; #100;
A = 8'h5C; B = 8'hB2; #100;
A = 8'h5C; B = 8'hB3; #100;
A = 8'h5C; B = 8'hB4; #100;
A = 8'h5C; B = 8'hB5; #100;
A = 8'h5C; B = 8'hB6; #100;
A = 8'h5C; B = 8'hB7; #100;
A = 8'h5C; B = 8'hB8; #100;
A = 8'h5C; B = 8'hB9; #100;
A = 8'h5C; B = 8'hBA; #100;
A = 8'h5C; B = 8'hBB; #100;
A = 8'h5C; B = 8'hBC; #100;
A = 8'h5C; B = 8'hBD; #100;
A = 8'h5C; B = 8'hBE; #100;
A = 8'h5C; B = 8'hBF; #100;
A = 8'h5C; B = 8'hC0; #100;
A = 8'h5C; B = 8'hC1; #100;
A = 8'h5C; B = 8'hC2; #100;
A = 8'h5C; B = 8'hC3; #100;
A = 8'h5C; B = 8'hC4; #100;
A = 8'h5C; B = 8'hC5; #100;
A = 8'h5C; B = 8'hC6; #100;
A = 8'h5C; B = 8'hC7; #100;
A = 8'h5C; B = 8'hC8; #100;
A = 8'h5C; B = 8'hC9; #100;
A = 8'h5C; B = 8'hCA; #100;
A = 8'h5C; B = 8'hCB; #100;
A = 8'h5C; B = 8'hCC; #100;
A = 8'h5C; B = 8'hCD; #100;
A = 8'h5C; B = 8'hCE; #100;
A = 8'h5C; B = 8'hCF; #100;
A = 8'h5C; B = 8'hD0; #100;
A = 8'h5C; B = 8'hD1; #100;
A = 8'h5C; B = 8'hD2; #100;
A = 8'h5C; B = 8'hD3; #100;
A = 8'h5C; B = 8'hD4; #100;
A = 8'h5C; B = 8'hD5; #100;
A = 8'h5C; B = 8'hD6; #100;
A = 8'h5C; B = 8'hD7; #100;
A = 8'h5C; B = 8'hD8; #100;
A = 8'h5C; B = 8'hD9; #100;
A = 8'h5C; B = 8'hDA; #100;
A = 8'h5C; B = 8'hDB; #100;
A = 8'h5C; B = 8'hDC; #100;
A = 8'h5C; B = 8'hDD; #100;
A = 8'h5C; B = 8'hDE; #100;
A = 8'h5C; B = 8'hDF; #100;
A = 8'h5C; B = 8'hE0; #100;
A = 8'h5C; B = 8'hE1; #100;
A = 8'h5C; B = 8'hE2; #100;
A = 8'h5C; B = 8'hE3; #100;
A = 8'h5C; B = 8'hE4; #100;
A = 8'h5C; B = 8'hE5; #100;
A = 8'h5C; B = 8'hE6; #100;
A = 8'h5C; B = 8'hE7; #100;
A = 8'h5C; B = 8'hE8; #100;
A = 8'h5C; B = 8'hE9; #100;
A = 8'h5C; B = 8'hEA; #100;
A = 8'h5C; B = 8'hEB; #100;
A = 8'h5C; B = 8'hEC; #100;
A = 8'h5C; B = 8'hED; #100;
A = 8'h5C; B = 8'hEE; #100;
A = 8'h5C; B = 8'hEF; #100;
A = 8'h5C; B = 8'hF0; #100;
A = 8'h5C; B = 8'hF1; #100;
A = 8'h5C; B = 8'hF2; #100;
A = 8'h5C; B = 8'hF3; #100;
A = 8'h5C; B = 8'hF4; #100;
A = 8'h5C; B = 8'hF5; #100;
A = 8'h5C; B = 8'hF6; #100;
A = 8'h5C; B = 8'hF7; #100;
A = 8'h5C; B = 8'hF8; #100;
A = 8'h5C; B = 8'hF9; #100;
A = 8'h5C; B = 8'hFA; #100;
A = 8'h5C; B = 8'hFB; #100;
A = 8'h5C; B = 8'hFC; #100;
A = 8'h5C; B = 8'hFD; #100;
A = 8'h5C; B = 8'hFE; #100;
A = 8'h5C; B = 8'hFF; #100;
A = 8'h5D; B = 8'h0; #100;
A = 8'h5D; B = 8'h1; #100;
A = 8'h5D; B = 8'h2; #100;
A = 8'h5D; B = 8'h3; #100;
A = 8'h5D; B = 8'h4; #100;
A = 8'h5D; B = 8'h5; #100;
A = 8'h5D; B = 8'h6; #100;
A = 8'h5D; B = 8'h7; #100;
A = 8'h5D; B = 8'h8; #100;
A = 8'h5D; B = 8'h9; #100;
A = 8'h5D; B = 8'hA; #100;
A = 8'h5D; B = 8'hB; #100;
A = 8'h5D; B = 8'hC; #100;
A = 8'h5D; B = 8'hD; #100;
A = 8'h5D; B = 8'hE; #100;
A = 8'h5D; B = 8'hF; #100;
A = 8'h5D; B = 8'h10; #100;
A = 8'h5D; B = 8'h11; #100;
A = 8'h5D; B = 8'h12; #100;
A = 8'h5D; B = 8'h13; #100;
A = 8'h5D; B = 8'h14; #100;
A = 8'h5D; B = 8'h15; #100;
A = 8'h5D; B = 8'h16; #100;
A = 8'h5D; B = 8'h17; #100;
A = 8'h5D; B = 8'h18; #100;
A = 8'h5D; B = 8'h19; #100;
A = 8'h5D; B = 8'h1A; #100;
A = 8'h5D; B = 8'h1B; #100;
A = 8'h5D; B = 8'h1C; #100;
A = 8'h5D; B = 8'h1D; #100;
A = 8'h5D; B = 8'h1E; #100;
A = 8'h5D; B = 8'h1F; #100;
A = 8'h5D; B = 8'h20; #100;
A = 8'h5D; B = 8'h21; #100;
A = 8'h5D; B = 8'h22; #100;
A = 8'h5D; B = 8'h23; #100;
A = 8'h5D; B = 8'h24; #100;
A = 8'h5D; B = 8'h25; #100;
A = 8'h5D; B = 8'h26; #100;
A = 8'h5D; B = 8'h27; #100;
A = 8'h5D; B = 8'h28; #100;
A = 8'h5D; B = 8'h29; #100;
A = 8'h5D; B = 8'h2A; #100;
A = 8'h5D; B = 8'h2B; #100;
A = 8'h5D; B = 8'h2C; #100;
A = 8'h5D; B = 8'h2D; #100;
A = 8'h5D; B = 8'h2E; #100;
A = 8'h5D; B = 8'h2F; #100;
A = 8'h5D; B = 8'h30; #100;
A = 8'h5D; B = 8'h31; #100;
A = 8'h5D; B = 8'h32; #100;
A = 8'h5D; B = 8'h33; #100;
A = 8'h5D; B = 8'h34; #100;
A = 8'h5D; B = 8'h35; #100;
A = 8'h5D; B = 8'h36; #100;
A = 8'h5D; B = 8'h37; #100;
A = 8'h5D; B = 8'h38; #100;
A = 8'h5D; B = 8'h39; #100;
A = 8'h5D; B = 8'h3A; #100;
A = 8'h5D; B = 8'h3B; #100;
A = 8'h5D; B = 8'h3C; #100;
A = 8'h5D; B = 8'h3D; #100;
A = 8'h5D; B = 8'h3E; #100;
A = 8'h5D; B = 8'h3F; #100;
A = 8'h5D; B = 8'h40; #100;
A = 8'h5D; B = 8'h41; #100;
A = 8'h5D; B = 8'h42; #100;
A = 8'h5D; B = 8'h43; #100;
A = 8'h5D; B = 8'h44; #100;
A = 8'h5D; B = 8'h45; #100;
A = 8'h5D; B = 8'h46; #100;
A = 8'h5D; B = 8'h47; #100;
A = 8'h5D; B = 8'h48; #100;
A = 8'h5D; B = 8'h49; #100;
A = 8'h5D; B = 8'h4A; #100;
A = 8'h5D; B = 8'h4B; #100;
A = 8'h5D; B = 8'h4C; #100;
A = 8'h5D; B = 8'h4D; #100;
A = 8'h5D; B = 8'h4E; #100;
A = 8'h5D; B = 8'h4F; #100;
A = 8'h5D; B = 8'h50; #100;
A = 8'h5D; B = 8'h51; #100;
A = 8'h5D; B = 8'h52; #100;
A = 8'h5D; B = 8'h53; #100;
A = 8'h5D; B = 8'h54; #100;
A = 8'h5D; B = 8'h55; #100;
A = 8'h5D; B = 8'h56; #100;
A = 8'h5D; B = 8'h57; #100;
A = 8'h5D; B = 8'h58; #100;
A = 8'h5D; B = 8'h59; #100;
A = 8'h5D; B = 8'h5A; #100;
A = 8'h5D; B = 8'h5B; #100;
A = 8'h5D; B = 8'h5C; #100;
A = 8'h5D; B = 8'h5D; #100;
A = 8'h5D; B = 8'h5E; #100;
A = 8'h5D; B = 8'h5F; #100;
A = 8'h5D; B = 8'h60; #100;
A = 8'h5D; B = 8'h61; #100;
A = 8'h5D; B = 8'h62; #100;
A = 8'h5D; B = 8'h63; #100;
A = 8'h5D; B = 8'h64; #100;
A = 8'h5D; B = 8'h65; #100;
A = 8'h5D; B = 8'h66; #100;
A = 8'h5D; B = 8'h67; #100;
A = 8'h5D; B = 8'h68; #100;
A = 8'h5D; B = 8'h69; #100;
A = 8'h5D; B = 8'h6A; #100;
A = 8'h5D; B = 8'h6B; #100;
A = 8'h5D; B = 8'h6C; #100;
A = 8'h5D; B = 8'h6D; #100;
A = 8'h5D; B = 8'h6E; #100;
A = 8'h5D; B = 8'h6F; #100;
A = 8'h5D; B = 8'h70; #100;
A = 8'h5D; B = 8'h71; #100;
A = 8'h5D; B = 8'h72; #100;
A = 8'h5D; B = 8'h73; #100;
A = 8'h5D; B = 8'h74; #100;
A = 8'h5D; B = 8'h75; #100;
A = 8'h5D; B = 8'h76; #100;
A = 8'h5D; B = 8'h77; #100;
A = 8'h5D; B = 8'h78; #100;
A = 8'h5D; B = 8'h79; #100;
A = 8'h5D; B = 8'h7A; #100;
A = 8'h5D; B = 8'h7B; #100;
A = 8'h5D; B = 8'h7C; #100;
A = 8'h5D; B = 8'h7D; #100;
A = 8'h5D; B = 8'h7E; #100;
A = 8'h5D; B = 8'h7F; #100;
A = 8'h5D; B = 8'h80; #100;
A = 8'h5D; B = 8'h81; #100;
A = 8'h5D; B = 8'h82; #100;
A = 8'h5D; B = 8'h83; #100;
A = 8'h5D; B = 8'h84; #100;
A = 8'h5D; B = 8'h85; #100;
A = 8'h5D; B = 8'h86; #100;
A = 8'h5D; B = 8'h87; #100;
A = 8'h5D; B = 8'h88; #100;
A = 8'h5D; B = 8'h89; #100;
A = 8'h5D; B = 8'h8A; #100;
A = 8'h5D; B = 8'h8B; #100;
A = 8'h5D; B = 8'h8C; #100;
A = 8'h5D; B = 8'h8D; #100;
A = 8'h5D; B = 8'h8E; #100;
A = 8'h5D; B = 8'h8F; #100;
A = 8'h5D; B = 8'h90; #100;
A = 8'h5D; B = 8'h91; #100;
A = 8'h5D; B = 8'h92; #100;
A = 8'h5D; B = 8'h93; #100;
A = 8'h5D; B = 8'h94; #100;
A = 8'h5D; B = 8'h95; #100;
A = 8'h5D; B = 8'h96; #100;
A = 8'h5D; B = 8'h97; #100;
A = 8'h5D; B = 8'h98; #100;
A = 8'h5D; B = 8'h99; #100;
A = 8'h5D; B = 8'h9A; #100;
A = 8'h5D; B = 8'h9B; #100;
A = 8'h5D; B = 8'h9C; #100;
A = 8'h5D; B = 8'h9D; #100;
A = 8'h5D; B = 8'h9E; #100;
A = 8'h5D; B = 8'h9F; #100;
A = 8'h5D; B = 8'hA0; #100;
A = 8'h5D; B = 8'hA1; #100;
A = 8'h5D; B = 8'hA2; #100;
A = 8'h5D; B = 8'hA3; #100;
A = 8'h5D; B = 8'hA4; #100;
A = 8'h5D; B = 8'hA5; #100;
A = 8'h5D; B = 8'hA6; #100;
A = 8'h5D; B = 8'hA7; #100;
A = 8'h5D; B = 8'hA8; #100;
A = 8'h5D; B = 8'hA9; #100;
A = 8'h5D; B = 8'hAA; #100;
A = 8'h5D; B = 8'hAB; #100;
A = 8'h5D; B = 8'hAC; #100;
A = 8'h5D; B = 8'hAD; #100;
A = 8'h5D; B = 8'hAE; #100;
A = 8'h5D; B = 8'hAF; #100;
A = 8'h5D; B = 8'hB0; #100;
A = 8'h5D; B = 8'hB1; #100;
A = 8'h5D; B = 8'hB2; #100;
A = 8'h5D; B = 8'hB3; #100;
A = 8'h5D; B = 8'hB4; #100;
A = 8'h5D; B = 8'hB5; #100;
A = 8'h5D; B = 8'hB6; #100;
A = 8'h5D; B = 8'hB7; #100;
A = 8'h5D; B = 8'hB8; #100;
A = 8'h5D; B = 8'hB9; #100;
A = 8'h5D; B = 8'hBA; #100;
A = 8'h5D; B = 8'hBB; #100;
A = 8'h5D; B = 8'hBC; #100;
A = 8'h5D; B = 8'hBD; #100;
A = 8'h5D; B = 8'hBE; #100;
A = 8'h5D; B = 8'hBF; #100;
A = 8'h5D; B = 8'hC0; #100;
A = 8'h5D; B = 8'hC1; #100;
A = 8'h5D; B = 8'hC2; #100;
A = 8'h5D; B = 8'hC3; #100;
A = 8'h5D; B = 8'hC4; #100;
A = 8'h5D; B = 8'hC5; #100;
A = 8'h5D; B = 8'hC6; #100;
A = 8'h5D; B = 8'hC7; #100;
A = 8'h5D; B = 8'hC8; #100;
A = 8'h5D; B = 8'hC9; #100;
A = 8'h5D; B = 8'hCA; #100;
A = 8'h5D; B = 8'hCB; #100;
A = 8'h5D; B = 8'hCC; #100;
A = 8'h5D; B = 8'hCD; #100;
A = 8'h5D; B = 8'hCE; #100;
A = 8'h5D; B = 8'hCF; #100;
A = 8'h5D; B = 8'hD0; #100;
A = 8'h5D; B = 8'hD1; #100;
A = 8'h5D; B = 8'hD2; #100;
A = 8'h5D; B = 8'hD3; #100;
A = 8'h5D; B = 8'hD4; #100;
A = 8'h5D; B = 8'hD5; #100;
A = 8'h5D; B = 8'hD6; #100;
A = 8'h5D; B = 8'hD7; #100;
A = 8'h5D; B = 8'hD8; #100;
A = 8'h5D; B = 8'hD9; #100;
A = 8'h5D; B = 8'hDA; #100;
A = 8'h5D; B = 8'hDB; #100;
A = 8'h5D; B = 8'hDC; #100;
A = 8'h5D; B = 8'hDD; #100;
A = 8'h5D; B = 8'hDE; #100;
A = 8'h5D; B = 8'hDF; #100;
A = 8'h5D; B = 8'hE0; #100;
A = 8'h5D; B = 8'hE1; #100;
A = 8'h5D; B = 8'hE2; #100;
A = 8'h5D; B = 8'hE3; #100;
A = 8'h5D; B = 8'hE4; #100;
A = 8'h5D; B = 8'hE5; #100;
A = 8'h5D; B = 8'hE6; #100;
A = 8'h5D; B = 8'hE7; #100;
A = 8'h5D; B = 8'hE8; #100;
A = 8'h5D; B = 8'hE9; #100;
A = 8'h5D; B = 8'hEA; #100;
A = 8'h5D; B = 8'hEB; #100;
A = 8'h5D; B = 8'hEC; #100;
A = 8'h5D; B = 8'hED; #100;
A = 8'h5D; B = 8'hEE; #100;
A = 8'h5D; B = 8'hEF; #100;
A = 8'h5D; B = 8'hF0; #100;
A = 8'h5D; B = 8'hF1; #100;
A = 8'h5D; B = 8'hF2; #100;
A = 8'h5D; B = 8'hF3; #100;
A = 8'h5D; B = 8'hF4; #100;
A = 8'h5D; B = 8'hF5; #100;
A = 8'h5D; B = 8'hF6; #100;
A = 8'h5D; B = 8'hF7; #100;
A = 8'h5D; B = 8'hF8; #100;
A = 8'h5D; B = 8'hF9; #100;
A = 8'h5D; B = 8'hFA; #100;
A = 8'h5D; B = 8'hFB; #100;
A = 8'h5D; B = 8'hFC; #100;
A = 8'h5D; B = 8'hFD; #100;
A = 8'h5D; B = 8'hFE; #100;
A = 8'h5D; B = 8'hFF; #100;
A = 8'h5E; B = 8'h0; #100;
A = 8'h5E; B = 8'h1; #100;
A = 8'h5E; B = 8'h2; #100;
A = 8'h5E; B = 8'h3; #100;
A = 8'h5E; B = 8'h4; #100;
A = 8'h5E; B = 8'h5; #100;
A = 8'h5E; B = 8'h6; #100;
A = 8'h5E; B = 8'h7; #100;
A = 8'h5E; B = 8'h8; #100;
A = 8'h5E; B = 8'h9; #100;
A = 8'h5E; B = 8'hA; #100;
A = 8'h5E; B = 8'hB; #100;
A = 8'h5E; B = 8'hC; #100;
A = 8'h5E; B = 8'hD; #100;
A = 8'h5E; B = 8'hE; #100;
A = 8'h5E; B = 8'hF; #100;
A = 8'h5E; B = 8'h10; #100;
A = 8'h5E; B = 8'h11; #100;
A = 8'h5E; B = 8'h12; #100;
A = 8'h5E; B = 8'h13; #100;
A = 8'h5E; B = 8'h14; #100;
A = 8'h5E; B = 8'h15; #100;
A = 8'h5E; B = 8'h16; #100;
A = 8'h5E; B = 8'h17; #100;
A = 8'h5E; B = 8'h18; #100;
A = 8'h5E; B = 8'h19; #100;
A = 8'h5E; B = 8'h1A; #100;
A = 8'h5E; B = 8'h1B; #100;
A = 8'h5E; B = 8'h1C; #100;
A = 8'h5E; B = 8'h1D; #100;
A = 8'h5E; B = 8'h1E; #100;
A = 8'h5E; B = 8'h1F; #100;
A = 8'h5E; B = 8'h20; #100;
A = 8'h5E; B = 8'h21; #100;
A = 8'h5E; B = 8'h22; #100;
A = 8'h5E; B = 8'h23; #100;
A = 8'h5E; B = 8'h24; #100;
A = 8'h5E; B = 8'h25; #100;
A = 8'h5E; B = 8'h26; #100;
A = 8'h5E; B = 8'h27; #100;
A = 8'h5E; B = 8'h28; #100;
A = 8'h5E; B = 8'h29; #100;
A = 8'h5E; B = 8'h2A; #100;
A = 8'h5E; B = 8'h2B; #100;
A = 8'h5E; B = 8'h2C; #100;
A = 8'h5E; B = 8'h2D; #100;
A = 8'h5E; B = 8'h2E; #100;
A = 8'h5E; B = 8'h2F; #100;
A = 8'h5E; B = 8'h30; #100;
A = 8'h5E; B = 8'h31; #100;
A = 8'h5E; B = 8'h32; #100;
A = 8'h5E; B = 8'h33; #100;
A = 8'h5E; B = 8'h34; #100;
A = 8'h5E; B = 8'h35; #100;
A = 8'h5E; B = 8'h36; #100;
A = 8'h5E; B = 8'h37; #100;
A = 8'h5E; B = 8'h38; #100;
A = 8'h5E; B = 8'h39; #100;
A = 8'h5E; B = 8'h3A; #100;
A = 8'h5E; B = 8'h3B; #100;
A = 8'h5E; B = 8'h3C; #100;
A = 8'h5E; B = 8'h3D; #100;
A = 8'h5E; B = 8'h3E; #100;
A = 8'h5E; B = 8'h3F; #100;
A = 8'h5E; B = 8'h40; #100;
A = 8'h5E; B = 8'h41; #100;
A = 8'h5E; B = 8'h42; #100;
A = 8'h5E; B = 8'h43; #100;
A = 8'h5E; B = 8'h44; #100;
A = 8'h5E; B = 8'h45; #100;
A = 8'h5E; B = 8'h46; #100;
A = 8'h5E; B = 8'h47; #100;
A = 8'h5E; B = 8'h48; #100;
A = 8'h5E; B = 8'h49; #100;
A = 8'h5E; B = 8'h4A; #100;
A = 8'h5E; B = 8'h4B; #100;
A = 8'h5E; B = 8'h4C; #100;
A = 8'h5E; B = 8'h4D; #100;
A = 8'h5E; B = 8'h4E; #100;
A = 8'h5E; B = 8'h4F; #100;
A = 8'h5E; B = 8'h50; #100;
A = 8'h5E; B = 8'h51; #100;
A = 8'h5E; B = 8'h52; #100;
A = 8'h5E; B = 8'h53; #100;
A = 8'h5E; B = 8'h54; #100;
A = 8'h5E; B = 8'h55; #100;
A = 8'h5E; B = 8'h56; #100;
A = 8'h5E; B = 8'h57; #100;
A = 8'h5E; B = 8'h58; #100;
A = 8'h5E; B = 8'h59; #100;
A = 8'h5E; B = 8'h5A; #100;
A = 8'h5E; B = 8'h5B; #100;
A = 8'h5E; B = 8'h5C; #100;
A = 8'h5E; B = 8'h5D; #100;
A = 8'h5E; B = 8'h5E; #100;
A = 8'h5E; B = 8'h5F; #100;
A = 8'h5E; B = 8'h60; #100;
A = 8'h5E; B = 8'h61; #100;
A = 8'h5E; B = 8'h62; #100;
A = 8'h5E; B = 8'h63; #100;
A = 8'h5E; B = 8'h64; #100;
A = 8'h5E; B = 8'h65; #100;
A = 8'h5E; B = 8'h66; #100;
A = 8'h5E; B = 8'h67; #100;
A = 8'h5E; B = 8'h68; #100;
A = 8'h5E; B = 8'h69; #100;
A = 8'h5E; B = 8'h6A; #100;
A = 8'h5E; B = 8'h6B; #100;
A = 8'h5E; B = 8'h6C; #100;
A = 8'h5E; B = 8'h6D; #100;
A = 8'h5E; B = 8'h6E; #100;
A = 8'h5E; B = 8'h6F; #100;
A = 8'h5E; B = 8'h70; #100;
A = 8'h5E; B = 8'h71; #100;
A = 8'h5E; B = 8'h72; #100;
A = 8'h5E; B = 8'h73; #100;
A = 8'h5E; B = 8'h74; #100;
A = 8'h5E; B = 8'h75; #100;
A = 8'h5E; B = 8'h76; #100;
A = 8'h5E; B = 8'h77; #100;
A = 8'h5E; B = 8'h78; #100;
A = 8'h5E; B = 8'h79; #100;
A = 8'h5E; B = 8'h7A; #100;
A = 8'h5E; B = 8'h7B; #100;
A = 8'h5E; B = 8'h7C; #100;
A = 8'h5E; B = 8'h7D; #100;
A = 8'h5E; B = 8'h7E; #100;
A = 8'h5E; B = 8'h7F; #100;
A = 8'h5E; B = 8'h80; #100;
A = 8'h5E; B = 8'h81; #100;
A = 8'h5E; B = 8'h82; #100;
A = 8'h5E; B = 8'h83; #100;
A = 8'h5E; B = 8'h84; #100;
A = 8'h5E; B = 8'h85; #100;
A = 8'h5E; B = 8'h86; #100;
A = 8'h5E; B = 8'h87; #100;
A = 8'h5E; B = 8'h88; #100;
A = 8'h5E; B = 8'h89; #100;
A = 8'h5E; B = 8'h8A; #100;
A = 8'h5E; B = 8'h8B; #100;
A = 8'h5E; B = 8'h8C; #100;
A = 8'h5E; B = 8'h8D; #100;
A = 8'h5E; B = 8'h8E; #100;
A = 8'h5E; B = 8'h8F; #100;
A = 8'h5E; B = 8'h90; #100;
A = 8'h5E; B = 8'h91; #100;
A = 8'h5E; B = 8'h92; #100;
A = 8'h5E; B = 8'h93; #100;
A = 8'h5E; B = 8'h94; #100;
A = 8'h5E; B = 8'h95; #100;
A = 8'h5E; B = 8'h96; #100;
A = 8'h5E; B = 8'h97; #100;
A = 8'h5E; B = 8'h98; #100;
A = 8'h5E; B = 8'h99; #100;
A = 8'h5E; B = 8'h9A; #100;
A = 8'h5E; B = 8'h9B; #100;
A = 8'h5E; B = 8'h9C; #100;
A = 8'h5E; B = 8'h9D; #100;
A = 8'h5E; B = 8'h9E; #100;
A = 8'h5E; B = 8'h9F; #100;
A = 8'h5E; B = 8'hA0; #100;
A = 8'h5E; B = 8'hA1; #100;
A = 8'h5E; B = 8'hA2; #100;
A = 8'h5E; B = 8'hA3; #100;
A = 8'h5E; B = 8'hA4; #100;
A = 8'h5E; B = 8'hA5; #100;
A = 8'h5E; B = 8'hA6; #100;
A = 8'h5E; B = 8'hA7; #100;
A = 8'h5E; B = 8'hA8; #100;
A = 8'h5E; B = 8'hA9; #100;
A = 8'h5E; B = 8'hAA; #100;
A = 8'h5E; B = 8'hAB; #100;
A = 8'h5E; B = 8'hAC; #100;
A = 8'h5E; B = 8'hAD; #100;
A = 8'h5E; B = 8'hAE; #100;
A = 8'h5E; B = 8'hAF; #100;
A = 8'h5E; B = 8'hB0; #100;
A = 8'h5E; B = 8'hB1; #100;
A = 8'h5E; B = 8'hB2; #100;
A = 8'h5E; B = 8'hB3; #100;
A = 8'h5E; B = 8'hB4; #100;
A = 8'h5E; B = 8'hB5; #100;
A = 8'h5E; B = 8'hB6; #100;
A = 8'h5E; B = 8'hB7; #100;
A = 8'h5E; B = 8'hB8; #100;
A = 8'h5E; B = 8'hB9; #100;
A = 8'h5E; B = 8'hBA; #100;
A = 8'h5E; B = 8'hBB; #100;
A = 8'h5E; B = 8'hBC; #100;
A = 8'h5E; B = 8'hBD; #100;
A = 8'h5E; B = 8'hBE; #100;
A = 8'h5E; B = 8'hBF; #100;
A = 8'h5E; B = 8'hC0; #100;
A = 8'h5E; B = 8'hC1; #100;
A = 8'h5E; B = 8'hC2; #100;
A = 8'h5E; B = 8'hC3; #100;
A = 8'h5E; B = 8'hC4; #100;
A = 8'h5E; B = 8'hC5; #100;
A = 8'h5E; B = 8'hC6; #100;
A = 8'h5E; B = 8'hC7; #100;
A = 8'h5E; B = 8'hC8; #100;
A = 8'h5E; B = 8'hC9; #100;
A = 8'h5E; B = 8'hCA; #100;
A = 8'h5E; B = 8'hCB; #100;
A = 8'h5E; B = 8'hCC; #100;
A = 8'h5E; B = 8'hCD; #100;
A = 8'h5E; B = 8'hCE; #100;
A = 8'h5E; B = 8'hCF; #100;
A = 8'h5E; B = 8'hD0; #100;
A = 8'h5E; B = 8'hD1; #100;
A = 8'h5E; B = 8'hD2; #100;
A = 8'h5E; B = 8'hD3; #100;
A = 8'h5E; B = 8'hD4; #100;
A = 8'h5E; B = 8'hD5; #100;
A = 8'h5E; B = 8'hD6; #100;
A = 8'h5E; B = 8'hD7; #100;
A = 8'h5E; B = 8'hD8; #100;
A = 8'h5E; B = 8'hD9; #100;
A = 8'h5E; B = 8'hDA; #100;
A = 8'h5E; B = 8'hDB; #100;
A = 8'h5E; B = 8'hDC; #100;
A = 8'h5E; B = 8'hDD; #100;
A = 8'h5E; B = 8'hDE; #100;
A = 8'h5E; B = 8'hDF; #100;
A = 8'h5E; B = 8'hE0; #100;
A = 8'h5E; B = 8'hE1; #100;
A = 8'h5E; B = 8'hE2; #100;
A = 8'h5E; B = 8'hE3; #100;
A = 8'h5E; B = 8'hE4; #100;
A = 8'h5E; B = 8'hE5; #100;
A = 8'h5E; B = 8'hE6; #100;
A = 8'h5E; B = 8'hE7; #100;
A = 8'h5E; B = 8'hE8; #100;
A = 8'h5E; B = 8'hE9; #100;
A = 8'h5E; B = 8'hEA; #100;
A = 8'h5E; B = 8'hEB; #100;
A = 8'h5E; B = 8'hEC; #100;
A = 8'h5E; B = 8'hED; #100;
A = 8'h5E; B = 8'hEE; #100;
A = 8'h5E; B = 8'hEF; #100;
A = 8'h5E; B = 8'hF0; #100;
A = 8'h5E; B = 8'hF1; #100;
A = 8'h5E; B = 8'hF2; #100;
A = 8'h5E; B = 8'hF3; #100;
A = 8'h5E; B = 8'hF4; #100;
A = 8'h5E; B = 8'hF5; #100;
A = 8'h5E; B = 8'hF6; #100;
A = 8'h5E; B = 8'hF7; #100;
A = 8'h5E; B = 8'hF8; #100;
A = 8'h5E; B = 8'hF9; #100;
A = 8'h5E; B = 8'hFA; #100;
A = 8'h5E; B = 8'hFB; #100;
A = 8'h5E; B = 8'hFC; #100;
A = 8'h5E; B = 8'hFD; #100;
A = 8'h5E; B = 8'hFE; #100;
A = 8'h5E; B = 8'hFF; #100;
A = 8'h5F; B = 8'h0; #100;
A = 8'h5F; B = 8'h1; #100;
A = 8'h5F; B = 8'h2; #100;
A = 8'h5F; B = 8'h3; #100;
A = 8'h5F; B = 8'h4; #100;
A = 8'h5F; B = 8'h5; #100;
A = 8'h5F; B = 8'h6; #100;
A = 8'h5F; B = 8'h7; #100;
A = 8'h5F; B = 8'h8; #100;
A = 8'h5F; B = 8'h9; #100;
A = 8'h5F; B = 8'hA; #100;
A = 8'h5F; B = 8'hB; #100;
A = 8'h5F; B = 8'hC; #100;
A = 8'h5F; B = 8'hD; #100;
A = 8'h5F; B = 8'hE; #100;
A = 8'h5F; B = 8'hF; #100;
A = 8'h5F; B = 8'h10; #100;
A = 8'h5F; B = 8'h11; #100;
A = 8'h5F; B = 8'h12; #100;
A = 8'h5F; B = 8'h13; #100;
A = 8'h5F; B = 8'h14; #100;
A = 8'h5F; B = 8'h15; #100;
A = 8'h5F; B = 8'h16; #100;
A = 8'h5F; B = 8'h17; #100;
A = 8'h5F; B = 8'h18; #100;
A = 8'h5F; B = 8'h19; #100;
A = 8'h5F; B = 8'h1A; #100;
A = 8'h5F; B = 8'h1B; #100;
A = 8'h5F; B = 8'h1C; #100;
A = 8'h5F; B = 8'h1D; #100;
A = 8'h5F; B = 8'h1E; #100;
A = 8'h5F; B = 8'h1F; #100;
A = 8'h5F; B = 8'h20; #100;
A = 8'h5F; B = 8'h21; #100;
A = 8'h5F; B = 8'h22; #100;
A = 8'h5F; B = 8'h23; #100;
A = 8'h5F; B = 8'h24; #100;
A = 8'h5F; B = 8'h25; #100;
A = 8'h5F; B = 8'h26; #100;
A = 8'h5F; B = 8'h27; #100;
A = 8'h5F; B = 8'h28; #100;
A = 8'h5F; B = 8'h29; #100;
A = 8'h5F; B = 8'h2A; #100;
A = 8'h5F; B = 8'h2B; #100;
A = 8'h5F; B = 8'h2C; #100;
A = 8'h5F; B = 8'h2D; #100;
A = 8'h5F; B = 8'h2E; #100;
A = 8'h5F; B = 8'h2F; #100;
A = 8'h5F; B = 8'h30; #100;
A = 8'h5F; B = 8'h31; #100;
A = 8'h5F; B = 8'h32; #100;
A = 8'h5F; B = 8'h33; #100;
A = 8'h5F; B = 8'h34; #100;
A = 8'h5F; B = 8'h35; #100;
A = 8'h5F; B = 8'h36; #100;
A = 8'h5F; B = 8'h37; #100;
A = 8'h5F; B = 8'h38; #100;
A = 8'h5F; B = 8'h39; #100;
A = 8'h5F; B = 8'h3A; #100;
A = 8'h5F; B = 8'h3B; #100;
A = 8'h5F; B = 8'h3C; #100;
A = 8'h5F; B = 8'h3D; #100;
A = 8'h5F; B = 8'h3E; #100;
A = 8'h5F; B = 8'h3F; #100;
A = 8'h5F; B = 8'h40; #100;
A = 8'h5F; B = 8'h41; #100;
A = 8'h5F; B = 8'h42; #100;
A = 8'h5F; B = 8'h43; #100;
A = 8'h5F; B = 8'h44; #100;
A = 8'h5F; B = 8'h45; #100;
A = 8'h5F; B = 8'h46; #100;
A = 8'h5F; B = 8'h47; #100;
A = 8'h5F; B = 8'h48; #100;
A = 8'h5F; B = 8'h49; #100;
A = 8'h5F; B = 8'h4A; #100;
A = 8'h5F; B = 8'h4B; #100;
A = 8'h5F; B = 8'h4C; #100;
A = 8'h5F; B = 8'h4D; #100;
A = 8'h5F; B = 8'h4E; #100;
A = 8'h5F; B = 8'h4F; #100;
A = 8'h5F; B = 8'h50; #100;
A = 8'h5F; B = 8'h51; #100;
A = 8'h5F; B = 8'h52; #100;
A = 8'h5F; B = 8'h53; #100;
A = 8'h5F; B = 8'h54; #100;
A = 8'h5F; B = 8'h55; #100;
A = 8'h5F; B = 8'h56; #100;
A = 8'h5F; B = 8'h57; #100;
A = 8'h5F; B = 8'h58; #100;
A = 8'h5F; B = 8'h59; #100;
A = 8'h5F; B = 8'h5A; #100;
A = 8'h5F; B = 8'h5B; #100;
A = 8'h5F; B = 8'h5C; #100;
A = 8'h5F; B = 8'h5D; #100;
A = 8'h5F; B = 8'h5E; #100;
A = 8'h5F; B = 8'h5F; #100;
A = 8'h5F; B = 8'h60; #100;
A = 8'h5F; B = 8'h61; #100;
A = 8'h5F; B = 8'h62; #100;
A = 8'h5F; B = 8'h63; #100;
A = 8'h5F; B = 8'h64; #100;
A = 8'h5F; B = 8'h65; #100;
A = 8'h5F; B = 8'h66; #100;
A = 8'h5F; B = 8'h67; #100;
A = 8'h5F; B = 8'h68; #100;
A = 8'h5F; B = 8'h69; #100;
A = 8'h5F; B = 8'h6A; #100;
A = 8'h5F; B = 8'h6B; #100;
A = 8'h5F; B = 8'h6C; #100;
A = 8'h5F; B = 8'h6D; #100;
A = 8'h5F; B = 8'h6E; #100;
A = 8'h5F; B = 8'h6F; #100;
A = 8'h5F; B = 8'h70; #100;
A = 8'h5F; B = 8'h71; #100;
A = 8'h5F; B = 8'h72; #100;
A = 8'h5F; B = 8'h73; #100;
A = 8'h5F; B = 8'h74; #100;
A = 8'h5F; B = 8'h75; #100;
A = 8'h5F; B = 8'h76; #100;
A = 8'h5F; B = 8'h77; #100;
A = 8'h5F; B = 8'h78; #100;
A = 8'h5F; B = 8'h79; #100;
A = 8'h5F; B = 8'h7A; #100;
A = 8'h5F; B = 8'h7B; #100;
A = 8'h5F; B = 8'h7C; #100;
A = 8'h5F; B = 8'h7D; #100;
A = 8'h5F; B = 8'h7E; #100;
A = 8'h5F; B = 8'h7F; #100;
A = 8'h5F; B = 8'h80; #100;
A = 8'h5F; B = 8'h81; #100;
A = 8'h5F; B = 8'h82; #100;
A = 8'h5F; B = 8'h83; #100;
A = 8'h5F; B = 8'h84; #100;
A = 8'h5F; B = 8'h85; #100;
A = 8'h5F; B = 8'h86; #100;
A = 8'h5F; B = 8'h87; #100;
A = 8'h5F; B = 8'h88; #100;
A = 8'h5F; B = 8'h89; #100;
A = 8'h5F; B = 8'h8A; #100;
A = 8'h5F; B = 8'h8B; #100;
A = 8'h5F; B = 8'h8C; #100;
A = 8'h5F; B = 8'h8D; #100;
A = 8'h5F; B = 8'h8E; #100;
A = 8'h5F; B = 8'h8F; #100;
A = 8'h5F; B = 8'h90; #100;
A = 8'h5F; B = 8'h91; #100;
A = 8'h5F; B = 8'h92; #100;
A = 8'h5F; B = 8'h93; #100;
A = 8'h5F; B = 8'h94; #100;
A = 8'h5F; B = 8'h95; #100;
A = 8'h5F; B = 8'h96; #100;
A = 8'h5F; B = 8'h97; #100;
A = 8'h5F; B = 8'h98; #100;
A = 8'h5F; B = 8'h99; #100;
A = 8'h5F; B = 8'h9A; #100;
A = 8'h5F; B = 8'h9B; #100;
A = 8'h5F; B = 8'h9C; #100;
A = 8'h5F; B = 8'h9D; #100;
A = 8'h5F; B = 8'h9E; #100;
A = 8'h5F; B = 8'h9F; #100;
A = 8'h5F; B = 8'hA0; #100;
A = 8'h5F; B = 8'hA1; #100;
A = 8'h5F; B = 8'hA2; #100;
A = 8'h5F; B = 8'hA3; #100;
A = 8'h5F; B = 8'hA4; #100;
A = 8'h5F; B = 8'hA5; #100;
A = 8'h5F; B = 8'hA6; #100;
A = 8'h5F; B = 8'hA7; #100;
A = 8'h5F; B = 8'hA8; #100;
A = 8'h5F; B = 8'hA9; #100;
A = 8'h5F; B = 8'hAA; #100;
A = 8'h5F; B = 8'hAB; #100;
A = 8'h5F; B = 8'hAC; #100;
A = 8'h5F; B = 8'hAD; #100;
A = 8'h5F; B = 8'hAE; #100;
A = 8'h5F; B = 8'hAF; #100;
A = 8'h5F; B = 8'hB0; #100;
A = 8'h5F; B = 8'hB1; #100;
A = 8'h5F; B = 8'hB2; #100;
A = 8'h5F; B = 8'hB3; #100;
A = 8'h5F; B = 8'hB4; #100;
A = 8'h5F; B = 8'hB5; #100;
A = 8'h5F; B = 8'hB6; #100;
A = 8'h5F; B = 8'hB7; #100;
A = 8'h5F; B = 8'hB8; #100;
A = 8'h5F; B = 8'hB9; #100;
A = 8'h5F; B = 8'hBA; #100;
A = 8'h5F; B = 8'hBB; #100;
A = 8'h5F; B = 8'hBC; #100;
A = 8'h5F; B = 8'hBD; #100;
A = 8'h5F; B = 8'hBE; #100;
A = 8'h5F; B = 8'hBF; #100;
A = 8'h5F; B = 8'hC0; #100;
A = 8'h5F; B = 8'hC1; #100;
A = 8'h5F; B = 8'hC2; #100;
A = 8'h5F; B = 8'hC3; #100;
A = 8'h5F; B = 8'hC4; #100;
A = 8'h5F; B = 8'hC5; #100;
A = 8'h5F; B = 8'hC6; #100;
A = 8'h5F; B = 8'hC7; #100;
A = 8'h5F; B = 8'hC8; #100;
A = 8'h5F; B = 8'hC9; #100;
A = 8'h5F; B = 8'hCA; #100;
A = 8'h5F; B = 8'hCB; #100;
A = 8'h5F; B = 8'hCC; #100;
A = 8'h5F; B = 8'hCD; #100;
A = 8'h5F; B = 8'hCE; #100;
A = 8'h5F; B = 8'hCF; #100;
A = 8'h5F; B = 8'hD0; #100;
A = 8'h5F; B = 8'hD1; #100;
A = 8'h5F; B = 8'hD2; #100;
A = 8'h5F; B = 8'hD3; #100;
A = 8'h5F; B = 8'hD4; #100;
A = 8'h5F; B = 8'hD5; #100;
A = 8'h5F; B = 8'hD6; #100;
A = 8'h5F; B = 8'hD7; #100;
A = 8'h5F; B = 8'hD8; #100;
A = 8'h5F; B = 8'hD9; #100;
A = 8'h5F; B = 8'hDA; #100;
A = 8'h5F; B = 8'hDB; #100;
A = 8'h5F; B = 8'hDC; #100;
A = 8'h5F; B = 8'hDD; #100;
A = 8'h5F; B = 8'hDE; #100;
A = 8'h5F; B = 8'hDF; #100;
A = 8'h5F; B = 8'hE0; #100;
A = 8'h5F; B = 8'hE1; #100;
A = 8'h5F; B = 8'hE2; #100;
A = 8'h5F; B = 8'hE3; #100;
A = 8'h5F; B = 8'hE4; #100;
A = 8'h5F; B = 8'hE5; #100;
A = 8'h5F; B = 8'hE6; #100;
A = 8'h5F; B = 8'hE7; #100;
A = 8'h5F; B = 8'hE8; #100;
A = 8'h5F; B = 8'hE9; #100;
A = 8'h5F; B = 8'hEA; #100;
A = 8'h5F; B = 8'hEB; #100;
A = 8'h5F; B = 8'hEC; #100;
A = 8'h5F; B = 8'hED; #100;
A = 8'h5F; B = 8'hEE; #100;
A = 8'h5F; B = 8'hEF; #100;
A = 8'h5F; B = 8'hF0; #100;
A = 8'h5F; B = 8'hF1; #100;
A = 8'h5F; B = 8'hF2; #100;
A = 8'h5F; B = 8'hF3; #100;
A = 8'h5F; B = 8'hF4; #100;
A = 8'h5F; B = 8'hF5; #100;
A = 8'h5F; B = 8'hF6; #100;
A = 8'h5F; B = 8'hF7; #100;
A = 8'h5F; B = 8'hF8; #100;
A = 8'h5F; B = 8'hF9; #100;
A = 8'h5F; B = 8'hFA; #100;
A = 8'h5F; B = 8'hFB; #100;
A = 8'h5F; B = 8'hFC; #100;
A = 8'h5F; B = 8'hFD; #100;
A = 8'h5F; B = 8'hFE; #100;
A = 8'h5F; B = 8'hFF; #100;
A = 8'h60; B = 8'h0; #100;
A = 8'h60; B = 8'h1; #100;
A = 8'h60; B = 8'h2; #100;
A = 8'h60; B = 8'h3; #100;
A = 8'h60; B = 8'h4; #100;
A = 8'h60; B = 8'h5; #100;
A = 8'h60; B = 8'h6; #100;
A = 8'h60; B = 8'h7; #100;
A = 8'h60; B = 8'h8; #100;
A = 8'h60; B = 8'h9; #100;
A = 8'h60; B = 8'hA; #100;
A = 8'h60; B = 8'hB; #100;
A = 8'h60; B = 8'hC; #100;
A = 8'h60; B = 8'hD; #100;
A = 8'h60; B = 8'hE; #100;
A = 8'h60; B = 8'hF; #100;
A = 8'h60; B = 8'h10; #100;
A = 8'h60; B = 8'h11; #100;
A = 8'h60; B = 8'h12; #100;
A = 8'h60; B = 8'h13; #100;
A = 8'h60; B = 8'h14; #100;
A = 8'h60; B = 8'h15; #100;
A = 8'h60; B = 8'h16; #100;
A = 8'h60; B = 8'h17; #100;
A = 8'h60; B = 8'h18; #100;
A = 8'h60; B = 8'h19; #100;
A = 8'h60; B = 8'h1A; #100;
A = 8'h60; B = 8'h1B; #100;
A = 8'h60; B = 8'h1C; #100;
A = 8'h60; B = 8'h1D; #100;
A = 8'h60; B = 8'h1E; #100;
A = 8'h60; B = 8'h1F; #100;
A = 8'h60; B = 8'h20; #100;
A = 8'h60; B = 8'h21; #100;
A = 8'h60; B = 8'h22; #100;
A = 8'h60; B = 8'h23; #100;
A = 8'h60; B = 8'h24; #100;
A = 8'h60; B = 8'h25; #100;
A = 8'h60; B = 8'h26; #100;
A = 8'h60; B = 8'h27; #100;
A = 8'h60; B = 8'h28; #100;
A = 8'h60; B = 8'h29; #100;
A = 8'h60; B = 8'h2A; #100;
A = 8'h60; B = 8'h2B; #100;
A = 8'h60; B = 8'h2C; #100;
A = 8'h60; B = 8'h2D; #100;
A = 8'h60; B = 8'h2E; #100;
A = 8'h60; B = 8'h2F; #100;
A = 8'h60; B = 8'h30; #100;
A = 8'h60; B = 8'h31; #100;
A = 8'h60; B = 8'h32; #100;
A = 8'h60; B = 8'h33; #100;
A = 8'h60; B = 8'h34; #100;
A = 8'h60; B = 8'h35; #100;
A = 8'h60; B = 8'h36; #100;
A = 8'h60; B = 8'h37; #100;
A = 8'h60; B = 8'h38; #100;
A = 8'h60; B = 8'h39; #100;
A = 8'h60; B = 8'h3A; #100;
A = 8'h60; B = 8'h3B; #100;
A = 8'h60; B = 8'h3C; #100;
A = 8'h60; B = 8'h3D; #100;
A = 8'h60; B = 8'h3E; #100;
A = 8'h60; B = 8'h3F; #100;
A = 8'h60; B = 8'h40; #100;
A = 8'h60; B = 8'h41; #100;
A = 8'h60; B = 8'h42; #100;
A = 8'h60; B = 8'h43; #100;
A = 8'h60; B = 8'h44; #100;
A = 8'h60; B = 8'h45; #100;
A = 8'h60; B = 8'h46; #100;
A = 8'h60; B = 8'h47; #100;
A = 8'h60; B = 8'h48; #100;
A = 8'h60; B = 8'h49; #100;
A = 8'h60; B = 8'h4A; #100;
A = 8'h60; B = 8'h4B; #100;
A = 8'h60; B = 8'h4C; #100;
A = 8'h60; B = 8'h4D; #100;
A = 8'h60; B = 8'h4E; #100;
A = 8'h60; B = 8'h4F; #100;
A = 8'h60; B = 8'h50; #100;
A = 8'h60; B = 8'h51; #100;
A = 8'h60; B = 8'h52; #100;
A = 8'h60; B = 8'h53; #100;
A = 8'h60; B = 8'h54; #100;
A = 8'h60; B = 8'h55; #100;
A = 8'h60; B = 8'h56; #100;
A = 8'h60; B = 8'h57; #100;
A = 8'h60; B = 8'h58; #100;
A = 8'h60; B = 8'h59; #100;
A = 8'h60; B = 8'h5A; #100;
A = 8'h60; B = 8'h5B; #100;
A = 8'h60; B = 8'h5C; #100;
A = 8'h60; B = 8'h5D; #100;
A = 8'h60; B = 8'h5E; #100;
A = 8'h60; B = 8'h5F; #100;
A = 8'h60; B = 8'h60; #100;
A = 8'h60; B = 8'h61; #100;
A = 8'h60; B = 8'h62; #100;
A = 8'h60; B = 8'h63; #100;
A = 8'h60; B = 8'h64; #100;
A = 8'h60; B = 8'h65; #100;
A = 8'h60; B = 8'h66; #100;
A = 8'h60; B = 8'h67; #100;
A = 8'h60; B = 8'h68; #100;
A = 8'h60; B = 8'h69; #100;
A = 8'h60; B = 8'h6A; #100;
A = 8'h60; B = 8'h6B; #100;
A = 8'h60; B = 8'h6C; #100;
A = 8'h60; B = 8'h6D; #100;
A = 8'h60; B = 8'h6E; #100;
A = 8'h60; B = 8'h6F; #100;
A = 8'h60; B = 8'h70; #100;
A = 8'h60; B = 8'h71; #100;
A = 8'h60; B = 8'h72; #100;
A = 8'h60; B = 8'h73; #100;
A = 8'h60; B = 8'h74; #100;
A = 8'h60; B = 8'h75; #100;
A = 8'h60; B = 8'h76; #100;
A = 8'h60; B = 8'h77; #100;
A = 8'h60; B = 8'h78; #100;
A = 8'h60; B = 8'h79; #100;
A = 8'h60; B = 8'h7A; #100;
A = 8'h60; B = 8'h7B; #100;
A = 8'h60; B = 8'h7C; #100;
A = 8'h60; B = 8'h7D; #100;
A = 8'h60; B = 8'h7E; #100;
A = 8'h60; B = 8'h7F; #100;
A = 8'h60; B = 8'h80; #100;
A = 8'h60; B = 8'h81; #100;
A = 8'h60; B = 8'h82; #100;
A = 8'h60; B = 8'h83; #100;
A = 8'h60; B = 8'h84; #100;
A = 8'h60; B = 8'h85; #100;
A = 8'h60; B = 8'h86; #100;
A = 8'h60; B = 8'h87; #100;
A = 8'h60; B = 8'h88; #100;
A = 8'h60; B = 8'h89; #100;
A = 8'h60; B = 8'h8A; #100;
A = 8'h60; B = 8'h8B; #100;
A = 8'h60; B = 8'h8C; #100;
A = 8'h60; B = 8'h8D; #100;
A = 8'h60; B = 8'h8E; #100;
A = 8'h60; B = 8'h8F; #100;
A = 8'h60; B = 8'h90; #100;
A = 8'h60; B = 8'h91; #100;
A = 8'h60; B = 8'h92; #100;
A = 8'h60; B = 8'h93; #100;
A = 8'h60; B = 8'h94; #100;
A = 8'h60; B = 8'h95; #100;
A = 8'h60; B = 8'h96; #100;
A = 8'h60; B = 8'h97; #100;
A = 8'h60; B = 8'h98; #100;
A = 8'h60; B = 8'h99; #100;
A = 8'h60; B = 8'h9A; #100;
A = 8'h60; B = 8'h9B; #100;
A = 8'h60; B = 8'h9C; #100;
A = 8'h60; B = 8'h9D; #100;
A = 8'h60; B = 8'h9E; #100;
A = 8'h60; B = 8'h9F; #100;
A = 8'h60; B = 8'hA0; #100;
A = 8'h60; B = 8'hA1; #100;
A = 8'h60; B = 8'hA2; #100;
A = 8'h60; B = 8'hA3; #100;
A = 8'h60; B = 8'hA4; #100;
A = 8'h60; B = 8'hA5; #100;
A = 8'h60; B = 8'hA6; #100;
A = 8'h60; B = 8'hA7; #100;
A = 8'h60; B = 8'hA8; #100;
A = 8'h60; B = 8'hA9; #100;
A = 8'h60; B = 8'hAA; #100;
A = 8'h60; B = 8'hAB; #100;
A = 8'h60; B = 8'hAC; #100;
A = 8'h60; B = 8'hAD; #100;
A = 8'h60; B = 8'hAE; #100;
A = 8'h60; B = 8'hAF; #100;
A = 8'h60; B = 8'hB0; #100;
A = 8'h60; B = 8'hB1; #100;
A = 8'h60; B = 8'hB2; #100;
A = 8'h60; B = 8'hB3; #100;
A = 8'h60; B = 8'hB4; #100;
A = 8'h60; B = 8'hB5; #100;
A = 8'h60; B = 8'hB6; #100;
A = 8'h60; B = 8'hB7; #100;
A = 8'h60; B = 8'hB8; #100;
A = 8'h60; B = 8'hB9; #100;
A = 8'h60; B = 8'hBA; #100;
A = 8'h60; B = 8'hBB; #100;
A = 8'h60; B = 8'hBC; #100;
A = 8'h60; B = 8'hBD; #100;
A = 8'h60; B = 8'hBE; #100;
A = 8'h60; B = 8'hBF; #100;
A = 8'h60; B = 8'hC0; #100;
A = 8'h60; B = 8'hC1; #100;
A = 8'h60; B = 8'hC2; #100;
A = 8'h60; B = 8'hC3; #100;
A = 8'h60; B = 8'hC4; #100;
A = 8'h60; B = 8'hC5; #100;
A = 8'h60; B = 8'hC6; #100;
A = 8'h60; B = 8'hC7; #100;
A = 8'h60; B = 8'hC8; #100;
A = 8'h60; B = 8'hC9; #100;
A = 8'h60; B = 8'hCA; #100;
A = 8'h60; B = 8'hCB; #100;
A = 8'h60; B = 8'hCC; #100;
A = 8'h60; B = 8'hCD; #100;
A = 8'h60; B = 8'hCE; #100;
A = 8'h60; B = 8'hCF; #100;
A = 8'h60; B = 8'hD0; #100;
A = 8'h60; B = 8'hD1; #100;
A = 8'h60; B = 8'hD2; #100;
A = 8'h60; B = 8'hD3; #100;
A = 8'h60; B = 8'hD4; #100;
A = 8'h60; B = 8'hD5; #100;
A = 8'h60; B = 8'hD6; #100;
A = 8'h60; B = 8'hD7; #100;
A = 8'h60; B = 8'hD8; #100;
A = 8'h60; B = 8'hD9; #100;
A = 8'h60; B = 8'hDA; #100;
A = 8'h60; B = 8'hDB; #100;
A = 8'h60; B = 8'hDC; #100;
A = 8'h60; B = 8'hDD; #100;
A = 8'h60; B = 8'hDE; #100;
A = 8'h60; B = 8'hDF; #100;
A = 8'h60; B = 8'hE0; #100;
A = 8'h60; B = 8'hE1; #100;
A = 8'h60; B = 8'hE2; #100;
A = 8'h60; B = 8'hE3; #100;
A = 8'h60; B = 8'hE4; #100;
A = 8'h60; B = 8'hE5; #100;
A = 8'h60; B = 8'hE6; #100;
A = 8'h60; B = 8'hE7; #100;
A = 8'h60; B = 8'hE8; #100;
A = 8'h60; B = 8'hE9; #100;
A = 8'h60; B = 8'hEA; #100;
A = 8'h60; B = 8'hEB; #100;
A = 8'h60; B = 8'hEC; #100;
A = 8'h60; B = 8'hED; #100;
A = 8'h60; B = 8'hEE; #100;
A = 8'h60; B = 8'hEF; #100;
A = 8'h60; B = 8'hF0; #100;
A = 8'h60; B = 8'hF1; #100;
A = 8'h60; B = 8'hF2; #100;
A = 8'h60; B = 8'hF3; #100;
A = 8'h60; B = 8'hF4; #100;
A = 8'h60; B = 8'hF5; #100;
A = 8'h60; B = 8'hF6; #100;
A = 8'h60; B = 8'hF7; #100;
A = 8'h60; B = 8'hF8; #100;
A = 8'h60; B = 8'hF9; #100;
A = 8'h60; B = 8'hFA; #100;
A = 8'h60; B = 8'hFB; #100;
A = 8'h60; B = 8'hFC; #100;
A = 8'h60; B = 8'hFD; #100;
A = 8'h60; B = 8'hFE; #100;
A = 8'h60; B = 8'hFF; #100;
A = 8'h61; B = 8'h0; #100;
A = 8'h61; B = 8'h1; #100;
A = 8'h61; B = 8'h2; #100;
A = 8'h61; B = 8'h3; #100;
A = 8'h61; B = 8'h4; #100;
A = 8'h61; B = 8'h5; #100;
A = 8'h61; B = 8'h6; #100;
A = 8'h61; B = 8'h7; #100;
A = 8'h61; B = 8'h8; #100;
A = 8'h61; B = 8'h9; #100;
A = 8'h61; B = 8'hA; #100;
A = 8'h61; B = 8'hB; #100;
A = 8'h61; B = 8'hC; #100;
A = 8'h61; B = 8'hD; #100;
A = 8'h61; B = 8'hE; #100;
A = 8'h61; B = 8'hF; #100;
A = 8'h61; B = 8'h10; #100;
A = 8'h61; B = 8'h11; #100;
A = 8'h61; B = 8'h12; #100;
A = 8'h61; B = 8'h13; #100;
A = 8'h61; B = 8'h14; #100;
A = 8'h61; B = 8'h15; #100;
A = 8'h61; B = 8'h16; #100;
A = 8'h61; B = 8'h17; #100;
A = 8'h61; B = 8'h18; #100;
A = 8'h61; B = 8'h19; #100;
A = 8'h61; B = 8'h1A; #100;
A = 8'h61; B = 8'h1B; #100;
A = 8'h61; B = 8'h1C; #100;
A = 8'h61; B = 8'h1D; #100;
A = 8'h61; B = 8'h1E; #100;
A = 8'h61; B = 8'h1F; #100;
A = 8'h61; B = 8'h20; #100;
A = 8'h61; B = 8'h21; #100;
A = 8'h61; B = 8'h22; #100;
A = 8'h61; B = 8'h23; #100;
A = 8'h61; B = 8'h24; #100;
A = 8'h61; B = 8'h25; #100;
A = 8'h61; B = 8'h26; #100;
A = 8'h61; B = 8'h27; #100;
A = 8'h61; B = 8'h28; #100;
A = 8'h61; B = 8'h29; #100;
A = 8'h61; B = 8'h2A; #100;
A = 8'h61; B = 8'h2B; #100;
A = 8'h61; B = 8'h2C; #100;
A = 8'h61; B = 8'h2D; #100;
A = 8'h61; B = 8'h2E; #100;
A = 8'h61; B = 8'h2F; #100;
A = 8'h61; B = 8'h30; #100;
A = 8'h61; B = 8'h31; #100;
A = 8'h61; B = 8'h32; #100;
A = 8'h61; B = 8'h33; #100;
A = 8'h61; B = 8'h34; #100;
A = 8'h61; B = 8'h35; #100;
A = 8'h61; B = 8'h36; #100;
A = 8'h61; B = 8'h37; #100;
A = 8'h61; B = 8'h38; #100;
A = 8'h61; B = 8'h39; #100;
A = 8'h61; B = 8'h3A; #100;
A = 8'h61; B = 8'h3B; #100;
A = 8'h61; B = 8'h3C; #100;
A = 8'h61; B = 8'h3D; #100;
A = 8'h61; B = 8'h3E; #100;
A = 8'h61; B = 8'h3F; #100;
A = 8'h61; B = 8'h40; #100;
A = 8'h61; B = 8'h41; #100;
A = 8'h61; B = 8'h42; #100;
A = 8'h61; B = 8'h43; #100;
A = 8'h61; B = 8'h44; #100;
A = 8'h61; B = 8'h45; #100;
A = 8'h61; B = 8'h46; #100;
A = 8'h61; B = 8'h47; #100;
A = 8'h61; B = 8'h48; #100;
A = 8'h61; B = 8'h49; #100;
A = 8'h61; B = 8'h4A; #100;
A = 8'h61; B = 8'h4B; #100;
A = 8'h61; B = 8'h4C; #100;
A = 8'h61; B = 8'h4D; #100;
A = 8'h61; B = 8'h4E; #100;
A = 8'h61; B = 8'h4F; #100;
A = 8'h61; B = 8'h50; #100;
A = 8'h61; B = 8'h51; #100;
A = 8'h61; B = 8'h52; #100;
A = 8'h61; B = 8'h53; #100;
A = 8'h61; B = 8'h54; #100;
A = 8'h61; B = 8'h55; #100;
A = 8'h61; B = 8'h56; #100;
A = 8'h61; B = 8'h57; #100;
A = 8'h61; B = 8'h58; #100;
A = 8'h61; B = 8'h59; #100;
A = 8'h61; B = 8'h5A; #100;
A = 8'h61; B = 8'h5B; #100;
A = 8'h61; B = 8'h5C; #100;
A = 8'h61; B = 8'h5D; #100;
A = 8'h61; B = 8'h5E; #100;
A = 8'h61; B = 8'h5F; #100;
A = 8'h61; B = 8'h60; #100;
A = 8'h61; B = 8'h61; #100;
A = 8'h61; B = 8'h62; #100;
A = 8'h61; B = 8'h63; #100;
A = 8'h61; B = 8'h64; #100;
A = 8'h61; B = 8'h65; #100;
A = 8'h61; B = 8'h66; #100;
A = 8'h61; B = 8'h67; #100;
A = 8'h61; B = 8'h68; #100;
A = 8'h61; B = 8'h69; #100;
A = 8'h61; B = 8'h6A; #100;
A = 8'h61; B = 8'h6B; #100;
A = 8'h61; B = 8'h6C; #100;
A = 8'h61; B = 8'h6D; #100;
A = 8'h61; B = 8'h6E; #100;
A = 8'h61; B = 8'h6F; #100;
A = 8'h61; B = 8'h70; #100;
A = 8'h61; B = 8'h71; #100;
A = 8'h61; B = 8'h72; #100;
A = 8'h61; B = 8'h73; #100;
A = 8'h61; B = 8'h74; #100;
A = 8'h61; B = 8'h75; #100;
A = 8'h61; B = 8'h76; #100;
A = 8'h61; B = 8'h77; #100;
A = 8'h61; B = 8'h78; #100;
A = 8'h61; B = 8'h79; #100;
A = 8'h61; B = 8'h7A; #100;
A = 8'h61; B = 8'h7B; #100;
A = 8'h61; B = 8'h7C; #100;
A = 8'h61; B = 8'h7D; #100;
A = 8'h61; B = 8'h7E; #100;
A = 8'h61; B = 8'h7F; #100;
A = 8'h61; B = 8'h80; #100;
A = 8'h61; B = 8'h81; #100;
A = 8'h61; B = 8'h82; #100;
A = 8'h61; B = 8'h83; #100;
A = 8'h61; B = 8'h84; #100;
A = 8'h61; B = 8'h85; #100;
A = 8'h61; B = 8'h86; #100;
A = 8'h61; B = 8'h87; #100;
A = 8'h61; B = 8'h88; #100;
A = 8'h61; B = 8'h89; #100;
A = 8'h61; B = 8'h8A; #100;
A = 8'h61; B = 8'h8B; #100;
A = 8'h61; B = 8'h8C; #100;
A = 8'h61; B = 8'h8D; #100;
A = 8'h61; B = 8'h8E; #100;
A = 8'h61; B = 8'h8F; #100;
A = 8'h61; B = 8'h90; #100;
A = 8'h61; B = 8'h91; #100;
A = 8'h61; B = 8'h92; #100;
A = 8'h61; B = 8'h93; #100;
A = 8'h61; B = 8'h94; #100;
A = 8'h61; B = 8'h95; #100;
A = 8'h61; B = 8'h96; #100;
A = 8'h61; B = 8'h97; #100;
A = 8'h61; B = 8'h98; #100;
A = 8'h61; B = 8'h99; #100;
A = 8'h61; B = 8'h9A; #100;
A = 8'h61; B = 8'h9B; #100;
A = 8'h61; B = 8'h9C; #100;
A = 8'h61; B = 8'h9D; #100;
A = 8'h61; B = 8'h9E; #100;
A = 8'h61; B = 8'h9F; #100;
A = 8'h61; B = 8'hA0; #100;
A = 8'h61; B = 8'hA1; #100;
A = 8'h61; B = 8'hA2; #100;
A = 8'h61; B = 8'hA3; #100;
A = 8'h61; B = 8'hA4; #100;
A = 8'h61; B = 8'hA5; #100;
A = 8'h61; B = 8'hA6; #100;
A = 8'h61; B = 8'hA7; #100;
A = 8'h61; B = 8'hA8; #100;
A = 8'h61; B = 8'hA9; #100;
A = 8'h61; B = 8'hAA; #100;
A = 8'h61; B = 8'hAB; #100;
A = 8'h61; B = 8'hAC; #100;
A = 8'h61; B = 8'hAD; #100;
A = 8'h61; B = 8'hAE; #100;
A = 8'h61; B = 8'hAF; #100;
A = 8'h61; B = 8'hB0; #100;
A = 8'h61; B = 8'hB1; #100;
A = 8'h61; B = 8'hB2; #100;
A = 8'h61; B = 8'hB3; #100;
A = 8'h61; B = 8'hB4; #100;
A = 8'h61; B = 8'hB5; #100;
A = 8'h61; B = 8'hB6; #100;
A = 8'h61; B = 8'hB7; #100;
A = 8'h61; B = 8'hB8; #100;
A = 8'h61; B = 8'hB9; #100;
A = 8'h61; B = 8'hBA; #100;
A = 8'h61; B = 8'hBB; #100;
A = 8'h61; B = 8'hBC; #100;
A = 8'h61; B = 8'hBD; #100;
A = 8'h61; B = 8'hBE; #100;
A = 8'h61; B = 8'hBF; #100;
A = 8'h61; B = 8'hC0; #100;
A = 8'h61; B = 8'hC1; #100;
A = 8'h61; B = 8'hC2; #100;
A = 8'h61; B = 8'hC3; #100;
A = 8'h61; B = 8'hC4; #100;
A = 8'h61; B = 8'hC5; #100;
A = 8'h61; B = 8'hC6; #100;
A = 8'h61; B = 8'hC7; #100;
A = 8'h61; B = 8'hC8; #100;
A = 8'h61; B = 8'hC9; #100;
A = 8'h61; B = 8'hCA; #100;
A = 8'h61; B = 8'hCB; #100;
A = 8'h61; B = 8'hCC; #100;
A = 8'h61; B = 8'hCD; #100;
A = 8'h61; B = 8'hCE; #100;
A = 8'h61; B = 8'hCF; #100;
A = 8'h61; B = 8'hD0; #100;
A = 8'h61; B = 8'hD1; #100;
A = 8'h61; B = 8'hD2; #100;
A = 8'h61; B = 8'hD3; #100;
A = 8'h61; B = 8'hD4; #100;
A = 8'h61; B = 8'hD5; #100;
A = 8'h61; B = 8'hD6; #100;
A = 8'h61; B = 8'hD7; #100;
A = 8'h61; B = 8'hD8; #100;
A = 8'h61; B = 8'hD9; #100;
A = 8'h61; B = 8'hDA; #100;
A = 8'h61; B = 8'hDB; #100;
A = 8'h61; B = 8'hDC; #100;
A = 8'h61; B = 8'hDD; #100;
A = 8'h61; B = 8'hDE; #100;
A = 8'h61; B = 8'hDF; #100;
A = 8'h61; B = 8'hE0; #100;
A = 8'h61; B = 8'hE1; #100;
A = 8'h61; B = 8'hE2; #100;
A = 8'h61; B = 8'hE3; #100;
A = 8'h61; B = 8'hE4; #100;
A = 8'h61; B = 8'hE5; #100;
A = 8'h61; B = 8'hE6; #100;
A = 8'h61; B = 8'hE7; #100;
A = 8'h61; B = 8'hE8; #100;
A = 8'h61; B = 8'hE9; #100;
A = 8'h61; B = 8'hEA; #100;
A = 8'h61; B = 8'hEB; #100;
A = 8'h61; B = 8'hEC; #100;
A = 8'h61; B = 8'hED; #100;
A = 8'h61; B = 8'hEE; #100;
A = 8'h61; B = 8'hEF; #100;
A = 8'h61; B = 8'hF0; #100;
A = 8'h61; B = 8'hF1; #100;
A = 8'h61; B = 8'hF2; #100;
A = 8'h61; B = 8'hF3; #100;
A = 8'h61; B = 8'hF4; #100;
A = 8'h61; B = 8'hF5; #100;
A = 8'h61; B = 8'hF6; #100;
A = 8'h61; B = 8'hF7; #100;
A = 8'h61; B = 8'hF8; #100;
A = 8'h61; B = 8'hF9; #100;
A = 8'h61; B = 8'hFA; #100;
A = 8'h61; B = 8'hFB; #100;
A = 8'h61; B = 8'hFC; #100;
A = 8'h61; B = 8'hFD; #100;
A = 8'h61; B = 8'hFE; #100;
A = 8'h61; B = 8'hFF; #100;
A = 8'h62; B = 8'h0; #100;
A = 8'h62; B = 8'h1; #100;
A = 8'h62; B = 8'h2; #100;
A = 8'h62; B = 8'h3; #100;
A = 8'h62; B = 8'h4; #100;
A = 8'h62; B = 8'h5; #100;
A = 8'h62; B = 8'h6; #100;
A = 8'h62; B = 8'h7; #100;
A = 8'h62; B = 8'h8; #100;
A = 8'h62; B = 8'h9; #100;
A = 8'h62; B = 8'hA; #100;
A = 8'h62; B = 8'hB; #100;
A = 8'h62; B = 8'hC; #100;
A = 8'h62; B = 8'hD; #100;
A = 8'h62; B = 8'hE; #100;
A = 8'h62; B = 8'hF; #100;
A = 8'h62; B = 8'h10; #100;
A = 8'h62; B = 8'h11; #100;
A = 8'h62; B = 8'h12; #100;
A = 8'h62; B = 8'h13; #100;
A = 8'h62; B = 8'h14; #100;
A = 8'h62; B = 8'h15; #100;
A = 8'h62; B = 8'h16; #100;
A = 8'h62; B = 8'h17; #100;
A = 8'h62; B = 8'h18; #100;
A = 8'h62; B = 8'h19; #100;
A = 8'h62; B = 8'h1A; #100;
A = 8'h62; B = 8'h1B; #100;
A = 8'h62; B = 8'h1C; #100;
A = 8'h62; B = 8'h1D; #100;
A = 8'h62; B = 8'h1E; #100;
A = 8'h62; B = 8'h1F; #100;
A = 8'h62; B = 8'h20; #100;
A = 8'h62; B = 8'h21; #100;
A = 8'h62; B = 8'h22; #100;
A = 8'h62; B = 8'h23; #100;
A = 8'h62; B = 8'h24; #100;
A = 8'h62; B = 8'h25; #100;
A = 8'h62; B = 8'h26; #100;
A = 8'h62; B = 8'h27; #100;
A = 8'h62; B = 8'h28; #100;
A = 8'h62; B = 8'h29; #100;
A = 8'h62; B = 8'h2A; #100;
A = 8'h62; B = 8'h2B; #100;
A = 8'h62; B = 8'h2C; #100;
A = 8'h62; B = 8'h2D; #100;
A = 8'h62; B = 8'h2E; #100;
A = 8'h62; B = 8'h2F; #100;
A = 8'h62; B = 8'h30; #100;
A = 8'h62; B = 8'h31; #100;
A = 8'h62; B = 8'h32; #100;
A = 8'h62; B = 8'h33; #100;
A = 8'h62; B = 8'h34; #100;
A = 8'h62; B = 8'h35; #100;
A = 8'h62; B = 8'h36; #100;
A = 8'h62; B = 8'h37; #100;
A = 8'h62; B = 8'h38; #100;
A = 8'h62; B = 8'h39; #100;
A = 8'h62; B = 8'h3A; #100;
A = 8'h62; B = 8'h3B; #100;
A = 8'h62; B = 8'h3C; #100;
A = 8'h62; B = 8'h3D; #100;
A = 8'h62; B = 8'h3E; #100;
A = 8'h62; B = 8'h3F; #100;
A = 8'h62; B = 8'h40; #100;
A = 8'h62; B = 8'h41; #100;
A = 8'h62; B = 8'h42; #100;
A = 8'h62; B = 8'h43; #100;
A = 8'h62; B = 8'h44; #100;
A = 8'h62; B = 8'h45; #100;
A = 8'h62; B = 8'h46; #100;
A = 8'h62; B = 8'h47; #100;
A = 8'h62; B = 8'h48; #100;
A = 8'h62; B = 8'h49; #100;
A = 8'h62; B = 8'h4A; #100;
A = 8'h62; B = 8'h4B; #100;
A = 8'h62; B = 8'h4C; #100;
A = 8'h62; B = 8'h4D; #100;
A = 8'h62; B = 8'h4E; #100;
A = 8'h62; B = 8'h4F; #100;
A = 8'h62; B = 8'h50; #100;
A = 8'h62; B = 8'h51; #100;
A = 8'h62; B = 8'h52; #100;
A = 8'h62; B = 8'h53; #100;
A = 8'h62; B = 8'h54; #100;
A = 8'h62; B = 8'h55; #100;
A = 8'h62; B = 8'h56; #100;
A = 8'h62; B = 8'h57; #100;
A = 8'h62; B = 8'h58; #100;
A = 8'h62; B = 8'h59; #100;
A = 8'h62; B = 8'h5A; #100;
A = 8'h62; B = 8'h5B; #100;
A = 8'h62; B = 8'h5C; #100;
A = 8'h62; B = 8'h5D; #100;
A = 8'h62; B = 8'h5E; #100;
A = 8'h62; B = 8'h5F; #100;
A = 8'h62; B = 8'h60; #100;
A = 8'h62; B = 8'h61; #100;
A = 8'h62; B = 8'h62; #100;
A = 8'h62; B = 8'h63; #100;
A = 8'h62; B = 8'h64; #100;
A = 8'h62; B = 8'h65; #100;
A = 8'h62; B = 8'h66; #100;
A = 8'h62; B = 8'h67; #100;
A = 8'h62; B = 8'h68; #100;
A = 8'h62; B = 8'h69; #100;
A = 8'h62; B = 8'h6A; #100;
A = 8'h62; B = 8'h6B; #100;
A = 8'h62; B = 8'h6C; #100;
A = 8'h62; B = 8'h6D; #100;
A = 8'h62; B = 8'h6E; #100;
A = 8'h62; B = 8'h6F; #100;
A = 8'h62; B = 8'h70; #100;
A = 8'h62; B = 8'h71; #100;
A = 8'h62; B = 8'h72; #100;
A = 8'h62; B = 8'h73; #100;
A = 8'h62; B = 8'h74; #100;
A = 8'h62; B = 8'h75; #100;
A = 8'h62; B = 8'h76; #100;
A = 8'h62; B = 8'h77; #100;
A = 8'h62; B = 8'h78; #100;
A = 8'h62; B = 8'h79; #100;
A = 8'h62; B = 8'h7A; #100;
A = 8'h62; B = 8'h7B; #100;
A = 8'h62; B = 8'h7C; #100;
A = 8'h62; B = 8'h7D; #100;
A = 8'h62; B = 8'h7E; #100;
A = 8'h62; B = 8'h7F; #100;
A = 8'h62; B = 8'h80; #100;
A = 8'h62; B = 8'h81; #100;
A = 8'h62; B = 8'h82; #100;
A = 8'h62; B = 8'h83; #100;
A = 8'h62; B = 8'h84; #100;
A = 8'h62; B = 8'h85; #100;
A = 8'h62; B = 8'h86; #100;
A = 8'h62; B = 8'h87; #100;
A = 8'h62; B = 8'h88; #100;
A = 8'h62; B = 8'h89; #100;
A = 8'h62; B = 8'h8A; #100;
A = 8'h62; B = 8'h8B; #100;
A = 8'h62; B = 8'h8C; #100;
A = 8'h62; B = 8'h8D; #100;
A = 8'h62; B = 8'h8E; #100;
A = 8'h62; B = 8'h8F; #100;
A = 8'h62; B = 8'h90; #100;
A = 8'h62; B = 8'h91; #100;
A = 8'h62; B = 8'h92; #100;
A = 8'h62; B = 8'h93; #100;
A = 8'h62; B = 8'h94; #100;
A = 8'h62; B = 8'h95; #100;
A = 8'h62; B = 8'h96; #100;
A = 8'h62; B = 8'h97; #100;
A = 8'h62; B = 8'h98; #100;
A = 8'h62; B = 8'h99; #100;
A = 8'h62; B = 8'h9A; #100;
A = 8'h62; B = 8'h9B; #100;
A = 8'h62; B = 8'h9C; #100;
A = 8'h62; B = 8'h9D; #100;
A = 8'h62; B = 8'h9E; #100;
A = 8'h62; B = 8'h9F; #100;
A = 8'h62; B = 8'hA0; #100;
A = 8'h62; B = 8'hA1; #100;
A = 8'h62; B = 8'hA2; #100;
A = 8'h62; B = 8'hA3; #100;
A = 8'h62; B = 8'hA4; #100;
A = 8'h62; B = 8'hA5; #100;
A = 8'h62; B = 8'hA6; #100;
A = 8'h62; B = 8'hA7; #100;
A = 8'h62; B = 8'hA8; #100;
A = 8'h62; B = 8'hA9; #100;
A = 8'h62; B = 8'hAA; #100;
A = 8'h62; B = 8'hAB; #100;
A = 8'h62; B = 8'hAC; #100;
A = 8'h62; B = 8'hAD; #100;
A = 8'h62; B = 8'hAE; #100;
A = 8'h62; B = 8'hAF; #100;
A = 8'h62; B = 8'hB0; #100;
A = 8'h62; B = 8'hB1; #100;
A = 8'h62; B = 8'hB2; #100;
A = 8'h62; B = 8'hB3; #100;
A = 8'h62; B = 8'hB4; #100;
A = 8'h62; B = 8'hB5; #100;
A = 8'h62; B = 8'hB6; #100;
A = 8'h62; B = 8'hB7; #100;
A = 8'h62; B = 8'hB8; #100;
A = 8'h62; B = 8'hB9; #100;
A = 8'h62; B = 8'hBA; #100;
A = 8'h62; B = 8'hBB; #100;
A = 8'h62; B = 8'hBC; #100;
A = 8'h62; B = 8'hBD; #100;
A = 8'h62; B = 8'hBE; #100;
A = 8'h62; B = 8'hBF; #100;
A = 8'h62; B = 8'hC0; #100;
A = 8'h62; B = 8'hC1; #100;
A = 8'h62; B = 8'hC2; #100;
A = 8'h62; B = 8'hC3; #100;
A = 8'h62; B = 8'hC4; #100;
A = 8'h62; B = 8'hC5; #100;
A = 8'h62; B = 8'hC6; #100;
A = 8'h62; B = 8'hC7; #100;
A = 8'h62; B = 8'hC8; #100;
A = 8'h62; B = 8'hC9; #100;
A = 8'h62; B = 8'hCA; #100;
A = 8'h62; B = 8'hCB; #100;
A = 8'h62; B = 8'hCC; #100;
A = 8'h62; B = 8'hCD; #100;
A = 8'h62; B = 8'hCE; #100;
A = 8'h62; B = 8'hCF; #100;
A = 8'h62; B = 8'hD0; #100;
A = 8'h62; B = 8'hD1; #100;
A = 8'h62; B = 8'hD2; #100;
A = 8'h62; B = 8'hD3; #100;
A = 8'h62; B = 8'hD4; #100;
A = 8'h62; B = 8'hD5; #100;
A = 8'h62; B = 8'hD6; #100;
A = 8'h62; B = 8'hD7; #100;
A = 8'h62; B = 8'hD8; #100;
A = 8'h62; B = 8'hD9; #100;
A = 8'h62; B = 8'hDA; #100;
A = 8'h62; B = 8'hDB; #100;
A = 8'h62; B = 8'hDC; #100;
A = 8'h62; B = 8'hDD; #100;
A = 8'h62; B = 8'hDE; #100;
A = 8'h62; B = 8'hDF; #100;
A = 8'h62; B = 8'hE0; #100;
A = 8'h62; B = 8'hE1; #100;
A = 8'h62; B = 8'hE2; #100;
A = 8'h62; B = 8'hE3; #100;
A = 8'h62; B = 8'hE4; #100;
A = 8'h62; B = 8'hE5; #100;
A = 8'h62; B = 8'hE6; #100;
A = 8'h62; B = 8'hE7; #100;
A = 8'h62; B = 8'hE8; #100;
A = 8'h62; B = 8'hE9; #100;
A = 8'h62; B = 8'hEA; #100;
A = 8'h62; B = 8'hEB; #100;
A = 8'h62; B = 8'hEC; #100;
A = 8'h62; B = 8'hED; #100;
A = 8'h62; B = 8'hEE; #100;
A = 8'h62; B = 8'hEF; #100;
A = 8'h62; B = 8'hF0; #100;
A = 8'h62; B = 8'hF1; #100;
A = 8'h62; B = 8'hF2; #100;
A = 8'h62; B = 8'hF3; #100;
A = 8'h62; B = 8'hF4; #100;
A = 8'h62; B = 8'hF5; #100;
A = 8'h62; B = 8'hF6; #100;
A = 8'h62; B = 8'hF7; #100;
A = 8'h62; B = 8'hF8; #100;
A = 8'h62; B = 8'hF9; #100;
A = 8'h62; B = 8'hFA; #100;
A = 8'h62; B = 8'hFB; #100;
A = 8'h62; B = 8'hFC; #100;
A = 8'h62; B = 8'hFD; #100;
A = 8'h62; B = 8'hFE; #100;
A = 8'h62; B = 8'hFF; #100;
A = 8'h63; B = 8'h0; #100;
A = 8'h63; B = 8'h1; #100;
A = 8'h63; B = 8'h2; #100;
A = 8'h63; B = 8'h3; #100;
A = 8'h63; B = 8'h4; #100;
A = 8'h63; B = 8'h5; #100;
A = 8'h63; B = 8'h6; #100;
A = 8'h63; B = 8'h7; #100;
A = 8'h63; B = 8'h8; #100;
A = 8'h63; B = 8'h9; #100;
A = 8'h63; B = 8'hA; #100;
A = 8'h63; B = 8'hB; #100;
A = 8'h63; B = 8'hC; #100;
A = 8'h63; B = 8'hD; #100;
A = 8'h63; B = 8'hE; #100;
A = 8'h63; B = 8'hF; #100;
A = 8'h63; B = 8'h10; #100;
A = 8'h63; B = 8'h11; #100;
A = 8'h63; B = 8'h12; #100;
A = 8'h63; B = 8'h13; #100;
A = 8'h63; B = 8'h14; #100;
A = 8'h63; B = 8'h15; #100;
A = 8'h63; B = 8'h16; #100;
A = 8'h63; B = 8'h17; #100;
A = 8'h63; B = 8'h18; #100;
A = 8'h63; B = 8'h19; #100;
A = 8'h63; B = 8'h1A; #100;
A = 8'h63; B = 8'h1B; #100;
A = 8'h63; B = 8'h1C; #100;
A = 8'h63; B = 8'h1D; #100;
A = 8'h63; B = 8'h1E; #100;
A = 8'h63; B = 8'h1F; #100;
A = 8'h63; B = 8'h20; #100;
A = 8'h63; B = 8'h21; #100;
A = 8'h63; B = 8'h22; #100;
A = 8'h63; B = 8'h23; #100;
A = 8'h63; B = 8'h24; #100;
A = 8'h63; B = 8'h25; #100;
A = 8'h63; B = 8'h26; #100;
A = 8'h63; B = 8'h27; #100;
A = 8'h63; B = 8'h28; #100;
A = 8'h63; B = 8'h29; #100;
A = 8'h63; B = 8'h2A; #100;
A = 8'h63; B = 8'h2B; #100;
A = 8'h63; B = 8'h2C; #100;
A = 8'h63; B = 8'h2D; #100;
A = 8'h63; B = 8'h2E; #100;
A = 8'h63; B = 8'h2F; #100;
A = 8'h63; B = 8'h30; #100;
A = 8'h63; B = 8'h31; #100;
A = 8'h63; B = 8'h32; #100;
A = 8'h63; B = 8'h33; #100;
A = 8'h63; B = 8'h34; #100;
A = 8'h63; B = 8'h35; #100;
A = 8'h63; B = 8'h36; #100;
A = 8'h63; B = 8'h37; #100;
A = 8'h63; B = 8'h38; #100;
A = 8'h63; B = 8'h39; #100;
A = 8'h63; B = 8'h3A; #100;
A = 8'h63; B = 8'h3B; #100;
A = 8'h63; B = 8'h3C; #100;
A = 8'h63; B = 8'h3D; #100;
A = 8'h63; B = 8'h3E; #100;
A = 8'h63; B = 8'h3F; #100;
A = 8'h63; B = 8'h40; #100;
A = 8'h63; B = 8'h41; #100;
A = 8'h63; B = 8'h42; #100;
A = 8'h63; B = 8'h43; #100;
A = 8'h63; B = 8'h44; #100;
A = 8'h63; B = 8'h45; #100;
A = 8'h63; B = 8'h46; #100;
A = 8'h63; B = 8'h47; #100;
A = 8'h63; B = 8'h48; #100;
A = 8'h63; B = 8'h49; #100;
A = 8'h63; B = 8'h4A; #100;
A = 8'h63; B = 8'h4B; #100;
A = 8'h63; B = 8'h4C; #100;
A = 8'h63; B = 8'h4D; #100;
A = 8'h63; B = 8'h4E; #100;
A = 8'h63; B = 8'h4F; #100;
A = 8'h63; B = 8'h50; #100;
A = 8'h63; B = 8'h51; #100;
A = 8'h63; B = 8'h52; #100;
A = 8'h63; B = 8'h53; #100;
A = 8'h63; B = 8'h54; #100;
A = 8'h63; B = 8'h55; #100;
A = 8'h63; B = 8'h56; #100;
A = 8'h63; B = 8'h57; #100;
A = 8'h63; B = 8'h58; #100;
A = 8'h63; B = 8'h59; #100;
A = 8'h63; B = 8'h5A; #100;
A = 8'h63; B = 8'h5B; #100;
A = 8'h63; B = 8'h5C; #100;
A = 8'h63; B = 8'h5D; #100;
A = 8'h63; B = 8'h5E; #100;
A = 8'h63; B = 8'h5F; #100;
A = 8'h63; B = 8'h60; #100;
A = 8'h63; B = 8'h61; #100;
A = 8'h63; B = 8'h62; #100;
A = 8'h63; B = 8'h63; #100;
A = 8'h63; B = 8'h64; #100;
A = 8'h63; B = 8'h65; #100;
A = 8'h63; B = 8'h66; #100;
A = 8'h63; B = 8'h67; #100;
A = 8'h63; B = 8'h68; #100;
A = 8'h63; B = 8'h69; #100;
A = 8'h63; B = 8'h6A; #100;
A = 8'h63; B = 8'h6B; #100;
A = 8'h63; B = 8'h6C; #100;
A = 8'h63; B = 8'h6D; #100;
A = 8'h63; B = 8'h6E; #100;
A = 8'h63; B = 8'h6F; #100;
A = 8'h63; B = 8'h70; #100;
A = 8'h63; B = 8'h71; #100;
A = 8'h63; B = 8'h72; #100;
A = 8'h63; B = 8'h73; #100;
A = 8'h63; B = 8'h74; #100;
A = 8'h63; B = 8'h75; #100;
A = 8'h63; B = 8'h76; #100;
A = 8'h63; B = 8'h77; #100;
A = 8'h63; B = 8'h78; #100;
A = 8'h63; B = 8'h79; #100;
A = 8'h63; B = 8'h7A; #100;
A = 8'h63; B = 8'h7B; #100;
A = 8'h63; B = 8'h7C; #100;
A = 8'h63; B = 8'h7D; #100;
A = 8'h63; B = 8'h7E; #100;
A = 8'h63; B = 8'h7F; #100;
A = 8'h63; B = 8'h80; #100;
A = 8'h63; B = 8'h81; #100;
A = 8'h63; B = 8'h82; #100;
A = 8'h63; B = 8'h83; #100;
A = 8'h63; B = 8'h84; #100;
A = 8'h63; B = 8'h85; #100;
A = 8'h63; B = 8'h86; #100;
A = 8'h63; B = 8'h87; #100;
A = 8'h63; B = 8'h88; #100;
A = 8'h63; B = 8'h89; #100;
A = 8'h63; B = 8'h8A; #100;
A = 8'h63; B = 8'h8B; #100;
A = 8'h63; B = 8'h8C; #100;
A = 8'h63; B = 8'h8D; #100;
A = 8'h63; B = 8'h8E; #100;
A = 8'h63; B = 8'h8F; #100;
A = 8'h63; B = 8'h90; #100;
A = 8'h63; B = 8'h91; #100;
A = 8'h63; B = 8'h92; #100;
A = 8'h63; B = 8'h93; #100;
A = 8'h63; B = 8'h94; #100;
A = 8'h63; B = 8'h95; #100;
A = 8'h63; B = 8'h96; #100;
A = 8'h63; B = 8'h97; #100;
A = 8'h63; B = 8'h98; #100;
A = 8'h63; B = 8'h99; #100;
A = 8'h63; B = 8'h9A; #100;
A = 8'h63; B = 8'h9B; #100;
A = 8'h63; B = 8'h9C; #100;
A = 8'h63; B = 8'h9D; #100;
A = 8'h63; B = 8'h9E; #100;
A = 8'h63; B = 8'h9F; #100;
A = 8'h63; B = 8'hA0; #100;
A = 8'h63; B = 8'hA1; #100;
A = 8'h63; B = 8'hA2; #100;
A = 8'h63; B = 8'hA3; #100;
A = 8'h63; B = 8'hA4; #100;
A = 8'h63; B = 8'hA5; #100;
A = 8'h63; B = 8'hA6; #100;
A = 8'h63; B = 8'hA7; #100;
A = 8'h63; B = 8'hA8; #100;
A = 8'h63; B = 8'hA9; #100;
A = 8'h63; B = 8'hAA; #100;
A = 8'h63; B = 8'hAB; #100;
A = 8'h63; B = 8'hAC; #100;
A = 8'h63; B = 8'hAD; #100;
A = 8'h63; B = 8'hAE; #100;
A = 8'h63; B = 8'hAF; #100;
A = 8'h63; B = 8'hB0; #100;
A = 8'h63; B = 8'hB1; #100;
A = 8'h63; B = 8'hB2; #100;
A = 8'h63; B = 8'hB3; #100;
A = 8'h63; B = 8'hB4; #100;
A = 8'h63; B = 8'hB5; #100;
A = 8'h63; B = 8'hB6; #100;
A = 8'h63; B = 8'hB7; #100;
A = 8'h63; B = 8'hB8; #100;
A = 8'h63; B = 8'hB9; #100;
A = 8'h63; B = 8'hBA; #100;
A = 8'h63; B = 8'hBB; #100;
A = 8'h63; B = 8'hBC; #100;
A = 8'h63; B = 8'hBD; #100;
A = 8'h63; B = 8'hBE; #100;
A = 8'h63; B = 8'hBF; #100;
A = 8'h63; B = 8'hC0; #100;
A = 8'h63; B = 8'hC1; #100;
A = 8'h63; B = 8'hC2; #100;
A = 8'h63; B = 8'hC3; #100;
A = 8'h63; B = 8'hC4; #100;
A = 8'h63; B = 8'hC5; #100;
A = 8'h63; B = 8'hC6; #100;
A = 8'h63; B = 8'hC7; #100;
A = 8'h63; B = 8'hC8; #100;
A = 8'h63; B = 8'hC9; #100;
A = 8'h63; B = 8'hCA; #100;
A = 8'h63; B = 8'hCB; #100;
A = 8'h63; B = 8'hCC; #100;
A = 8'h63; B = 8'hCD; #100;
A = 8'h63; B = 8'hCE; #100;
A = 8'h63; B = 8'hCF; #100;
A = 8'h63; B = 8'hD0; #100;
A = 8'h63; B = 8'hD1; #100;
A = 8'h63; B = 8'hD2; #100;
A = 8'h63; B = 8'hD3; #100;
A = 8'h63; B = 8'hD4; #100;
A = 8'h63; B = 8'hD5; #100;
A = 8'h63; B = 8'hD6; #100;
A = 8'h63; B = 8'hD7; #100;
A = 8'h63; B = 8'hD8; #100;
A = 8'h63; B = 8'hD9; #100;
A = 8'h63; B = 8'hDA; #100;
A = 8'h63; B = 8'hDB; #100;
A = 8'h63; B = 8'hDC; #100;
A = 8'h63; B = 8'hDD; #100;
A = 8'h63; B = 8'hDE; #100;
A = 8'h63; B = 8'hDF; #100;
A = 8'h63; B = 8'hE0; #100;
A = 8'h63; B = 8'hE1; #100;
A = 8'h63; B = 8'hE2; #100;
A = 8'h63; B = 8'hE3; #100;
A = 8'h63; B = 8'hE4; #100;
A = 8'h63; B = 8'hE5; #100;
A = 8'h63; B = 8'hE6; #100;
A = 8'h63; B = 8'hE7; #100;
A = 8'h63; B = 8'hE8; #100;
A = 8'h63; B = 8'hE9; #100;
A = 8'h63; B = 8'hEA; #100;
A = 8'h63; B = 8'hEB; #100;
A = 8'h63; B = 8'hEC; #100;
A = 8'h63; B = 8'hED; #100;
A = 8'h63; B = 8'hEE; #100;
A = 8'h63; B = 8'hEF; #100;
A = 8'h63; B = 8'hF0; #100;
A = 8'h63; B = 8'hF1; #100;
A = 8'h63; B = 8'hF2; #100;
A = 8'h63; B = 8'hF3; #100;
A = 8'h63; B = 8'hF4; #100;
A = 8'h63; B = 8'hF5; #100;
A = 8'h63; B = 8'hF6; #100;
A = 8'h63; B = 8'hF7; #100;
A = 8'h63; B = 8'hF8; #100;
A = 8'h63; B = 8'hF9; #100;
A = 8'h63; B = 8'hFA; #100;
A = 8'h63; B = 8'hFB; #100;
A = 8'h63; B = 8'hFC; #100;
A = 8'h63; B = 8'hFD; #100;
A = 8'h63; B = 8'hFE; #100;
A = 8'h63; B = 8'hFF; #100;
A = 8'h64; B = 8'h0; #100;
A = 8'h64; B = 8'h1; #100;
A = 8'h64; B = 8'h2; #100;
A = 8'h64; B = 8'h3; #100;
A = 8'h64; B = 8'h4; #100;
A = 8'h64; B = 8'h5; #100;
A = 8'h64; B = 8'h6; #100;
A = 8'h64; B = 8'h7; #100;
A = 8'h64; B = 8'h8; #100;
A = 8'h64; B = 8'h9; #100;
A = 8'h64; B = 8'hA; #100;
A = 8'h64; B = 8'hB; #100;
A = 8'h64; B = 8'hC; #100;
A = 8'h64; B = 8'hD; #100;
A = 8'h64; B = 8'hE; #100;
A = 8'h64; B = 8'hF; #100;
A = 8'h64; B = 8'h10; #100;
A = 8'h64; B = 8'h11; #100;
A = 8'h64; B = 8'h12; #100;
A = 8'h64; B = 8'h13; #100;
A = 8'h64; B = 8'h14; #100;
A = 8'h64; B = 8'h15; #100;
A = 8'h64; B = 8'h16; #100;
A = 8'h64; B = 8'h17; #100;
A = 8'h64; B = 8'h18; #100;
A = 8'h64; B = 8'h19; #100;
A = 8'h64; B = 8'h1A; #100;
A = 8'h64; B = 8'h1B; #100;
A = 8'h64; B = 8'h1C; #100;
A = 8'h64; B = 8'h1D; #100;
A = 8'h64; B = 8'h1E; #100;
A = 8'h64; B = 8'h1F; #100;
A = 8'h64; B = 8'h20; #100;
A = 8'h64; B = 8'h21; #100;
A = 8'h64; B = 8'h22; #100;
A = 8'h64; B = 8'h23; #100;
A = 8'h64; B = 8'h24; #100;
A = 8'h64; B = 8'h25; #100;
A = 8'h64; B = 8'h26; #100;
A = 8'h64; B = 8'h27; #100;
A = 8'h64; B = 8'h28; #100;
A = 8'h64; B = 8'h29; #100;
A = 8'h64; B = 8'h2A; #100;
A = 8'h64; B = 8'h2B; #100;
A = 8'h64; B = 8'h2C; #100;
A = 8'h64; B = 8'h2D; #100;
A = 8'h64; B = 8'h2E; #100;
A = 8'h64; B = 8'h2F; #100;
A = 8'h64; B = 8'h30; #100;
A = 8'h64; B = 8'h31; #100;
A = 8'h64; B = 8'h32; #100;
A = 8'h64; B = 8'h33; #100;
A = 8'h64; B = 8'h34; #100;
A = 8'h64; B = 8'h35; #100;
A = 8'h64; B = 8'h36; #100;
A = 8'h64; B = 8'h37; #100;
A = 8'h64; B = 8'h38; #100;
A = 8'h64; B = 8'h39; #100;
A = 8'h64; B = 8'h3A; #100;
A = 8'h64; B = 8'h3B; #100;
A = 8'h64; B = 8'h3C; #100;
A = 8'h64; B = 8'h3D; #100;
A = 8'h64; B = 8'h3E; #100;
A = 8'h64; B = 8'h3F; #100;
A = 8'h64; B = 8'h40; #100;
A = 8'h64; B = 8'h41; #100;
A = 8'h64; B = 8'h42; #100;
A = 8'h64; B = 8'h43; #100;
A = 8'h64; B = 8'h44; #100;
A = 8'h64; B = 8'h45; #100;
A = 8'h64; B = 8'h46; #100;
A = 8'h64; B = 8'h47; #100;
A = 8'h64; B = 8'h48; #100;
A = 8'h64; B = 8'h49; #100;
A = 8'h64; B = 8'h4A; #100;
A = 8'h64; B = 8'h4B; #100;
A = 8'h64; B = 8'h4C; #100;
A = 8'h64; B = 8'h4D; #100;
A = 8'h64; B = 8'h4E; #100;
A = 8'h64; B = 8'h4F; #100;
A = 8'h64; B = 8'h50; #100;
A = 8'h64; B = 8'h51; #100;
A = 8'h64; B = 8'h52; #100;
A = 8'h64; B = 8'h53; #100;
A = 8'h64; B = 8'h54; #100;
A = 8'h64; B = 8'h55; #100;
A = 8'h64; B = 8'h56; #100;
A = 8'h64; B = 8'h57; #100;
A = 8'h64; B = 8'h58; #100;
A = 8'h64; B = 8'h59; #100;
A = 8'h64; B = 8'h5A; #100;
A = 8'h64; B = 8'h5B; #100;
A = 8'h64; B = 8'h5C; #100;
A = 8'h64; B = 8'h5D; #100;
A = 8'h64; B = 8'h5E; #100;
A = 8'h64; B = 8'h5F; #100;
A = 8'h64; B = 8'h60; #100;
A = 8'h64; B = 8'h61; #100;
A = 8'h64; B = 8'h62; #100;
A = 8'h64; B = 8'h63; #100;
A = 8'h64; B = 8'h64; #100;
A = 8'h64; B = 8'h65; #100;
A = 8'h64; B = 8'h66; #100;
A = 8'h64; B = 8'h67; #100;
A = 8'h64; B = 8'h68; #100;
A = 8'h64; B = 8'h69; #100;
A = 8'h64; B = 8'h6A; #100;
A = 8'h64; B = 8'h6B; #100;
A = 8'h64; B = 8'h6C; #100;
A = 8'h64; B = 8'h6D; #100;
A = 8'h64; B = 8'h6E; #100;
A = 8'h64; B = 8'h6F; #100;
A = 8'h64; B = 8'h70; #100;
A = 8'h64; B = 8'h71; #100;
A = 8'h64; B = 8'h72; #100;
A = 8'h64; B = 8'h73; #100;
A = 8'h64; B = 8'h74; #100;
A = 8'h64; B = 8'h75; #100;
A = 8'h64; B = 8'h76; #100;
A = 8'h64; B = 8'h77; #100;
A = 8'h64; B = 8'h78; #100;
A = 8'h64; B = 8'h79; #100;
A = 8'h64; B = 8'h7A; #100;
A = 8'h64; B = 8'h7B; #100;
A = 8'h64; B = 8'h7C; #100;
A = 8'h64; B = 8'h7D; #100;
A = 8'h64; B = 8'h7E; #100;
A = 8'h64; B = 8'h7F; #100;
A = 8'h64; B = 8'h80; #100;
A = 8'h64; B = 8'h81; #100;
A = 8'h64; B = 8'h82; #100;
A = 8'h64; B = 8'h83; #100;
A = 8'h64; B = 8'h84; #100;
A = 8'h64; B = 8'h85; #100;
A = 8'h64; B = 8'h86; #100;
A = 8'h64; B = 8'h87; #100;
A = 8'h64; B = 8'h88; #100;
A = 8'h64; B = 8'h89; #100;
A = 8'h64; B = 8'h8A; #100;
A = 8'h64; B = 8'h8B; #100;
A = 8'h64; B = 8'h8C; #100;
A = 8'h64; B = 8'h8D; #100;
A = 8'h64; B = 8'h8E; #100;
A = 8'h64; B = 8'h8F; #100;
A = 8'h64; B = 8'h90; #100;
A = 8'h64; B = 8'h91; #100;
A = 8'h64; B = 8'h92; #100;
A = 8'h64; B = 8'h93; #100;
A = 8'h64; B = 8'h94; #100;
A = 8'h64; B = 8'h95; #100;
A = 8'h64; B = 8'h96; #100;
A = 8'h64; B = 8'h97; #100;
A = 8'h64; B = 8'h98; #100;
A = 8'h64; B = 8'h99; #100;
A = 8'h64; B = 8'h9A; #100;
A = 8'h64; B = 8'h9B; #100;
A = 8'h64; B = 8'h9C; #100;
A = 8'h64; B = 8'h9D; #100;
A = 8'h64; B = 8'h9E; #100;
A = 8'h64; B = 8'h9F; #100;
A = 8'h64; B = 8'hA0; #100;
A = 8'h64; B = 8'hA1; #100;
A = 8'h64; B = 8'hA2; #100;
A = 8'h64; B = 8'hA3; #100;
A = 8'h64; B = 8'hA4; #100;
A = 8'h64; B = 8'hA5; #100;
A = 8'h64; B = 8'hA6; #100;
A = 8'h64; B = 8'hA7; #100;
A = 8'h64; B = 8'hA8; #100;
A = 8'h64; B = 8'hA9; #100;
A = 8'h64; B = 8'hAA; #100;
A = 8'h64; B = 8'hAB; #100;
A = 8'h64; B = 8'hAC; #100;
A = 8'h64; B = 8'hAD; #100;
A = 8'h64; B = 8'hAE; #100;
A = 8'h64; B = 8'hAF; #100;
A = 8'h64; B = 8'hB0; #100;
A = 8'h64; B = 8'hB1; #100;
A = 8'h64; B = 8'hB2; #100;
A = 8'h64; B = 8'hB3; #100;
A = 8'h64; B = 8'hB4; #100;
A = 8'h64; B = 8'hB5; #100;
A = 8'h64; B = 8'hB6; #100;
A = 8'h64; B = 8'hB7; #100;
A = 8'h64; B = 8'hB8; #100;
A = 8'h64; B = 8'hB9; #100;
A = 8'h64; B = 8'hBA; #100;
A = 8'h64; B = 8'hBB; #100;
A = 8'h64; B = 8'hBC; #100;
A = 8'h64; B = 8'hBD; #100;
A = 8'h64; B = 8'hBE; #100;
A = 8'h64; B = 8'hBF; #100;
A = 8'h64; B = 8'hC0; #100;
A = 8'h64; B = 8'hC1; #100;
A = 8'h64; B = 8'hC2; #100;
A = 8'h64; B = 8'hC3; #100;
A = 8'h64; B = 8'hC4; #100;
A = 8'h64; B = 8'hC5; #100;
A = 8'h64; B = 8'hC6; #100;
A = 8'h64; B = 8'hC7; #100;
A = 8'h64; B = 8'hC8; #100;
A = 8'h64; B = 8'hC9; #100;
A = 8'h64; B = 8'hCA; #100;
A = 8'h64; B = 8'hCB; #100;
A = 8'h64; B = 8'hCC; #100;
A = 8'h64; B = 8'hCD; #100;
A = 8'h64; B = 8'hCE; #100;
A = 8'h64; B = 8'hCF; #100;
A = 8'h64; B = 8'hD0; #100;
A = 8'h64; B = 8'hD1; #100;
A = 8'h64; B = 8'hD2; #100;
A = 8'h64; B = 8'hD3; #100;
A = 8'h64; B = 8'hD4; #100;
A = 8'h64; B = 8'hD5; #100;
A = 8'h64; B = 8'hD6; #100;
A = 8'h64; B = 8'hD7; #100;
A = 8'h64; B = 8'hD8; #100;
A = 8'h64; B = 8'hD9; #100;
A = 8'h64; B = 8'hDA; #100;
A = 8'h64; B = 8'hDB; #100;
A = 8'h64; B = 8'hDC; #100;
A = 8'h64; B = 8'hDD; #100;
A = 8'h64; B = 8'hDE; #100;
A = 8'h64; B = 8'hDF; #100;
A = 8'h64; B = 8'hE0; #100;
A = 8'h64; B = 8'hE1; #100;
A = 8'h64; B = 8'hE2; #100;
A = 8'h64; B = 8'hE3; #100;
A = 8'h64; B = 8'hE4; #100;
A = 8'h64; B = 8'hE5; #100;
A = 8'h64; B = 8'hE6; #100;
A = 8'h64; B = 8'hE7; #100;
A = 8'h64; B = 8'hE8; #100;
A = 8'h64; B = 8'hE9; #100;
A = 8'h64; B = 8'hEA; #100;
A = 8'h64; B = 8'hEB; #100;
A = 8'h64; B = 8'hEC; #100;
A = 8'h64; B = 8'hED; #100;
A = 8'h64; B = 8'hEE; #100;
A = 8'h64; B = 8'hEF; #100;
A = 8'h64; B = 8'hF0; #100;
A = 8'h64; B = 8'hF1; #100;
A = 8'h64; B = 8'hF2; #100;
A = 8'h64; B = 8'hF3; #100;
A = 8'h64; B = 8'hF4; #100;
A = 8'h64; B = 8'hF5; #100;
A = 8'h64; B = 8'hF6; #100;
A = 8'h64; B = 8'hF7; #100;
A = 8'h64; B = 8'hF8; #100;
A = 8'h64; B = 8'hF9; #100;
A = 8'h64; B = 8'hFA; #100;
A = 8'h64; B = 8'hFB; #100;
A = 8'h64; B = 8'hFC; #100;
A = 8'h64; B = 8'hFD; #100;
A = 8'h64; B = 8'hFE; #100;
A = 8'h64; B = 8'hFF; #100;
A = 8'h65; B = 8'h0; #100;
A = 8'h65; B = 8'h1; #100;
A = 8'h65; B = 8'h2; #100;
A = 8'h65; B = 8'h3; #100;
A = 8'h65; B = 8'h4; #100;
A = 8'h65; B = 8'h5; #100;
A = 8'h65; B = 8'h6; #100;
A = 8'h65; B = 8'h7; #100;
A = 8'h65; B = 8'h8; #100;
A = 8'h65; B = 8'h9; #100;
A = 8'h65; B = 8'hA; #100;
A = 8'h65; B = 8'hB; #100;
A = 8'h65; B = 8'hC; #100;
A = 8'h65; B = 8'hD; #100;
A = 8'h65; B = 8'hE; #100;
A = 8'h65; B = 8'hF; #100;
A = 8'h65; B = 8'h10; #100;
A = 8'h65; B = 8'h11; #100;
A = 8'h65; B = 8'h12; #100;
A = 8'h65; B = 8'h13; #100;
A = 8'h65; B = 8'h14; #100;
A = 8'h65; B = 8'h15; #100;
A = 8'h65; B = 8'h16; #100;
A = 8'h65; B = 8'h17; #100;
A = 8'h65; B = 8'h18; #100;
A = 8'h65; B = 8'h19; #100;
A = 8'h65; B = 8'h1A; #100;
A = 8'h65; B = 8'h1B; #100;
A = 8'h65; B = 8'h1C; #100;
A = 8'h65; B = 8'h1D; #100;
A = 8'h65; B = 8'h1E; #100;
A = 8'h65; B = 8'h1F; #100;
A = 8'h65; B = 8'h20; #100;
A = 8'h65; B = 8'h21; #100;
A = 8'h65; B = 8'h22; #100;
A = 8'h65; B = 8'h23; #100;
A = 8'h65; B = 8'h24; #100;
A = 8'h65; B = 8'h25; #100;
A = 8'h65; B = 8'h26; #100;
A = 8'h65; B = 8'h27; #100;
A = 8'h65; B = 8'h28; #100;
A = 8'h65; B = 8'h29; #100;
A = 8'h65; B = 8'h2A; #100;
A = 8'h65; B = 8'h2B; #100;
A = 8'h65; B = 8'h2C; #100;
A = 8'h65; B = 8'h2D; #100;
A = 8'h65; B = 8'h2E; #100;
A = 8'h65; B = 8'h2F; #100;
A = 8'h65; B = 8'h30; #100;
A = 8'h65; B = 8'h31; #100;
A = 8'h65; B = 8'h32; #100;
A = 8'h65; B = 8'h33; #100;
A = 8'h65; B = 8'h34; #100;
A = 8'h65; B = 8'h35; #100;
A = 8'h65; B = 8'h36; #100;
A = 8'h65; B = 8'h37; #100;
A = 8'h65; B = 8'h38; #100;
A = 8'h65; B = 8'h39; #100;
A = 8'h65; B = 8'h3A; #100;
A = 8'h65; B = 8'h3B; #100;
A = 8'h65; B = 8'h3C; #100;
A = 8'h65; B = 8'h3D; #100;
A = 8'h65; B = 8'h3E; #100;
A = 8'h65; B = 8'h3F; #100;
A = 8'h65; B = 8'h40; #100;
A = 8'h65; B = 8'h41; #100;
A = 8'h65; B = 8'h42; #100;
A = 8'h65; B = 8'h43; #100;
A = 8'h65; B = 8'h44; #100;
A = 8'h65; B = 8'h45; #100;
A = 8'h65; B = 8'h46; #100;
A = 8'h65; B = 8'h47; #100;
A = 8'h65; B = 8'h48; #100;
A = 8'h65; B = 8'h49; #100;
A = 8'h65; B = 8'h4A; #100;
A = 8'h65; B = 8'h4B; #100;
A = 8'h65; B = 8'h4C; #100;
A = 8'h65; B = 8'h4D; #100;
A = 8'h65; B = 8'h4E; #100;
A = 8'h65; B = 8'h4F; #100;
A = 8'h65; B = 8'h50; #100;
A = 8'h65; B = 8'h51; #100;
A = 8'h65; B = 8'h52; #100;
A = 8'h65; B = 8'h53; #100;
A = 8'h65; B = 8'h54; #100;
A = 8'h65; B = 8'h55; #100;
A = 8'h65; B = 8'h56; #100;
A = 8'h65; B = 8'h57; #100;
A = 8'h65; B = 8'h58; #100;
A = 8'h65; B = 8'h59; #100;
A = 8'h65; B = 8'h5A; #100;
A = 8'h65; B = 8'h5B; #100;
A = 8'h65; B = 8'h5C; #100;
A = 8'h65; B = 8'h5D; #100;
A = 8'h65; B = 8'h5E; #100;
A = 8'h65; B = 8'h5F; #100;
A = 8'h65; B = 8'h60; #100;
A = 8'h65; B = 8'h61; #100;
A = 8'h65; B = 8'h62; #100;
A = 8'h65; B = 8'h63; #100;
A = 8'h65; B = 8'h64; #100;
A = 8'h65; B = 8'h65; #100;
A = 8'h65; B = 8'h66; #100;
A = 8'h65; B = 8'h67; #100;
A = 8'h65; B = 8'h68; #100;
A = 8'h65; B = 8'h69; #100;
A = 8'h65; B = 8'h6A; #100;
A = 8'h65; B = 8'h6B; #100;
A = 8'h65; B = 8'h6C; #100;
A = 8'h65; B = 8'h6D; #100;
A = 8'h65; B = 8'h6E; #100;
A = 8'h65; B = 8'h6F; #100;
A = 8'h65; B = 8'h70; #100;
A = 8'h65; B = 8'h71; #100;
A = 8'h65; B = 8'h72; #100;
A = 8'h65; B = 8'h73; #100;
A = 8'h65; B = 8'h74; #100;
A = 8'h65; B = 8'h75; #100;
A = 8'h65; B = 8'h76; #100;
A = 8'h65; B = 8'h77; #100;
A = 8'h65; B = 8'h78; #100;
A = 8'h65; B = 8'h79; #100;
A = 8'h65; B = 8'h7A; #100;
A = 8'h65; B = 8'h7B; #100;
A = 8'h65; B = 8'h7C; #100;
A = 8'h65; B = 8'h7D; #100;
A = 8'h65; B = 8'h7E; #100;
A = 8'h65; B = 8'h7F; #100;
A = 8'h65; B = 8'h80; #100;
A = 8'h65; B = 8'h81; #100;
A = 8'h65; B = 8'h82; #100;
A = 8'h65; B = 8'h83; #100;
A = 8'h65; B = 8'h84; #100;
A = 8'h65; B = 8'h85; #100;
A = 8'h65; B = 8'h86; #100;
A = 8'h65; B = 8'h87; #100;
A = 8'h65; B = 8'h88; #100;
A = 8'h65; B = 8'h89; #100;
A = 8'h65; B = 8'h8A; #100;
A = 8'h65; B = 8'h8B; #100;
A = 8'h65; B = 8'h8C; #100;
A = 8'h65; B = 8'h8D; #100;
A = 8'h65; B = 8'h8E; #100;
A = 8'h65; B = 8'h8F; #100;
A = 8'h65; B = 8'h90; #100;
A = 8'h65; B = 8'h91; #100;
A = 8'h65; B = 8'h92; #100;
A = 8'h65; B = 8'h93; #100;
A = 8'h65; B = 8'h94; #100;
A = 8'h65; B = 8'h95; #100;
A = 8'h65; B = 8'h96; #100;
A = 8'h65; B = 8'h97; #100;
A = 8'h65; B = 8'h98; #100;
A = 8'h65; B = 8'h99; #100;
A = 8'h65; B = 8'h9A; #100;
A = 8'h65; B = 8'h9B; #100;
A = 8'h65; B = 8'h9C; #100;
A = 8'h65; B = 8'h9D; #100;
A = 8'h65; B = 8'h9E; #100;
A = 8'h65; B = 8'h9F; #100;
A = 8'h65; B = 8'hA0; #100;
A = 8'h65; B = 8'hA1; #100;
A = 8'h65; B = 8'hA2; #100;
A = 8'h65; B = 8'hA3; #100;
A = 8'h65; B = 8'hA4; #100;
A = 8'h65; B = 8'hA5; #100;
A = 8'h65; B = 8'hA6; #100;
A = 8'h65; B = 8'hA7; #100;
A = 8'h65; B = 8'hA8; #100;
A = 8'h65; B = 8'hA9; #100;
A = 8'h65; B = 8'hAA; #100;
A = 8'h65; B = 8'hAB; #100;
A = 8'h65; B = 8'hAC; #100;
A = 8'h65; B = 8'hAD; #100;
A = 8'h65; B = 8'hAE; #100;
A = 8'h65; B = 8'hAF; #100;
A = 8'h65; B = 8'hB0; #100;
A = 8'h65; B = 8'hB1; #100;
A = 8'h65; B = 8'hB2; #100;
A = 8'h65; B = 8'hB3; #100;
A = 8'h65; B = 8'hB4; #100;
A = 8'h65; B = 8'hB5; #100;
A = 8'h65; B = 8'hB6; #100;
A = 8'h65; B = 8'hB7; #100;
A = 8'h65; B = 8'hB8; #100;
A = 8'h65; B = 8'hB9; #100;
A = 8'h65; B = 8'hBA; #100;
A = 8'h65; B = 8'hBB; #100;
A = 8'h65; B = 8'hBC; #100;
A = 8'h65; B = 8'hBD; #100;
A = 8'h65; B = 8'hBE; #100;
A = 8'h65; B = 8'hBF; #100;
A = 8'h65; B = 8'hC0; #100;
A = 8'h65; B = 8'hC1; #100;
A = 8'h65; B = 8'hC2; #100;
A = 8'h65; B = 8'hC3; #100;
A = 8'h65; B = 8'hC4; #100;
A = 8'h65; B = 8'hC5; #100;
A = 8'h65; B = 8'hC6; #100;
A = 8'h65; B = 8'hC7; #100;
A = 8'h65; B = 8'hC8; #100;
A = 8'h65; B = 8'hC9; #100;
A = 8'h65; B = 8'hCA; #100;
A = 8'h65; B = 8'hCB; #100;
A = 8'h65; B = 8'hCC; #100;
A = 8'h65; B = 8'hCD; #100;
A = 8'h65; B = 8'hCE; #100;
A = 8'h65; B = 8'hCF; #100;
A = 8'h65; B = 8'hD0; #100;
A = 8'h65; B = 8'hD1; #100;
A = 8'h65; B = 8'hD2; #100;
A = 8'h65; B = 8'hD3; #100;
A = 8'h65; B = 8'hD4; #100;
A = 8'h65; B = 8'hD5; #100;
A = 8'h65; B = 8'hD6; #100;
A = 8'h65; B = 8'hD7; #100;
A = 8'h65; B = 8'hD8; #100;
A = 8'h65; B = 8'hD9; #100;
A = 8'h65; B = 8'hDA; #100;
A = 8'h65; B = 8'hDB; #100;
A = 8'h65; B = 8'hDC; #100;
A = 8'h65; B = 8'hDD; #100;
A = 8'h65; B = 8'hDE; #100;
A = 8'h65; B = 8'hDF; #100;
A = 8'h65; B = 8'hE0; #100;
A = 8'h65; B = 8'hE1; #100;
A = 8'h65; B = 8'hE2; #100;
A = 8'h65; B = 8'hE3; #100;
A = 8'h65; B = 8'hE4; #100;
A = 8'h65; B = 8'hE5; #100;
A = 8'h65; B = 8'hE6; #100;
A = 8'h65; B = 8'hE7; #100;
A = 8'h65; B = 8'hE8; #100;
A = 8'h65; B = 8'hE9; #100;
A = 8'h65; B = 8'hEA; #100;
A = 8'h65; B = 8'hEB; #100;
A = 8'h65; B = 8'hEC; #100;
A = 8'h65; B = 8'hED; #100;
A = 8'h65; B = 8'hEE; #100;
A = 8'h65; B = 8'hEF; #100;
A = 8'h65; B = 8'hF0; #100;
A = 8'h65; B = 8'hF1; #100;
A = 8'h65; B = 8'hF2; #100;
A = 8'h65; B = 8'hF3; #100;
A = 8'h65; B = 8'hF4; #100;
A = 8'h65; B = 8'hF5; #100;
A = 8'h65; B = 8'hF6; #100;
A = 8'h65; B = 8'hF7; #100;
A = 8'h65; B = 8'hF8; #100;
A = 8'h65; B = 8'hF9; #100;
A = 8'h65; B = 8'hFA; #100;
A = 8'h65; B = 8'hFB; #100;
A = 8'h65; B = 8'hFC; #100;
A = 8'h65; B = 8'hFD; #100;
A = 8'h65; B = 8'hFE; #100;
A = 8'h65; B = 8'hFF; #100;
A = 8'h66; B = 8'h0; #100;
A = 8'h66; B = 8'h1; #100;
A = 8'h66; B = 8'h2; #100;
A = 8'h66; B = 8'h3; #100;
A = 8'h66; B = 8'h4; #100;
A = 8'h66; B = 8'h5; #100;
A = 8'h66; B = 8'h6; #100;
A = 8'h66; B = 8'h7; #100;
A = 8'h66; B = 8'h8; #100;
A = 8'h66; B = 8'h9; #100;
A = 8'h66; B = 8'hA; #100;
A = 8'h66; B = 8'hB; #100;
A = 8'h66; B = 8'hC; #100;
A = 8'h66; B = 8'hD; #100;
A = 8'h66; B = 8'hE; #100;
A = 8'h66; B = 8'hF; #100;
A = 8'h66; B = 8'h10; #100;
A = 8'h66; B = 8'h11; #100;
A = 8'h66; B = 8'h12; #100;
A = 8'h66; B = 8'h13; #100;
A = 8'h66; B = 8'h14; #100;
A = 8'h66; B = 8'h15; #100;
A = 8'h66; B = 8'h16; #100;
A = 8'h66; B = 8'h17; #100;
A = 8'h66; B = 8'h18; #100;
A = 8'h66; B = 8'h19; #100;
A = 8'h66; B = 8'h1A; #100;
A = 8'h66; B = 8'h1B; #100;
A = 8'h66; B = 8'h1C; #100;
A = 8'h66; B = 8'h1D; #100;
A = 8'h66; B = 8'h1E; #100;
A = 8'h66; B = 8'h1F; #100;
A = 8'h66; B = 8'h20; #100;
A = 8'h66; B = 8'h21; #100;
A = 8'h66; B = 8'h22; #100;
A = 8'h66; B = 8'h23; #100;
A = 8'h66; B = 8'h24; #100;
A = 8'h66; B = 8'h25; #100;
A = 8'h66; B = 8'h26; #100;
A = 8'h66; B = 8'h27; #100;
A = 8'h66; B = 8'h28; #100;
A = 8'h66; B = 8'h29; #100;
A = 8'h66; B = 8'h2A; #100;
A = 8'h66; B = 8'h2B; #100;
A = 8'h66; B = 8'h2C; #100;
A = 8'h66; B = 8'h2D; #100;
A = 8'h66; B = 8'h2E; #100;
A = 8'h66; B = 8'h2F; #100;
A = 8'h66; B = 8'h30; #100;
A = 8'h66; B = 8'h31; #100;
A = 8'h66; B = 8'h32; #100;
A = 8'h66; B = 8'h33; #100;
A = 8'h66; B = 8'h34; #100;
A = 8'h66; B = 8'h35; #100;
A = 8'h66; B = 8'h36; #100;
A = 8'h66; B = 8'h37; #100;
A = 8'h66; B = 8'h38; #100;
A = 8'h66; B = 8'h39; #100;
A = 8'h66; B = 8'h3A; #100;
A = 8'h66; B = 8'h3B; #100;
A = 8'h66; B = 8'h3C; #100;
A = 8'h66; B = 8'h3D; #100;
A = 8'h66; B = 8'h3E; #100;
A = 8'h66; B = 8'h3F; #100;
A = 8'h66; B = 8'h40; #100;
A = 8'h66; B = 8'h41; #100;
A = 8'h66; B = 8'h42; #100;
A = 8'h66; B = 8'h43; #100;
A = 8'h66; B = 8'h44; #100;
A = 8'h66; B = 8'h45; #100;
A = 8'h66; B = 8'h46; #100;
A = 8'h66; B = 8'h47; #100;
A = 8'h66; B = 8'h48; #100;
A = 8'h66; B = 8'h49; #100;
A = 8'h66; B = 8'h4A; #100;
A = 8'h66; B = 8'h4B; #100;
A = 8'h66; B = 8'h4C; #100;
A = 8'h66; B = 8'h4D; #100;
A = 8'h66; B = 8'h4E; #100;
A = 8'h66; B = 8'h4F; #100;
A = 8'h66; B = 8'h50; #100;
A = 8'h66; B = 8'h51; #100;
A = 8'h66; B = 8'h52; #100;
A = 8'h66; B = 8'h53; #100;
A = 8'h66; B = 8'h54; #100;
A = 8'h66; B = 8'h55; #100;
A = 8'h66; B = 8'h56; #100;
A = 8'h66; B = 8'h57; #100;
A = 8'h66; B = 8'h58; #100;
A = 8'h66; B = 8'h59; #100;
A = 8'h66; B = 8'h5A; #100;
A = 8'h66; B = 8'h5B; #100;
A = 8'h66; B = 8'h5C; #100;
A = 8'h66; B = 8'h5D; #100;
A = 8'h66; B = 8'h5E; #100;
A = 8'h66; B = 8'h5F; #100;
A = 8'h66; B = 8'h60; #100;
A = 8'h66; B = 8'h61; #100;
A = 8'h66; B = 8'h62; #100;
A = 8'h66; B = 8'h63; #100;
A = 8'h66; B = 8'h64; #100;
A = 8'h66; B = 8'h65; #100;
A = 8'h66; B = 8'h66; #100;
A = 8'h66; B = 8'h67; #100;
A = 8'h66; B = 8'h68; #100;
A = 8'h66; B = 8'h69; #100;
A = 8'h66; B = 8'h6A; #100;
A = 8'h66; B = 8'h6B; #100;
A = 8'h66; B = 8'h6C; #100;
A = 8'h66; B = 8'h6D; #100;
A = 8'h66; B = 8'h6E; #100;
A = 8'h66; B = 8'h6F; #100;
A = 8'h66; B = 8'h70; #100;
A = 8'h66; B = 8'h71; #100;
A = 8'h66; B = 8'h72; #100;
A = 8'h66; B = 8'h73; #100;
A = 8'h66; B = 8'h74; #100;
A = 8'h66; B = 8'h75; #100;
A = 8'h66; B = 8'h76; #100;
A = 8'h66; B = 8'h77; #100;
A = 8'h66; B = 8'h78; #100;
A = 8'h66; B = 8'h79; #100;
A = 8'h66; B = 8'h7A; #100;
A = 8'h66; B = 8'h7B; #100;
A = 8'h66; B = 8'h7C; #100;
A = 8'h66; B = 8'h7D; #100;
A = 8'h66; B = 8'h7E; #100;
A = 8'h66; B = 8'h7F; #100;
A = 8'h66; B = 8'h80; #100;
A = 8'h66; B = 8'h81; #100;
A = 8'h66; B = 8'h82; #100;
A = 8'h66; B = 8'h83; #100;
A = 8'h66; B = 8'h84; #100;
A = 8'h66; B = 8'h85; #100;
A = 8'h66; B = 8'h86; #100;
A = 8'h66; B = 8'h87; #100;
A = 8'h66; B = 8'h88; #100;
A = 8'h66; B = 8'h89; #100;
A = 8'h66; B = 8'h8A; #100;
A = 8'h66; B = 8'h8B; #100;
A = 8'h66; B = 8'h8C; #100;
A = 8'h66; B = 8'h8D; #100;
A = 8'h66; B = 8'h8E; #100;
A = 8'h66; B = 8'h8F; #100;
A = 8'h66; B = 8'h90; #100;
A = 8'h66; B = 8'h91; #100;
A = 8'h66; B = 8'h92; #100;
A = 8'h66; B = 8'h93; #100;
A = 8'h66; B = 8'h94; #100;
A = 8'h66; B = 8'h95; #100;
A = 8'h66; B = 8'h96; #100;
A = 8'h66; B = 8'h97; #100;
A = 8'h66; B = 8'h98; #100;
A = 8'h66; B = 8'h99; #100;
A = 8'h66; B = 8'h9A; #100;
A = 8'h66; B = 8'h9B; #100;
A = 8'h66; B = 8'h9C; #100;
A = 8'h66; B = 8'h9D; #100;
A = 8'h66; B = 8'h9E; #100;
A = 8'h66; B = 8'h9F; #100;
A = 8'h66; B = 8'hA0; #100;
A = 8'h66; B = 8'hA1; #100;
A = 8'h66; B = 8'hA2; #100;
A = 8'h66; B = 8'hA3; #100;
A = 8'h66; B = 8'hA4; #100;
A = 8'h66; B = 8'hA5; #100;
A = 8'h66; B = 8'hA6; #100;
A = 8'h66; B = 8'hA7; #100;
A = 8'h66; B = 8'hA8; #100;
A = 8'h66; B = 8'hA9; #100;
A = 8'h66; B = 8'hAA; #100;
A = 8'h66; B = 8'hAB; #100;
A = 8'h66; B = 8'hAC; #100;
A = 8'h66; B = 8'hAD; #100;
A = 8'h66; B = 8'hAE; #100;
A = 8'h66; B = 8'hAF; #100;
A = 8'h66; B = 8'hB0; #100;
A = 8'h66; B = 8'hB1; #100;
A = 8'h66; B = 8'hB2; #100;
A = 8'h66; B = 8'hB3; #100;
A = 8'h66; B = 8'hB4; #100;
A = 8'h66; B = 8'hB5; #100;
A = 8'h66; B = 8'hB6; #100;
A = 8'h66; B = 8'hB7; #100;
A = 8'h66; B = 8'hB8; #100;
A = 8'h66; B = 8'hB9; #100;
A = 8'h66; B = 8'hBA; #100;
A = 8'h66; B = 8'hBB; #100;
A = 8'h66; B = 8'hBC; #100;
A = 8'h66; B = 8'hBD; #100;
A = 8'h66; B = 8'hBE; #100;
A = 8'h66; B = 8'hBF; #100;
A = 8'h66; B = 8'hC0; #100;
A = 8'h66; B = 8'hC1; #100;
A = 8'h66; B = 8'hC2; #100;
A = 8'h66; B = 8'hC3; #100;
A = 8'h66; B = 8'hC4; #100;
A = 8'h66; B = 8'hC5; #100;
A = 8'h66; B = 8'hC6; #100;
A = 8'h66; B = 8'hC7; #100;
A = 8'h66; B = 8'hC8; #100;
A = 8'h66; B = 8'hC9; #100;
A = 8'h66; B = 8'hCA; #100;
A = 8'h66; B = 8'hCB; #100;
A = 8'h66; B = 8'hCC; #100;
A = 8'h66; B = 8'hCD; #100;
A = 8'h66; B = 8'hCE; #100;
A = 8'h66; B = 8'hCF; #100;
A = 8'h66; B = 8'hD0; #100;
A = 8'h66; B = 8'hD1; #100;
A = 8'h66; B = 8'hD2; #100;
A = 8'h66; B = 8'hD3; #100;
A = 8'h66; B = 8'hD4; #100;
A = 8'h66; B = 8'hD5; #100;
A = 8'h66; B = 8'hD6; #100;
A = 8'h66; B = 8'hD7; #100;
A = 8'h66; B = 8'hD8; #100;
A = 8'h66; B = 8'hD9; #100;
A = 8'h66; B = 8'hDA; #100;
A = 8'h66; B = 8'hDB; #100;
A = 8'h66; B = 8'hDC; #100;
A = 8'h66; B = 8'hDD; #100;
A = 8'h66; B = 8'hDE; #100;
A = 8'h66; B = 8'hDF; #100;
A = 8'h66; B = 8'hE0; #100;
A = 8'h66; B = 8'hE1; #100;
A = 8'h66; B = 8'hE2; #100;
A = 8'h66; B = 8'hE3; #100;
A = 8'h66; B = 8'hE4; #100;
A = 8'h66; B = 8'hE5; #100;
A = 8'h66; B = 8'hE6; #100;
A = 8'h66; B = 8'hE7; #100;
A = 8'h66; B = 8'hE8; #100;
A = 8'h66; B = 8'hE9; #100;
A = 8'h66; B = 8'hEA; #100;
A = 8'h66; B = 8'hEB; #100;
A = 8'h66; B = 8'hEC; #100;
A = 8'h66; B = 8'hED; #100;
A = 8'h66; B = 8'hEE; #100;
A = 8'h66; B = 8'hEF; #100;
A = 8'h66; B = 8'hF0; #100;
A = 8'h66; B = 8'hF1; #100;
A = 8'h66; B = 8'hF2; #100;
A = 8'h66; B = 8'hF3; #100;
A = 8'h66; B = 8'hF4; #100;
A = 8'h66; B = 8'hF5; #100;
A = 8'h66; B = 8'hF6; #100;
A = 8'h66; B = 8'hF7; #100;
A = 8'h66; B = 8'hF8; #100;
A = 8'h66; B = 8'hF9; #100;
A = 8'h66; B = 8'hFA; #100;
A = 8'h66; B = 8'hFB; #100;
A = 8'h66; B = 8'hFC; #100;
A = 8'h66; B = 8'hFD; #100;
A = 8'h66; B = 8'hFE; #100;
A = 8'h66; B = 8'hFF; #100;
A = 8'h67; B = 8'h0; #100;
A = 8'h67; B = 8'h1; #100;
A = 8'h67; B = 8'h2; #100;
A = 8'h67; B = 8'h3; #100;
A = 8'h67; B = 8'h4; #100;
A = 8'h67; B = 8'h5; #100;
A = 8'h67; B = 8'h6; #100;
A = 8'h67; B = 8'h7; #100;
A = 8'h67; B = 8'h8; #100;
A = 8'h67; B = 8'h9; #100;
A = 8'h67; B = 8'hA; #100;
A = 8'h67; B = 8'hB; #100;
A = 8'h67; B = 8'hC; #100;
A = 8'h67; B = 8'hD; #100;
A = 8'h67; B = 8'hE; #100;
A = 8'h67; B = 8'hF; #100;
A = 8'h67; B = 8'h10; #100;
A = 8'h67; B = 8'h11; #100;
A = 8'h67; B = 8'h12; #100;
A = 8'h67; B = 8'h13; #100;
A = 8'h67; B = 8'h14; #100;
A = 8'h67; B = 8'h15; #100;
A = 8'h67; B = 8'h16; #100;
A = 8'h67; B = 8'h17; #100;
A = 8'h67; B = 8'h18; #100;
A = 8'h67; B = 8'h19; #100;
A = 8'h67; B = 8'h1A; #100;
A = 8'h67; B = 8'h1B; #100;
A = 8'h67; B = 8'h1C; #100;
A = 8'h67; B = 8'h1D; #100;
A = 8'h67; B = 8'h1E; #100;
A = 8'h67; B = 8'h1F; #100;
A = 8'h67; B = 8'h20; #100;
A = 8'h67; B = 8'h21; #100;
A = 8'h67; B = 8'h22; #100;
A = 8'h67; B = 8'h23; #100;
A = 8'h67; B = 8'h24; #100;
A = 8'h67; B = 8'h25; #100;
A = 8'h67; B = 8'h26; #100;
A = 8'h67; B = 8'h27; #100;
A = 8'h67; B = 8'h28; #100;
A = 8'h67; B = 8'h29; #100;
A = 8'h67; B = 8'h2A; #100;
A = 8'h67; B = 8'h2B; #100;
A = 8'h67; B = 8'h2C; #100;
A = 8'h67; B = 8'h2D; #100;
A = 8'h67; B = 8'h2E; #100;
A = 8'h67; B = 8'h2F; #100;
A = 8'h67; B = 8'h30; #100;
A = 8'h67; B = 8'h31; #100;
A = 8'h67; B = 8'h32; #100;
A = 8'h67; B = 8'h33; #100;
A = 8'h67; B = 8'h34; #100;
A = 8'h67; B = 8'h35; #100;
A = 8'h67; B = 8'h36; #100;
A = 8'h67; B = 8'h37; #100;
A = 8'h67; B = 8'h38; #100;
A = 8'h67; B = 8'h39; #100;
A = 8'h67; B = 8'h3A; #100;
A = 8'h67; B = 8'h3B; #100;
A = 8'h67; B = 8'h3C; #100;
A = 8'h67; B = 8'h3D; #100;
A = 8'h67; B = 8'h3E; #100;
A = 8'h67; B = 8'h3F; #100;
A = 8'h67; B = 8'h40; #100;
A = 8'h67; B = 8'h41; #100;
A = 8'h67; B = 8'h42; #100;
A = 8'h67; B = 8'h43; #100;
A = 8'h67; B = 8'h44; #100;
A = 8'h67; B = 8'h45; #100;
A = 8'h67; B = 8'h46; #100;
A = 8'h67; B = 8'h47; #100;
A = 8'h67; B = 8'h48; #100;
A = 8'h67; B = 8'h49; #100;
A = 8'h67; B = 8'h4A; #100;
A = 8'h67; B = 8'h4B; #100;
A = 8'h67; B = 8'h4C; #100;
A = 8'h67; B = 8'h4D; #100;
A = 8'h67; B = 8'h4E; #100;
A = 8'h67; B = 8'h4F; #100;
A = 8'h67; B = 8'h50; #100;
A = 8'h67; B = 8'h51; #100;
A = 8'h67; B = 8'h52; #100;
A = 8'h67; B = 8'h53; #100;
A = 8'h67; B = 8'h54; #100;
A = 8'h67; B = 8'h55; #100;
A = 8'h67; B = 8'h56; #100;
A = 8'h67; B = 8'h57; #100;
A = 8'h67; B = 8'h58; #100;
A = 8'h67; B = 8'h59; #100;
A = 8'h67; B = 8'h5A; #100;
A = 8'h67; B = 8'h5B; #100;
A = 8'h67; B = 8'h5C; #100;
A = 8'h67; B = 8'h5D; #100;
A = 8'h67; B = 8'h5E; #100;
A = 8'h67; B = 8'h5F; #100;
A = 8'h67; B = 8'h60; #100;
A = 8'h67; B = 8'h61; #100;
A = 8'h67; B = 8'h62; #100;
A = 8'h67; B = 8'h63; #100;
A = 8'h67; B = 8'h64; #100;
A = 8'h67; B = 8'h65; #100;
A = 8'h67; B = 8'h66; #100;
A = 8'h67; B = 8'h67; #100;
A = 8'h67; B = 8'h68; #100;
A = 8'h67; B = 8'h69; #100;
A = 8'h67; B = 8'h6A; #100;
A = 8'h67; B = 8'h6B; #100;
A = 8'h67; B = 8'h6C; #100;
A = 8'h67; B = 8'h6D; #100;
A = 8'h67; B = 8'h6E; #100;
A = 8'h67; B = 8'h6F; #100;
A = 8'h67; B = 8'h70; #100;
A = 8'h67; B = 8'h71; #100;
A = 8'h67; B = 8'h72; #100;
A = 8'h67; B = 8'h73; #100;
A = 8'h67; B = 8'h74; #100;
A = 8'h67; B = 8'h75; #100;
A = 8'h67; B = 8'h76; #100;
A = 8'h67; B = 8'h77; #100;
A = 8'h67; B = 8'h78; #100;
A = 8'h67; B = 8'h79; #100;
A = 8'h67; B = 8'h7A; #100;
A = 8'h67; B = 8'h7B; #100;
A = 8'h67; B = 8'h7C; #100;
A = 8'h67; B = 8'h7D; #100;
A = 8'h67; B = 8'h7E; #100;
A = 8'h67; B = 8'h7F; #100;
A = 8'h67; B = 8'h80; #100;
A = 8'h67; B = 8'h81; #100;
A = 8'h67; B = 8'h82; #100;
A = 8'h67; B = 8'h83; #100;
A = 8'h67; B = 8'h84; #100;
A = 8'h67; B = 8'h85; #100;
A = 8'h67; B = 8'h86; #100;
A = 8'h67; B = 8'h87; #100;
A = 8'h67; B = 8'h88; #100;
A = 8'h67; B = 8'h89; #100;
A = 8'h67; B = 8'h8A; #100;
A = 8'h67; B = 8'h8B; #100;
A = 8'h67; B = 8'h8C; #100;
A = 8'h67; B = 8'h8D; #100;
A = 8'h67; B = 8'h8E; #100;
A = 8'h67; B = 8'h8F; #100;
A = 8'h67; B = 8'h90; #100;
A = 8'h67; B = 8'h91; #100;
A = 8'h67; B = 8'h92; #100;
A = 8'h67; B = 8'h93; #100;
A = 8'h67; B = 8'h94; #100;
A = 8'h67; B = 8'h95; #100;
A = 8'h67; B = 8'h96; #100;
A = 8'h67; B = 8'h97; #100;
A = 8'h67; B = 8'h98; #100;
A = 8'h67; B = 8'h99; #100;
A = 8'h67; B = 8'h9A; #100;
A = 8'h67; B = 8'h9B; #100;
A = 8'h67; B = 8'h9C; #100;
A = 8'h67; B = 8'h9D; #100;
A = 8'h67; B = 8'h9E; #100;
A = 8'h67; B = 8'h9F; #100;
A = 8'h67; B = 8'hA0; #100;
A = 8'h67; B = 8'hA1; #100;
A = 8'h67; B = 8'hA2; #100;
A = 8'h67; B = 8'hA3; #100;
A = 8'h67; B = 8'hA4; #100;
A = 8'h67; B = 8'hA5; #100;
A = 8'h67; B = 8'hA6; #100;
A = 8'h67; B = 8'hA7; #100;
A = 8'h67; B = 8'hA8; #100;
A = 8'h67; B = 8'hA9; #100;
A = 8'h67; B = 8'hAA; #100;
A = 8'h67; B = 8'hAB; #100;
A = 8'h67; B = 8'hAC; #100;
A = 8'h67; B = 8'hAD; #100;
A = 8'h67; B = 8'hAE; #100;
A = 8'h67; B = 8'hAF; #100;
A = 8'h67; B = 8'hB0; #100;
A = 8'h67; B = 8'hB1; #100;
A = 8'h67; B = 8'hB2; #100;
A = 8'h67; B = 8'hB3; #100;
A = 8'h67; B = 8'hB4; #100;
A = 8'h67; B = 8'hB5; #100;
A = 8'h67; B = 8'hB6; #100;
A = 8'h67; B = 8'hB7; #100;
A = 8'h67; B = 8'hB8; #100;
A = 8'h67; B = 8'hB9; #100;
A = 8'h67; B = 8'hBA; #100;
A = 8'h67; B = 8'hBB; #100;
A = 8'h67; B = 8'hBC; #100;
A = 8'h67; B = 8'hBD; #100;
A = 8'h67; B = 8'hBE; #100;
A = 8'h67; B = 8'hBF; #100;
A = 8'h67; B = 8'hC0; #100;
A = 8'h67; B = 8'hC1; #100;
A = 8'h67; B = 8'hC2; #100;
A = 8'h67; B = 8'hC3; #100;
A = 8'h67; B = 8'hC4; #100;
A = 8'h67; B = 8'hC5; #100;
A = 8'h67; B = 8'hC6; #100;
A = 8'h67; B = 8'hC7; #100;
A = 8'h67; B = 8'hC8; #100;
A = 8'h67; B = 8'hC9; #100;
A = 8'h67; B = 8'hCA; #100;
A = 8'h67; B = 8'hCB; #100;
A = 8'h67; B = 8'hCC; #100;
A = 8'h67; B = 8'hCD; #100;
A = 8'h67; B = 8'hCE; #100;
A = 8'h67; B = 8'hCF; #100;
A = 8'h67; B = 8'hD0; #100;
A = 8'h67; B = 8'hD1; #100;
A = 8'h67; B = 8'hD2; #100;
A = 8'h67; B = 8'hD3; #100;
A = 8'h67; B = 8'hD4; #100;
A = 8'h67; B = 8'hD5; #100;
A = 8'h67; B = 8'hD6; #100;
A = 8'h67; B = 8'hD7; #100;
A = 8'h67; B = 8'hD8; #100;
A = 8'h67; B = 8'hD9; #100;
A = 8'h67; B = 8'hDA; #100;
A = 8'h67; B = 8'hDB; #100;
A = 8'h67; B = 8'hDC; #100;
A = 8'h67; B = 8'hDD; #100;
A = 8'h67; B = 8'hDE; #100;
A = 8'h67; B = 8'hDF; #100;
A = 8'h67; B = 8'hE0; #100;
A = 8'h67; B = 8'hE1; #100;
A = 8'h67; B = 8'hE2; #100;
A = 8'h67; B = 8'hE3; #100;
A = 8'h67; B = 8'hE4; #100;
A = 8'h67; B = 8'hE5; #100;
A = 8'h67; B = 8'hE6; #100;
A = 8'h67; B = 8'hE7; #100;
A = 8'h67; B = 8'hE8; #100;
A = 8'h67; B = 8'hE9; #100;
A = 8'h67; B = 8'hEA; #100;
A = 8'h67; B = 8'hEB; #100;
A = 8'h67; B = 8'hEC; #100;
A = 8'h67; B = 8'hED; #100;
A = 8'h67; B = 8'hEE; #100;
A = 8'h67; B = 8'hEF; #100;
A = 8'h67; B = 8'hF0; #100;
A = 8'h67; B = 8'hF1; #100;
A = 8'h67; B = 8'hF2; #100;
A = 8'h67; B = 8'hF3; #100;
A = 8'h67; B = 8'hF4; #100;
A = 8'h67; B = 8'hF5; #100;
A = 8'h67; B = 8'hF6; #100;
A = 8'h67; B = 8'hF7; #100;
A = 8'h67; B = 8'hF8; #100;
A = 8'h67; B = 8'hF9; #100;
A = 8'h67; B = 8'hFA; #100;
A = 8'h67; B = 8'hFB; #100;
A = 8'h67; B = 8'hFC; #100;
A = 8'h67; B = 8'hFD; #100;
A = 8'h67; B = 8'hFE; #100;
A = 8'h67; B = 8'hFF; #100;
A = 8'h68; B = 8'h0; #100;
A = 8'h68; B = 8'h1; #100;
A = 8'h68; B = 8'h2; #100;
A = 8'h68; B = 8'h3; #100;
A = 8'h68; B = 8'h4; #100;
A = 8'h68; B = 8'h5; #100;
A = 8'h68; B = 8'h6; #100;
A = 8'h68; B = 8'h7; #100;
A = 8'h68; B = 8'h8; #100;
A = 8'h68; B = 8'h9; #100;
A = 8'h68; B = 8'hA; #100;
A = 8'h68; B = 8'hB; #100;
A = 8'h68; B = 8'hC; #100;
A = 8'h68; B = 8'hD; #100;
A = 8'h68; B = 8'hE; #100;
A = 8'h68; B = 8'hF; #100;
A = 8'h68; B = 8'h10; #100;
A = 8'h68; B = 8'h11; #100;
A = 8'h68; B = 8'h12; #100;
A = 8'h68; B = 8'h13; #100;
A = 8'h68; B = 8'h14; #100;
A = 8'h68; B = 8'h15; #100;
A = 8'h68; B = 8'h16; #100;
A = 8'h68; B = 8'h17; #100;
A = 8'h68; B = 8'h18; #100;
A = 8'h68; B = 8'h19; #100;
A = 8'h68; B = 8'h1A; #100;
A = 8'h68; B = 8'h1B; #100;
A = 8'h68; B = 8'h1C; #100;
A = 8'h68; B = 8'h1D; #100;
A = 8'h68; B = 8'h1E; #100;
A = 8'h68; B = 8'h1F; #100;
A = 8'h68; B = 8'h20; #100;
A = 8'h68; B = 8'h21; #100;
A = 8'h68; B = 8'h22; #100;
A = 8'h68; B = 8'h23; #100;
A = 8'h68; B = 8'h24; #100;
A = 8'h68; B = 8'h25; #100;
A = 8'h68; B = 8'h26; #100;
A = 8'h68; B = 8'h27; #100;
A = 8'h68; B = 8'h28; #100;
A = 8'h68; B = 8'h29; #100;
A = 8'h68; B = 8'h2A; #100;
A = 8'h68; B = 8'h2B; #100;
A = 8'h68; B = 8'h2C; #100;
A = 8'h68; B = 8'h2D; #100;
A = 8'h68; B = 8'h2E; #100;
A = 8'h68; B = 8'h2F; #100;
A = 8'h68; B = 8'h30; #100;
A = 8'h68; B = 8'h31; #100;
A = 8'h68; B = 8'h32; #100;
A = 8'h68; B = 8'h33; #100;
A = 8'h68; B = 8'h34; #100;
A = 8'h68; B = 8'h35; #100;
A = 8'h68; B = 8'h36; #100;
A = 8'h68; B = 8'h37; #100;
A = 8'h68; B = 8'h38; #100;
A = 8'h68; B = 8'h39; #100;
A = 8'h68; B = 8'h3A; #100;
A = 8'h68; B = 8'h3B; #100;
A = 8'h68; B = 8'h3C; #100;
A = 8'h68; B = 8'h3D; #100;
A = 8'h68; B = 8'h3E; #100;
A = 8'h68; B = 8'h3F; #100;
A = 8'h68; B = 8'h40; #100;
A = 8'h68; B = 8'h41; #100;
A = 8'h68; B = 8'h42; #100;
A = 8'h68; B = 8'h43; #100;
A = 8'h68; B = 8'h44; #100;
A = 8'h68; B = 8'h45; #100;
A = 8'h68; B = 8'h46; #100;
A = 8'h68; B = 8'h47; #100;
A = 8'h68; B = 8'h48; #100;
A = 8'h68; B = 8'h49; #100;
A = 8'h68; B = 8'h4A; #100;
A = 8'h68; B = 8'h4B; #100;
A = 8'h68; B = 8'h4C; #100;
A = 8'h68; B = 8'h4D; #100;
A = 8'h68; B = 8'h4E; #100;
A = 8'h68; B = 8'h4F; #100;
A = 8'h68; B = 8'h50; #100;
A = 8'h68; B = 8'h51; #100;
A = 8'h68; B = 8'h52; #100;
A = 8'h68; B = 8'h53; #100;
A = 8'h68; B = 8'h54; #100;
A = 8'h68; B = 8'h55; #100;
A = 8'h68; B = 8'h56; #100;
A = 8'h68; B = 8'h57; #100;
A = 8'h68; B = 8'h58; #100;
A = 8'h68; B = 8'h59; #100;
A = 8'h68; B = 8'h5A; #100;
A = 8'h68; B = 8'h5B; #100;
A = 8'h68; B = 8'h5C; #100;
A = 8'h68; B = 8'h5D; #100;
A = 8'h68; B = 8'h5E; #100;
A = 8'h68; B = 8'h5F; #100;
A = 8'h68; B = 8'h60; #100;
A = 8'h68; B = 8'h61; #100;
A = 8'h68; B = 8'h62; #100;
A = 8'h68; B = 8'h63; #100;
A = 8'h68; B = 8'h64; #100;
A = 8'h68; B = 8'h65; #100;
A = 8'h68; B = 8'h66; #100;
A = 8'h68; B = 8'h67; #100;
A = 8'h68; B = 8'h68; #100;
A = 8'h68; B = 8'h69; #100;
A = 8'h68; B = 8'h6A; #100;
A = 8'h68; B = 8'h6B; #100;
A = 8'h68; B = 8'h6C; #100;
A = 8'h68; B = 8'h6D; #100;
A = 8'h68; B = 8'h6E; #100;
A = 8'h68; B = 8'h6F; #100;
A = 8'h68; B = 8'h70; #100;
A = 8'h68; B = 8'h71; #100;
A = 8'h68; B = 8'h72; #100;
A = 8'h68; B = 8'h73; #100;
A = 8'h68; B = 8'h74; #100;
A = 8'h68; B = 8'h75; #100;
A = 8'h68; B = 8'h76; #100;
A = 8'h68; B = 8'h77; #100;
A = 8'h68; B = 8'h78; #100;
A = 8'h68; B = 8'h79; #100;
A = 8'h68; B = 8'h7A; #100;
A = 8'h68; B = 8'h7B; #100;
A = 8'h68; B = 8'h7C; #100;
A = 8'h68; B = 8'h7D; #100;
A = 8'h68; B = 8'h7E; #100;
A = 8'h68; B = 8'h7F; #100;
A = 8'h68; B = 8'h80; #100;
A = 8'h68; B = 8'h81; #100;
A = 8'h68; B = 8'h82; #100;
A = 8'h68; B = 8'h83; #100;
A = 8'h68; B = 8'h84; #100;
A = 8'h68; B = 8'h85; #100;
A = 8'h68; B = 8'h86; #100;
A = 8'h68; B = 8'h87; #100;
A = 8'h68; B = 8'h88; #100;
A = 8'h68; B = 8'h89; #100;
A = 8'h68; B = 8'h8A; #100;
A = 8'h68; B = 8'h8B; #100;
A = 8'h68; B = 8'h8C; #100;
A = 8'h68; B = 8'h8D; #100;
A = 8'h68; B = 8'h8E; #100;
A = 8'h68; B = 8'h8F; #100;
A = 8'h68; B = 8'h90; #100;
A = 8'h68; B = 8'h91; #100;
A = 8'h68; B = 8'h92; #100;
A = 8'h68; B = 8'h93; #100;
A = 8'h68; B = 8'h94; #100;
A = 8'h68; B = 8'h95; #100;
A = 8'h68; B = 8'h96; #100;
A = 8'h68; B = 8'h97; #100;
A = 8'h68; B = 8'h98; #100;
A = 8'h68; B = 8'h99; #100;
A = 8'h68; B = 8'h9A; #100;
A = 8'h68; B = 8'h9B; #100;
A = 8'h68; B = 8'h9C; #100;
A = 8'h68; B = 8'h9D; #100;
A = 8'h68; B = 8'h9E; #100;
A = 8'h68; B = 8'h9F; #100;
A = 8'h68; B = 8'hA0; #100;
A = 8'h68; B = 8'hA1; #100;
A = 8'h68; B = 8'hA2; #100;
A = 8'h68; B = 8'hA3; #100;
A = 8'h68; B = 8'hA4; #100;
A = 8'h68; B = 8'hA5; #100;
A = 8'h68; B = 8'hA6; #100;
A = 8'h68; B = 8'hA7; #100;
A = 8'h68; B = 8'hA8; #100;
A = 8'h68; B = 8'hA9; #100;
A = 8'h68; B = 8'hAA; #100;
A = 8'h68; B = 8'hAB; #100;
A = 8'h68; B = 8'hAC; #100;
A = 8'h68; B = 8'hAD; #100;
A = 8'h68; B = 8'hAE; #100;
A = 8'h68; B = 8'hAF; #100;
A = 8'h68; B = 8'hB0; #100;
A = 8'h68; B = 8'hB1; #100;
A = 8'h68; B = 8'hB2; #100;
A = 8'h68; B = 8'hB3; #100;
A = 8'h68; B = 8'hB4; #100;
A = 8'h68; B = 8'hB5; #100;
A = 8'h68; B = 8'hB6; #100;
A = 8'h68; B = 8'hB7; #100;
A = 8'h68; B = 8'hB8; #100;
A = 8'h68; B = 8'hB9; #100;
A = 8'h68; B = 8'hBA; #100;
A = 8'h68; B = 8'hBB; #100;
A = 8'h68; B = 8'hBC; #100;
A = 8'h68; B = 8'hBD; #100;
A = 8'h68; B = 8'hBE; #100;
A = 8'h68; B = 8'hBF; #100;
A = 8'h68; B = 8'hC0; #100;
A = 8'h68; B = 8'hC1; #100;
A = 8'h68; B = 8'hC2; #100;
A = 8'h68; B = 8'hC3; #100;
A = 8'h68; B = 8'hC4; #100;
A = 8'h68; B = 8'hC5; #100;
A = 8'h68; B = 8'hC6; #100;
A = 8'h68; B = 8'hC7; #100;
A = 8'h68; B = 8'hC8; #100;
A = 8'h68; B = 8'hC9; #100;
A = 8'h68; B = 8'hCA; #100;
A = 8'h68; B = 8'hCB; #100;
A = 8'h68; B = 8'hCC; #100;
A = 8'h68; B = 8'hCD; #100;
A = 8'h68; B = 8'hCE; #100;
A = 8'h68; B = 8'hCF; #100;
A = 8'h68; B = 8'hD0; #100;
A = 8'h68; B = 8'hD1; #100;
A = 8'h68; B = 8'hD2; #100;
A = 8'h68; B = 8'hD3; #100;
A = 8'h68; B = 8'hD4; #100;
A = 8'h68; B = 8'hD5; #100;
A = 8'h68; B = 8'hD6; #100;
A = 8'h68; B = 8'hD7; #100;
A = 8'h68; B = 8'hD8; #100;
A = 8'h68; B = 8'hD9; #100;
A = 8'h68; B = 8'hDA; #100;
A = 8'h68; B = 8'hDB; #100;
A = 8'h68; B = 8'hDC; #100;
A = 8'h68; B = 8'hDD; #100;
A = 8'h68; B = 8'hDE; #100;
A = 8'h68; B = 8'hDF; #100;
A = 8'h68; B = 8'hE0; #100;
A = 8'h68; B = 8'hE1; #100;
A = 8'h68; B = 8'hE2; #100;
A = 8'h68; B = 8'hE3; #100;
A = 8'h68; B = 8'hE4; #100;
A = 8'h68; B = 8'hE5; #100;
A = 8'h68; B = 8'hE6; #100;
A = 8'h68; B = 8'hE7; #100;
A = 8'h68; B = 8'hE8; #100;
A = 8'h68; B = 8'hE9; #100;
A = 8'h68; B = 8'hEA; #100;
A = 8'h68; B = 8'hEB; #100;
A = 8'h68; B = 8'hEC; #100;
A = 8'h68; B = 8'hED; #100;
A = 8'h68; B = 8'hEE; #100;
A = 8'h68; B = 8'hEF; #100;
A = 8'h68; B = 8'hF0; #100;
A = 8'h68; B = 8'hF1; #100;
A = 8'h68; B = 8'hF2; #100;
A = 8'h68; B = 8'hF3; #100;
A = 8'h68; B = 8'hF4; #100;
A = 8'h68; B = 8'hF5; #100;
A = 8'h68; B = 8'hF6; #100;
A = 8'h68; B = 8'hF7; #100;
A = 8'h68; B = 8'hF8; #100;
A = 8'h68; B = 8'hF9; #100;
A = 8'h68; B = 8'hFA; #100;
A = 8'h68; B = 8'hFB; #100;
A = 8'h68; B = 8'hFC; #100;
A = 8'h68; B = 8'hFD; #100;
A = 8'h68; B = 8'hFE; #100;
A = 8'h68; B = 8'hFF; #100;
A = 8'h69; B = 8'h0; #100;
A = 8'h69; B = 8'h1; #100;
A = 8'h69; B = 8'h2; #100;
A = 8'h69; B = 8'h3; #100;
A = 8'h69; B = 8'h4; #100;
A = 8'h69; B = 8'h5; #100;
A = 8'h69; B = 8'h6; #100;
A = 8'h69; B = 8'h7; #100;
A = 8'h69; B = 8'h8; #100;
A = 8'h69; B = 8'h9; #100;
A = 8'h69; B = 8'hA; #100;
A = 8'h69; B = 8'hB; #100;
A = 8'h69; B = 8'hC; #100;
A = 8'h69; B = 8'hD; #100;
A = 8'h69; B = 8'hE; #100;
A = 8'h69; B = 8'hF; #100;
A = 8'h69; B = 8'h10; #100;
A = 8'h69; B = 8'h11; #100;
A = 8'h69; B = 8'h12; #100;
A = 8'h69; B = 8'h13; #100;
A = 8'h69; B = 8'h14; #100;
A = 8'h69; B = 8'h15; #100;
A = 8'h69; B = 8'h16; #100;
A = 8'h69; B = 8'h17; #100;
A = 8'h69; B = 8'h18; #100;
A = 8'h69; B = 8'h19; #100;
A = 8'h69; B = 8'h1A; #100;
A = 8'h69; B = 8'h1B; #100;
A = 8'h69; B = 8'h1C; #100;
A = 8'h69; B = 8'h1D; #100;
A = 8'h69; B = 8'h1E; #100;
A = 8'h69; B = 8'h1F; #100;
A = 8'h69; B = 8'h20; #100;
A = 8'h69; B = 8'h21; #100;
A = 8'h69; B = 8'h22; #100;
A = 8'h69; B = 8'h23; #100;
A = 8'h69; B = 8'h24; #100;
A = 8'h69; B = 8'h25; #100;
A = 8'h69; B = 8'h26; #100;
A = 8'h69; B = 8'h27; #100;
A = 8'h69; B = 8'h28; #100;
A = 8'h69; B = 8'h29; #100;
A = 8'h69; B = 8'h2A; #100;
A = 8'h69; B = 8'h2B; #100;
A = 8'h69; B = 8'h2C; #100;
A = 8'h69; B = 8'h2D; #100;
A = 8'h69; B = 8'h2E; #100;
A = 8'h69; B = 8'h2F; #100;
A = 8'h69; B = 8'h30; #100;
A = 8'h69; B = 8'h31; #100;
A = 8'h69; B = 8'h32; #100;
A = 8'h69; B = 8'h33; #100;
A = 8'h69; B = 8'h34; #100;
A = 8'h69; B = 8'h35; #100;
A = 8'h69; B = 8'h36; #100;
A = 8'h69; B = 8'h37; #100;
A = 8'h69; B = 8'h38; #100;
A = 8'h69; B = 8'h39; #100;
A = 8'h69; B = 8'h3A; #100;
A = 8'h69; B = 8'h3B; #100;
A = 8'h69; B = 8'h3C; #100;
A = 8'h69; B = 8'h3D; #100;
A = 8'h69; B = 8'h3E; #100;
A = 8'h69; B = 8'h3F; #100;
A = 8'h69; B = 8'h40; #100;
A = 8'h69; B = 8'h41; #100;
A = 8'h69; B = 8'h42; #100;
A = 8'h69; B = 8'h43; #100;
A = 8'h69; B = 8'h44; #100;
A = 8'h69; B = 8'h45; #100;
A = 8'h69; B = 8'h46; #100;
A = 8'h69; B = 8'h47; #100;
A = 8'h69; B = 8'h48; #100;
A = 8'h69; B = 8'h49; #100;
A = 8'h69; B = 8'h4A; #100;
A = 8'h69; B = 8'h4B; #100;
A = 8'h69; B = 8'h4C; #100;
A = 8'h69; B = 8'h4D; #100;
A = 8'h69; B = 8'h4E; #100;
A = 8'h69; B = 8'h4F; #100;
A = 8'h69; B = 8'h50; #100;
A = 8'h69; B = 8'h51; #100;
A = 8'h69; B = 8'h52; #100;
A = 8'h69; B = 8'h53; #100;
A = 8'h69; B = 8'h54; #100;
A = 8'h69; B = 8'h55; #100;
A = 8'h69; B = 8'h56; #100;
A = 8'h69; B = 8'h57; #100;
A = 8'h69; B = 8'h58; #100;
A = 8'h69; B = 8'h59; #100;
A = 8'h69; B = 8'h5A; #100;
A = 8'h69; B = 8'h5B; #100;
A = 8'h69; B = 8'h5C; #100;
A = 8'h69; B = 8'h5D; #100;
A = 8'h69; B = 8'h5E; #100;
A = 8'h69; B = 8'h5F; #100;
A = 8'h69; B = 8'h60; #100;
A = 8'h69; B = 8'h61; #100;
A = 8'h69; B = 8'h62; #100;
A = 8'h69; B = 8'h63; #100;
A = 8'h69; B = 8'h64; #100;
A = 8'h69; B = 8'h65; #100;
A = 8'h69; B = 8'h66; #100;
A = 8'h69; B = 8'h67; #100;
A = 8'h69; B = 8'h68; #100;
A = 8'h69; B = 8'h69; #100;
A = 8'h69; B = 8'h6A; #100;
A = 8'h69; B = 8'h6B; #100;
A = 8'h69; B = 8'h6C; #100;
A = 8'h69; B = 8'h6D; #100;
A = 8'h69; B = 8'h6E; #100;
A = 8'h69; B = 8'h6F; #100;
A = 8'h69; B = 8'h70; #100;
A = 8'h69; B = 8'h71; #100;
A = 8'h69; B = 8'h72; #100;
A = 8'h69; B = 8'h73; #100;
A = 8'h69; B = 8'h74; #100;
A = 8'h69; B = 8'h75; #100;
A = 8'h69; B = 8'h76; #100;
A = 8'h69; B = 8'h77; #100;
A = 8'h69; B = 8'h78; #100;
A = 8'h69; B = 8'h79; #100;
A = 8'h69; B = 8'h7A; #100;
A = 8'h69; B = 8'h7B; #100;
A = 8'h69; B = 8'h7C; #100;
A = 8'h69; B = 8'h7D; #100;
A = 8'h69; B = 8'h7E; #100;
A = 8'h69; B = 8'h7F; #100;
A = 8'h69; B = 8'h80; #100;
A = 8'h69; B = 8'h81; #100;
A = 8'h69; B = 8'h82; #100;
A = 8'h69; B = 8'h83; #100;
A = 8'h69; B = 8'h84; #100;
A = 8'h69; B = 8'h85; #100;
A = 8'h69; B = 8'h86; #100;
A = 8'h69; B = 8'h87; #100;
A = 8'h69; B = 8'h88; #100;
A = 8'h69; B = 8'h89; #100;
A = 8'h69; B = 8'h8A; #100;
A = 8'h69; B = 8'h8B; #100;
A = 8'h69; B = 8'h8C; #100;
A = 8'h69; B = 8'h8D; #100;
A = 8'h69; B = 8'h8E; #100;
A = 8'h69; B = 8'h8F; #100;
A = 8'h69; B = 8'h90; #100;
A = 8'h69; B = 8'h91; #100;
A = 8'h69; B = 8'h92; #100;
A = 8'h69; B = 8'h93; #100;
A = 8'h69; B = 8'h94; #100;
A = 8'h69; B = 8'h95; #100;
A = 8'h69; B = 8'h96; #100;
A = 8'h69; B = 8'h97; #100;
A = 8'h69; B = 8'h98; #100;
A = 8'h69; B = 8'h99; #100;
A = 8'h69; B = 8'h9A; #100;
A = 8'h69; B = 8'h9B; #100;
A = 8'h69; B = 8'h9C; #100;
A = 8'h69; B = 8'h9D; #100;
A = 8'h69; B = 8'h9E; #100;
A = 8'h69; B = 8'h9F; #100;
A = 8'h69; B = 8'hA0; #100;
A = 8'h69; B = 8'hA1; #100;
A = 8'h69; B = 8'hA2; #100;
A = 8'h69; B = 8'hA3; #100;
A = 8'h69; B = 8'hA4; #100;
A = 8'h69; B = 8'hA5; #100;
A = 8'h69; B = 8'hA6; #100;
A = 8'h69; B = 8'hA7; #100;
A = 8'h69; B = 8'hA8; #100;
A = 8'h69; B = 8'hA9; #100;
A = 8'h69; B = 8'hAA; #100;
A = 8'h69; B = 8'hAB; #100;
A = 8'h69; B = 8'hAC; #100;
A = 8'h69; B = 8'hAD; #100;
A = 8'h69; B = 8'hAE; #100;
A = 8'h69; B = 8'hAF; #100;
A = 8'h69; B = 8'hB0; #100;
A = 8'h69; B = 8'hB1; #100;
A = 8'h69; B = 8'hB2; #100;
A = 8'h69; B = 8'hB3; #100;
A = 8'h69; B = 8'hB4; #100;
A = 8'h69; B = 8'hB5; #100;
A = 8'h69; B = 8'hB6; #100;
A = 8'h69; B = 8'hB7; #100;
A = 8'h69; B = 8'hB8; #100;
A = 8'h69; B = 8'hB9; #100;
A = 8'h69; B = 8'hBA; #100;
A = 8'h69; B = 8'hBB; #100;
A = 8'h69; B = 8'hBC; #100;
A = 8'h69; B = 8'hBD; #100;
A = 8'h69; B = 8'hBE; #100;
A = 8'h69; B = 8'hBF; #100;
A = 8'h69; B = 8'hC0; #100;
A = 8'h69; B = 8'hC1; #100;
A = 8'h69; B = 8'hC2; #100;
A = 8'h69; B = 8'hC3; #100;
A = 8'h69; B = 8'hC4; #100;
A = 8'h69; B = 8'hC5; #100;
A = 8'h69; B = 8'hC6; #100;
A = 8'h69; B = 8'hC7; #100;
A = 8'h69; B = 8'hC8; #100;
A = 8'h69; B = 8'hC9; #100;
A = 8'h69; B = 8'hCA; #100;
A = 8'h69; B = 8'hCB; #100;
A = 8'h69; B = 8'hCC; #100;
A = 8'h69; B = 8'hCD; #100;
A = 8'h69; B = 8'hCE; #100;
A = 8'h69; B = 8'hCF; #100;
A = 8'h69; B = 8'hD0; #100;
A = 8'h69; B = 8'hD1; #100;
A = 8'h69; B = 8'hD2; #100;
A = 8'h69; B = 8'hD3; #100;
A = 8'h69; B = 8'hD4; #100;
A = 8'h69; B = 8'hD5; #100;
A = 8'h69; B = 8'hD6; #100;
A = 8'h69; B = 8'hD7; #100;
A = 8'h69; B = 8'hD8; #100;
A = 8'h69; B = 8'hD9; #100;
A = 8'h69; B = 8'hDA; #100;
A = 8'h69; B = 8'hDB; #100;
A = 8'h69; B = 8'hDC; #100;
A = 8'h69; B = 8'hDD; #100;
A = 8'h69; B = 8'hDE; #100;
A = 8'h69; B = 8'hDF; #100;
A = 8'h69; B = 8'hE0; #100;
A = 8'h69; B = 8'hE1; #100;
A = 8'h69; B = 8'hE2; #100;
A = 8'h69; B = 8'hE3; #100;
A = 8'h69; B = 8'hE4; #100;
A = 8'h69; B = 8'hE5; #100;
A = 8'h69; B = 8'hE6; #100;
A = 8'h69; B = 8'hE7; #100;
A = 8'h69; B = 8'hE8; #100;
A = 8'h69; B = 8'hE9; #100;
A = 8'h69; B = 8'hEA; #100;
A = 8'h69; B = 8'hEB; #100;
A = 8'h69; B = 8'hEC; #100;
A = 8'h69; B = 8'hED; #100;
A = 8'h69; B = 8'hEE; #100;
A = 8'h69; B = 8'hEF; #100;
A = 8'h69; B = 8'hF0; #100;
A = 8'h69; B = 8'hF1; #100;
A = 8'h69; B = 8'hF2; #100;
A = 8'h69; B = 8'hF3; #100;
A = 8'h69; B = 8'hF4; #100;
A = 8'h69; B = 8'hF5; #100;
A = 8'h69; B = 8'hF6; #100;
A = 8'h69; B = 8'hF7; #100;
A = 8'h69; B = 8'hF8; #100;
A = 8'h69; B = 8'hF9; #100;
A = 8'h69; B = 8'hFA; #100;
A = 8'h69; B = 8'hFB; #100;
A = 8'h69; B = 8'hFC; #100;
A = 8'h69; B = 8'hFD; #100;
A = 8'h69; B = 8'hFE; #100;
A = 8'h69; B = 8'hFF; #100;
A = 8'h6A; B = 8'h0; #100;
A = 8'h6A; B = 8'h1; #100;
A = 8'h6A; B = 8'h2; #100;
A = 8'h6A; B = 8'h3; #100;
A = 8'h6A; B = 8'h4; #100;
A = 8'h6A; B = 8'h5; #100;
A = 8'h6A; B = 8'h6; #100;
A = 8'h6A; B = 8'h7; #100;
A = 8'h6A; B = 8'h8; #100;
A = 8'h6A; B = 8'h9; #100;
A = 8'h6A; B = 8'hA; #100;
A = 8'h6A; B = 8'hB; #100;
A = 8'h6A; B = 8'hC; #100;
A = 8'h6A; B = 8'hD; #100;
A = 8'h6A; B = 8'hE; #100;
A = 8'h6A; B = 8'hF; #100;
A = 8'h6A; B = 8'h10; #100;
A = 8'h6A; B = 8'h11; #100;
A = 8'h6A; B = 8'h12; #100;
A = 8'h6A; B = 8'h13; #100;
A = 8'h6A; B = 8'h14; #100;
A = 8'h6A; B = 8'h15; #100;
A = 8'h6A; B = 8'h16; #100;
A = 8'h6A; B = 8'h17; #100;
A = 8'h6A; B = 8'h18; #100;
A = 8'h6A; B = 8'h19; #100;
A = 8'h6A; B = 8'h1A; #100;
A = 8'h6A; B = 8'h1B; #100;
A = 8'h6A; B = 8'h1C; #100;
A = 8'h6A; B = 8'h1D; #100;
A = 8'h6A; B = 8'h1E; #100;
A = 8'h6A; B = 8'h1F; #100;
A = 8'h6A; B = 8'h20; #100;
A = 8'h6A; B = 8'h21; #100;
A = 8'h6A; B = 8'h22; #100;
A = 8'h6A; B = 8'h23; #100;
A = 8'h6A; B = 8'h24; #100;
A = 8'h6A; B = 8'h25; #100;
A = 8'h6A; B = 8'h26; #100;
A = 8'h6A; B = 8'h27; #100;
A = 8'h6A; B = 8'h28; #100;
A = 8'h6A; B = 8'h29; #100;
A = 8'h6A; B = 8'h2A; #100;
A = 8'h6A; B = 8'h2B; #100;
A = 8'h6A; B = 8'h2C; #100;
A = 8'h6A; B = 8'h2D; #100;
A = 8'h6A; B = 8'h2E; #100;
A = 8'h6A; B = 8'h2F; #100;
A = 8'h6A; B = 8'h30; #100;
A = 8'h6A; B = 8'h31; #100;
A = 8'h6A; B = 8'h32; #100;
A = 8'h6A; B = 8'h33; #100;
A = 8'h6A; B = 8'h34; #100;
A = 8'h6A; B = 8'h35; #100;
A = 8'h6A; B = 8'h36; #100;
A = 8'h6A; B = 8'h37; #100;
A = 8'h6A; B = 8'h38; #100;
A = 8'h6A; B = 8'h39; #100;
A = 8'h6A; B = 8'h3A; #100;
A = 8'h6A; B = 8'h3B; #100;
A = 8'h6A; B = 8'h3C; #100;
A = 8'h6A; B = 8'h3D; #100;
A = 8'h6A; B = 8'h3E; #100;
A = 8'h6A; B = 8'h3F; #100;
A = 8'h6A; B = 8'h40; #100;
A = 8'h6A; B = 8'h41; #100;
A = 8'h6A; B = 8'h42; #100;
A = 8'h6A; B = 8'h43; #100;
A = 8'h6A; B = 8'h44; #100;
A = 8'h6A; B = 8'h45; #100;
A = 8'h6A; B = 8'h46; #100;
A = 8'h6A; B = 8'h47; #100;
A = 8'h6A; B = 8'h48; #100;
A = 8'h6A; B = 8'h49; #100;
A = 8'h6A; B = 8'h4A; #100;
A = 8'h6A; B = 8'h4B; #100;
A = 8'h6A; B = 8'h4C; #100;
A = 8'h6A; B = 8'h4D; #100;
A = 8'h6A; B = 8'h4E; #100;
A = 8'h6A; B = 8'h4F; #100;
A = 8'h6A; B = 8'h50; #100;
A = 8'h6A; B = 8'h51; #100;
A = 8'h6A; B = 8'h52; #100;
A = 8'h6A; B = 8'h53; #100;
A = 8'h6A; B = 8'h54; #100;
A = 8'h6A; B = 8'h55; #100;
A = 8'h6A; B = 8'h56; #100;
A = 8'h6A; B = 8'h57; #100;
A = 8'h6A; B = 8'h58; #100;
A = 8'h6A; B = 8'h59; #100;
A = 8'h6A; B = 8'h5A; #100;
A = 8'h6A; B = 8'h5B; #100;
A = 8'h6A; B = 8'h5C; #100;
A = 8'h6A; B = 8'h5D; #100;
A = 8'h6A; B = 8'h5E; #100;
A = 8'h6A; B = 8'h5F; #100;
A = 8'h6A; B = 8'h60; #100;
A = 8'h6A; B = 8'h61; #100;
A = 8'h6A; B = 8'h62; #100;
A = 8'h6A; B = 8'h63; #100;
A = 8'h6A; B = 8'h64; #100;
A = 8'h6A; B = 8'h65; #100;
A = 8'h6A; B = 8'h66; #100;
A = 8'h6A; B = 8'h67; #100;
A = 8'h6A; B = 8'h68; #100;
A = 8'h6A; B = 8'h69; #100;
A = 8'h6A; B = 8'h6A; #100;
A = 8'h6A; B = 8'h6B; #100;
A = 8'h6A; B = 8'h6C; #100;
A = 8'h6A; B = 8'h6D; #100;
A = 8'h6A; B = 8'h6E; #100;
A = 8'h6A; B = 8'h6F; #100;
A = 8'h6A; B = 8'h70; #100;
A = 8'h6A; B = 8'h71; #100;
A = 8'h6A; B = 8'h72; #100;
A = 8'h6A; B = 8'h73; #100;
A = 8'h6A; B = 8'h74; #100;
A = 8'h6A; B = 8'h75; #100;
A = 8'h6A; B = 8'h76; #100;
A = 8'h6A; B = 8'h77; #100;
A = 8'h6A; B = 8'h78; #100;
A = 8'h6A; B = 8'h79; #100;
A = 8'h6A; B = 8'h7A; #100;
A = 8'h6A; B = 8'h7B; #100;
A = 8'h6A; B = 8'h7C; #100;
A = 8'h6A; B = 8'h7D; #100;
A = 8'h6A; B = 8'h7E; #100;
A = 8'h6A; B = 8'h7F; #100;
A = 8'h6A; B = 8'h80; #100;
A = 8'h6A; B = 8'h81; #100;
A = 8'h6A; B = 8'h82; #100;
A = 8'h6A; B = 8'h83; #100;
A = 8'h6A; B = 8'h84; #100;
A = 8'h6A; B = 8'h85; #100;
A = 8'h6A; B = 8'h86; #100;
A = 8'h6A; B = 8'h87; #100;
A = 8'h6A; B = 8'h88; #100;
A = 8'h6A; B = 8'h89; #100;
A = 8'h6A; B = 8'h8A; #100;
A = 8'h6A; B = 8'h8B; #100;
A = 8'h6A; B = 8'h8C; #100;
A = 8'h6A; B = 8'h8D; #100;
A = 8'h6A; B = 8'h8E; #100;
A = 8'h6A; B = 8'h8F; #100;
A = 8'h6A; B = 8'h90; #100;
A = 8'h6A; B = 8'h91; #100;
A = 8'h6A; B = 8'h92; #100;
A = 8'h6A; B = 8'h93; #100;
A = 8'h6A; B = 8'h94; #100;
A = 8'h6A; B = 8'h95; #100;
A = 8'h6A; B = 8'h96; #100;
A = 8'h6A; B = 8'h97; #100;
A = 8'h6A; B = 8'h98; #100;
A = 8'h6A; B = 8'h99; #100;
A = 8'h6A; B = 8'h9A; #100;
A = 8'h6A; B = 8'h9B; #100;
A = 8'h6A; B = 8'h9C; #100;
A = 8'h6A; B = 8'h9D; #100;
A = 8'h6A; B = 8'h9E; #100;
A = 8'h6A; B = 8'h9F; #100;
A = 8'h6A; B = 8'hA0; #100;
A = 8'h6A; B = 8'hA1; #100;
A = 8'h6A; B = 8'hA2; #100;
A = 8'h6A; B = 8'hA3; #100;
A = 8'h6A; B = 8'hA4; #100;
A = 8'h6A; B = 8'hA5; #100;
A = 8'h6A; B = 8'hA6; #100;
A = 8'h6A; B = 8'hA7; #100;
A = 8'h6A; B = 8'hA8; #100;
A = 8'h6A; B = 8'hA9; #100;
A = 8'h6A; B = 8'hAA; #100;
A = 8'h6A; B = 8'hAB; #100;
A = 8'h6A; B = 8'hAC; #100;
A = 8'h6A; B = 8'hAD; #100;
A = 8'h6A; B = 8'hAE; #100;
A = 8'h6A; B = 8'hAF; #100;
A = 8'h6A; B = 8'hB0; #100;
A = 8'h6A; B = 8'hB1; #100;
A = 8'h6A; B = 8'hB2; #100;
A = 8'h6A; B = 8'hB3; #100;
A = 8'h6A; B = 8'hB4; #100;
A = 8'h6A; B = 8'hB5; #100;
A = 8'h6A; B = 8'hB6; #100;
A = 8'h6A; B = 8'hB7; #100;
A = 8'h6A; B = 8'hB8; #100;
A = 8'h6A; B = 8'hB9; #100;
A = 8'h6A; B = 8'hBA; #100;
A = 8'h6A; B = 8'hBB; #100;
A = 8'h6A; B = 8'hBC; #100;
A = 8'h6A; B = 8'hBD; #100;
A = 8'h6A; B = 8'hBE; #100;
A = 8'h6A; B = 8'hBF; #100;
A = 8'h6A; B = 8'hC0; #100;
A = 8'h6A; B = 8'hC1; #100;
A = 8'h6A; B = 8'hC2; #100;
A = 8'h6A; B = 8'hC3; #100;
A = 8'h6A; B = 8'hC4; #100;
A = 8'h6A; B = 8'hC5; #100;
A = 8'h6A; B = 8'hC6; #100;
A = 8'h6A; B = 8'hC7; #100;
A = 8'h6A; B = 8'hC8; #100;
A = 8'h6A; B = 8'hC9; #100;
A = 8'h6A; B = 8'hCA; #100;
A = 8'h6A; B = 8'hCB; #100;
A = 8'h6A; B = 8'hCC; #100;
A = 8'h6A; B = 8'hCD; #100;
A = 8'h6A; B = 8'hCE; #100;
A = 8'h6A; B = 8'hCF; #100;
A = 8'h6A; B = 8'hD0; #100;
A = 8'h6A; B = 8'hD1; #100;
A = 8'h6A; B = 8'hD2; #100;
A = 8'h6A; B = 8'hD3; #100;
A = 8'h6A; B = 8'hD4; #100;
A = 8'h6A; B = 8'hD5; #100;
A = 8'h6A; B = 8'hD6; #100;
A = 8'h6A; B = 8'hD7; #100;
A = 8'h6A; B = 8'hD8; #100;
A = 8'h6A; B = 8'hD9; #100;
A = 8'h6A; B = 8'hDA; #100;
A = 8'h6A; B = 8'hDB; #100;
A = 8'h6A; B = 8'hDC; #100;
A = 8'h6A; B = 8'hDD; #100;
A = 8'h6A; B = 8'hDE; #100;
A = 8'h6A; B = 8'hDF; #100;
A = 8'h6A; B = 8'hE0; #100;
A = 8'h6A; B = 8'hE1; #100;
A = 8'h6A; B = 8'hE2; #100;
A = 8'h6A; B = 8'hE3; #100;
A = 8'h6A; B = 8'hE4; #100;
A = 8'h6A; B = 8'hE5; #100;
A = 8'h6A; B = 8'hE6; #100;
A = 8'h6A; B = 8'hE7; #100;
A = 8'h6A; B = 8'hE8; #100;
A = 8'h6A; B = 8'hE9; #100;
A = 8'h6A; B = 8'hEA; #100;
A = 8'h6A; B = 8'hEB; #100;
A = 8'h6A; B = 8'hEC; #100;
A = 8'h6A; B = 8'hED; #100;
A = 8'h6A; B = 8'hEE; #100;
A = 8'h6A; B = 8'hEF; #100;
A = 8'h6A; B = 8'hF0; #100;
A = 8'h6A; B = 8'hF1; #100;
A = 8'h6A; B = 8'hF2; #100;
A = 8'h6A; B = 8'hF3; #100;
A = 8'h6A; B = 8'hF4; #100;
A = 8'h6A; B = 8'hF5; #100;
A = 8'h6A; B = 8'hF6; #100;
A = 8'h6A; B = 8'hF7; #100;
A = 8'h6A; B = 8'hF8; #100;
A = 8'h6A; B = 8'hF9; #100;
A = 8'h6A; B = 8'hFA; #100;
A = 8'h6A; B = 8'hFB; #100;
A = 8'h6A; B = 8'hFC; #100;
A = 8'h6A; B = 8'hFD; #100;
A = 8'h6A; B = 8'hFE; #100;
A = 8'h6A; B = 8'hFF; #100;
A = 8'h6B; B = 8'h0; #100;
A = 8'h6B; B = 8'h1; #100;
A = 8'h6B; B = 8'h2; #100;
A = 8'h6B; B = 8'h3; #100;
A = 8'h6B; B = 8'h4; #100;
A = 8'h6B; B = 8'h5; #100;
A = 8'h6B; B = 8'h6; #100;
A = 8'h6B; B = 8'h7; #100;
A = 8'h6B; B = 8'h8; #100;
A = 8'h6B; B = 8'h9; #100;
A = 8'h6B; B = 8'hA; #100;
A = 8'h6B; B = 8'hB; #100;
A = 8'h6B; B = 8'hC; #100;
A = 8'h6B; B = 8'hD; #100;
A = 8'h6B; B = 8'hE; #100;
A = 8'h6B; B = 8'hF; #100;
A = 8'h6B; B = 8'h10; #100;
A = 8'h6B; B = 8'h11; #100;
A = 8'h6B; B = 8'h12; #100;
A = 8'h6B; B = 8'h13; #100;
A = 8'h6B; B = 8'h14; #100;
A = 8'h6B; B = 8'h15; #100;
A = 8'h6B; B = 8'h16; #100;
A = 8'h6B; B = 8'h17; #100;
A = 8'h6B; B = 8'h18; #100;
A = 8'h6B; B = 8'h19; #100;
A = 8'h6B; B = 8'h1A; #100;
A = 8'h6B; B = 8'h1B; #100;
A = 8'h6B; B = 8'h1C; #100;
A = 8'h6B; B = 8'h1D; #100;
A = 8'h6B; B = 8'h1E; #100;
A = 8'h6B; B = 8'h1F; #100;
A = 8'h6B; B = 8'h20; #100;
A = 8'h6B; B = 8'h21; #100;
A = 8'h6B; B = 8'h22; #100;
A = 8'h6B; B = 8'h23; #100;
A = 8'h6B; B = 8'h24; #100;
A = 8'h6B; B = 8'h25; #100;
A = 8'h6B; B = 8'h26; #100;
A = 8'h6B; B = 8'h27; #100;
A = 8'h6B; B = 8'h28; #100;
A = 8'h6B; B = 8'h29; #100;
A = 8'h6B; B = 8'h2A; #100;
A = 8'h6B; B = 8'h2B; #100;
A = 8'h6B; B = 8'h2C; #100;
A = 8'h6B; B = 8'h2D; #100;
A = 8'h6B; B = 8'h2E; #100;
A = 8'h6B; B = 8'h2F; #100;
A = 8'h6B; B = 8'h30; #100;
A = 8'h6B; B = 8'h31; #100;
A = 8'h6B; B = 8'h32; #100;
A = 8'h6B; B = 8'h33; #100;
A = 8'h6B; B = 8'h34; #100;
A = 8'h6B; B = 8'h35; #100;
A = 8'h6B; B = 8'h36; #100;
A = 8'h6B; B = 8'h37; #100;
A = 8'h6B; B = 8'h38; #100;
A = 8'h6B; B = 8'h39; #100;
A = 8'h6B; B = 8'h3A; #100;
A = 8'h6B; B = 8'h3B; #100;
A = 8'h6B; B = 8'h3C; #100;
A = 8'h6B; B = 8'h3D; #100;
A = 8'h6B; B = 8'h3E; #100;
A = 8'h6B; B = 8'h3F; #100;
A = 8'h6B; B = 8'h40; #100;
A = 8'h6B; B = 8'h41; #100;
A = 8'h6B; B = 8'h42; #100;
A = 8'h6B; B = 8'h43; #100;
A = 8'h6B; B = 8'h44; #100;
A = 8'h6B; B = 8'h45; #100;
A = 8'h6B; B = 8'h46; #100;
A = 8'h6B; B = 8'h47; #100;
A = 8'h6B; B = 8'h48; #100;
A = 8'h6B; B = 8'h49; #100;
A = 8'h6B; B = 8'h4A; #100;
A = 8'h6B; B = 8'h4B; #100;
A = 8'h6B; B = 8'h4C; #100;
A = 8'h6B; B = 8'h4D; #100;
A = 8'h6B; B = 8'h4E; #100;
A = 8'h6B; B = 8'h4F; #100;
A = 8'h6B; B = 8'h50; #100;
A = 8'h6B; B = 8'h51; #100;
A = 8'h6B; B = 8'h52; #100;
A = 8'h6B; B = 8'h53; #100;
A = 8'h6B; B = 8'h54; #100;
A = 8'h6B; B = 8'h55; #100;
A = 8'h6B; B = 8'h56; #100;
A = 8'h6B; B = 8'h57; #100;
A = 8'h6B; B = 8'h58; #100;
A = 8'h6B; B = 8'h59; #100;
A = 8'h6B; B = 8'h5A; #100;
A = 8'h6B; B = 8'h5B; #100;
A = 8'h6B; B = 8'h5C; #100;
A = 8'h6B; B = 8'h5D; #100;
A = 8'h6B; B = 8'h5E; #100;
A = 8'h6B; B = 8'h5F; #100;
A = 8'h6B; B = 8'h60; #100;
A = 8'h6B; B = 8'h61; #100;
A = 8'h6B; B = 8'h62; #100;
A = 8'h6B; B = 8'h63; #100;
A = 8'h6B; B = 8'h64; #100;
A = 8'h6B; B = 8'h65; #100;
A = 8'h6B; B = 8'h66; #100;
A = 8'h6B; B = 8'h67; #100;
A = 8'h6B; B = 8'h68; #100;
A = 8'h6B; B = 8'h69; #100;
A = 8'h6B; B = 8'h6A; #100;
A = 8'h6B; B = 8'h6B; #100;
A = 8'h6B; B = 8'h6C; #100;
A = 8'h6B; B = 8'h6D; #100;
A = 8'h6B; B = 8'h6E; #100;
A = 8'h6B; B = 8'h6F; #100;
A = 8'h6B; B = 8'h70; #100;
A = 8'h6B; B = 8'h71; #100;
A = 8'h6B; B = 8'h72; #100;
A = 8'h6B; B = 8'h73; #100;
A = 8'h6B; B = 8'h74; #100;
A = 8'h6B; B = 8'h75; #100;
A = 8'h6B; B = 8'h76; #100;
A = 8'h6B; B = 8'h77; #100;
A = 8'h6B; B = 8'h78; #100;
A = 8'h6B; B = 8'h79; #100;
A = 8'h6B; B = 8'h7A; #100;
A = 8'h6B; B = 8'h7B; #100;
A = 8'h6B; B = 8'h7C; #100;
A = 8'h6B; B = 8'h7D; #100;
A = 8'h6B; B = 8'h7E; #100;
A = 8'h6B; B = 8'h7F; #100;
A = 8'h6B; B = 8'h80; #100;
A = 8'h6B; B = 8'h81; #100;
A = 8'h6B; B = 8'h82; #100;
A = 8'h6B; B = 8'h83; #100;
A = 8'h6B; B = 8'h84; #100;
A = 8'h6B; B = 8'h85; #100;
A = 8'h6B; B = 8'h86; #100;
A = 8'h6B; B = 8'h87; #100;
A = 8'h6B; B = 8'h88; #100;
A = 8'h6B; B = 8'h89; #100;
A = 8'h6B; B = 8'h8A; #100;
A = 8'h6B; B = 8'h8B; #100;
A = 8'h6B; B = 8'h8C; #100;
A = 8'h6B; B = 8'h8D; #100;
A = 8'h6B; B = 8'h8E; #100;
A = 8'h6B; B = 8'h8F; #100;
A = 8'h6B; B = 8'h90; #100;
A = 8'h6B; B = 8'h91; #100;
A = 8'h6B; B = 8'h92; #100;
A = 8'h6B; B = 8'h93; #100;
A = 8'h6B; B = 8'h94; #100;
A = 8'h6B; B = 8'h95; #100;
A = 8'h6B; B = 8'h96; #100;
A = 8'h6B; B = 8'h97; #100;
A = 8'h6B; B = 8'h98; #100;
A = 8'h6B; B = 8'h99; #100;
A = 8'h6B; B = 8'h9A; #100;
A = 8'h6B; B = 8'h9B; #100;
A = 8'h6B; B = 8'h9C; #100;
A = 8'h6B; B = 8'h9D; #100;
A = 8'h6B; B = 8'h9E; #100;
A = 8'h6B; B = 8'h9F; #100;
A = 8'h6B; B = 8'hA0; #100;
A = 8'h6B; B = 8'hA1; #100;
A = 8'h6B; B = 8'hA2; #100;
A = 8'h6B; B = 8'hA3; #100;
A = 8'h6B; B = 8'hA4; #100;
A = 8'h6B; B = 8'hA5; #100;
A = 8'h6B; B = 8'hA6; #100;
A = 8'h6B; B = 8'hA7; #100;
A = 8'h6B; B = 8'hA8; #100;
A = 8'h6B; B = 8'hA9; #100;
A = 8'h6B; B = 8'hAA; #100;
A = 8'h6B; B = 8'hAB; #100;
A = 8'h6B; B = 8'hAC; #100;
A = 8'h6B; B = 8'hAD; #100;
A = 8'h6B; B = 8'hAE; #100;
A = 8'h6B; B = 8'hAF; #100;
A = 8'h6B; B = 8'hB0; #100;
A = 8'h6B; B = 8'hB1; #100;
A = 8'h6B; B = 8'hB2; #100;
A = 8'h6B; B = 8'hB3; #100;
A = 8'h6B; B = 8'hB4; #100;
A = 8'h6B; B = 8'hB5; #100;
A = 8'h6B; B = 8'hB6; #100;
A = 8'h6B; B = 8'hB7; #100;
A = 8'h6B; B = 8'hB8; #100;
A = 8'h6B; B = 8'hB9; #100;
A = 8'h6B; B = 8'hBA; #100;
A = 8'h6B; B = 8'hBB; #100;
A = 8'h6B; B = 8'hBC; #100;
A = 8'h6B; B = 8'hBD; #100;
A = 8'h6B; B = 8'hBE; #100;
A = 8'h6B; B = 8'hBF; #100;
A = 8'h6B; B = 8'hC0; #100;
A = 8'h6B; B = 8'hC1; #100;
A = 8'h6B; B = 8'hC2; #100;
A = 8'h6B; B = 8'hC3; #100;
A = 8'h6B; B = 8'hC4; #100;
A = 8'h6B; B = 8'hC5; #100;
A = 8'h6B; B = 8'hC6; #100;
A = 8'h6B; B = 8'hC7; #100;
A = 8'h6B; B = 8'hC8; #100;
A = 8'h6B; B = 8'hC9; #100;
A = 8'h6B; B = 8'hCA; #100;
A = 8'h6B; B = 8'hCB; #100;
A = 8'h6B; B = 8'hCC; #100;
A = 8'h6B; B = 8'hCD; #100;
A = 8'h6B; B = 8'hCE; #100;
A = 8'h6B; B = 8'hCF; #100;
A = 8'h6B; B = 8'hD0; #100;
A = 8'h6B; B = 8'hD1; #100;
A = 8'h6B; B = 8'hD2; #100;
A = 8'h6B; B = 8'hD3; #100;
A = 8'h6B; B = 8'hD4; #100;
A = 8'h6B; B = 8'hD5; #100;
A = 8'h6B; B = 8'hD6; #100;
A = 8'h6B; B = 8'hD7; #100;
A = 8'h6B; B = 8'hD8; #100;
A = 8'h6B; B = 8'hD9; #100;
A = 8'h6B; B = 8'hDA; #100;
A = 8'h6B; B = 8'hDB; #100;
A = 8'h6B; B = 8'hDC; #100;
A = 8'h6B; B = 8'hDD; #100;
A = 8'h6B; B = 8'hDE; #100;
A = 8'h6B; B = 8'hDF; #100;
A = 8'h6B; B = 8'hE0; #100;
A = 8'h6B; B = 8'hE1; #100;
A = 8'h6B; B = 8'hE2; #100;
A = 8'h6B; B = 8'hE3; #100;
A = 8'h6B; B = 8'hE4; #100;
A = 8'h6B; B = 8'hE5; #100;
A = 8'h6B; B = 8'hE6; #100;
A = 8'h6B; B = 8'hE7; #100;
A = 8'h6B; B = 8'hE8; #100;
A = 8'h6B; B = 8'hE9; #100;
A = 8'h6B; B = 8'hEA; #100;
A = 8'h6B; B = 8'hEB; #100;
A = 8'h6B; B = 8'hEC; #100;
A = 8'h6B; B = 8'hED; #100;
A = 8'h6B; B = 8'hEE; #100;
A = 8'h6B; B = 8'hEF; #100;
A = 8'h6B; B = 8'hF0; #100;
A = 8'h6B; B = 8'hF1; #100;
A = 8'h6B; B = 8'hF2; #100;
A = 8'h6B; B = 8'hF3; #100;
A = 8'h6B; B = 8'hF4; #100;
A = 8'h6B; B = 8'hF5; #100;
A = 8'h6B; B = 8'hF6; #100;
A = 8'h6B; B = 8'hF7; #100;
A = 8'h6B; B = 8'hF8; #100;
A = 8'h6B; B = 8'hF9; #100;
A = 8'h6B; B = 8'hFA; #100;
A = 8'h6B; B = 8'hFB; #100;
A = 8'h6B; B = 8'hFC; #100;
A = 8'h6B; B = 8'hFD; #100;
A = 8'h6B; B = 8'hFE; #100;
A = 8'h6B; B = 8'hFF; #100;
A = 8'h6C; B = 8'h0; #100;
A = 8'h6C; B = 8'h1; #100;
A = 8'h6C; B = 8'h2; #100;
A = 8'h6C; B = 8'h3; #100;
A = 8'h6C; B = 8'h4; #100;
A = 8'h6C; B = 8'h5; #100;
A = 8'h6C; B = 8'h6; #100;
A = 8'h6C; B = 8'h7; #100;
A = 8'h6C; B = 8'h8; #100;
A = 8'h6C; B = 8'h9; #100;
A = 8'h6C; B = 8'hA; #100;
A = 8'h6C; B = 8'hB; #100;
A = 8'h6C; B = 8'hC; #100;
A = 8'h6C; B = 8'hD; #100;
A = 8'h6C; B = 8'hE; #100;
A = 8'h6C; B = 8'hF; #100;
A = 8'h6C; B = 8'h10; #100;
A = 8'h6C; B = 8'h11; #100;
A = 8'h6C; B = 8'h12; #100;
A = 8'h6C; B = 8'h13; #100;
A = 8'h6C; B = 8'h14; #100;
A = 8'h6C; B = 8'h15; #100;
A = 8'h6C; B = 8'h16; #100;
A = 8'h6C; B = 8'h17; #100;
A = 8'h6C; B = 8'h18; #100;
A = 8'h6C; B = 8'h19; #100;
A = 8'h6C; B = 8'h1A; #100;
A = 8'h6C; B = 8'h1B; #100;
A = 8'h6C; B = 8'h1C; #100;
A = 8'h6C; B = 8'h1D; #100;
A = 8'h6C; B = 8'h1E; #100;
A = 8'h6C; B = 8'h1F; #100;
A = 8'h6C; B = 8'h20; #100;
A = 8'h6C; B = 8'h21; #100;
A = 8'h6C; B = 8'h22; #100;
A = 8'h6C; B = 8'h23; #100;
A = 8'h6C; B = 8'h24; #100;
A = 8'h6C; B = 8'h25; #100;
A = 8'h6C; B = 8'h26; #100;
A = 8'h6C; B = 8'h27; #100;
A = 8'h6C; B = 8'h28; #100;
A = 8'h6C; B = 8'h29; #100;
A = 8'h6C; B = 8'h2A; #100;
A = 8'h6C; B = 8'h2B; #100;
A = 8'h6C; B = 8'h2C; #100;
A = 8'h6C; B = 8'h2D; #100;
A = 8'h6C; B = 8'h2E; #100;
A = 8'h6C; B = 8'h2F; #100;
A = 8'h6C; B = 8'h30; #100;
A = 8'h6C; B = 8'h31; #100;
A = 8'h6C; B = 8'h32; #100;
A = 8'h6C; B = 8'h33; #100;
A = 8'h6C; B = 8'h34; #100;
A = 8'h6C; B = 8'h35; #100;
A = 8'h6C; B = 8'h36; #100;
A = 8'h6C; B = 8'h37; #100;
A = 8'h6C; B = 8'h38; #100;
A = 8'h6C; B = 8'h39; #100;
A = 8'h6C; B = 8'h3A; #100;
A = 8'h6C; B = 8'h3B; #100;
A = 8'h6C; B = 8'h3C; #100;
A = 8'h6C; B = 8'h3D; #100;
A = 8'h6C; B = 8'h3E; #100;
A = 8'h6C; B = 8'h3F; #100;
A = 8'h6C; B = 8'h40; #100;
A = 8'h6C; B = 8'h41; #100;
A = 8'h6C; B = 8'h42; #100;
A = 8'h6C; B = 8'h43; #100;
A = 8'h6C; B = 8'h44; #100;
A = 8'h6C; B = 8'h45; #100;
A = 8'h6C; B = 8'h46; #100;
A = 8'h6C; B = 8'h47; #100;
A = 8'h6C; B = 8'h48; #100;
A = 8'h6C; B = 8'h49; #100;
A = 8'h6C; B = 8'h4A; #100;
A = 8'h6C; B = 8'h4B; #100;
A = 8'h6C; B = 8'h4C; #100;
A = 8'h6C; B = 8'h4D; #100;
A = 8'h6C; B = 8'h4E; #100;
A = 8'h6C; B = 8'h4F; #100;
A = 8'h6C; B = 8'h50; #100;
A = 8'h6C; B = 8'h51; #100;
A = 8'h6C; B = 8'h52; #100;
A = 8'h6C; B = 8'h53; #100;
A = 8'h6C; B = 8'h54; #100;
A = 8'h6C; B = 8'h55; #100;
A = 8'h6C; B = 8'h56; #100;
A = 8'h6C; B = 8'h57; #100;
A = 8'h6C; B = 8'h58; #100;
A = 8'h6C; B = 8'h59; #100;
A = 8'h6C; B = 8'h5A; #100;
A = 8'h6C; B = 8'h5B; #100;
A = 8'h6C; B = 8'h5C; #100;
A = 8'h6C; B = 8'h5D; #100;
A = 8'h6C; B = 8'h5E; #100;
A = 8'h6C; B = 8'h5F; #100;
A = 8'h6C; B = 8'h60; #100;
A = 8'h6C; B = 8'h61; #100;
A = 8'h6C; B = 8'h62; #100;
A = 8'h6C; B = 8'h63; #100;
A = 8'h6C; B = 8'h64; #100;
A = 8'h6C; B = 8'h65; #100;
A = 8'h6C; B = 8'h66; #100;
A = 8'h6C; B = 8'h67; #100;
A = 8'h6C; B = 8'h68; #100;
A = 8'h6C; B = 8'h69; #100;
A = 8'h6C; B = 8'h6A; #100;
A = 8'h6C; B = 8'h6B; #100;
A = 8'h6C; B = 8'h6C; #100;
A = 8'h6C; B = 8'h6D; #100;
A = 8'h6C; B = 8'h6E; #100;
A = 8'h6C; B = 8'h6F; #100;
A = 8'h6C; B = 8'h70; #100;
A = 8'h6C; B = 8'h71; #100;
A = 8'h6C; B = 8'h72; #100;
A = 8'h6C; B = 8'h73; #100;
A = 8'h6C; B = 8'h74; #100;
A = 8'h6C; B = 8'h75; #100;
A = 8'h6C; B = 8'h76; #100;
A = 8'h6C; B = 8'h77; #100;
A = 8'h6C; B = 8'h78; #100;
A = 8'h6C; B = 8'h79; #100;
A = 8'h6C; B = 8'h7A; #100;
A = 8'h6C; B = 8'h7B; #100;
A = 8'h6C; B = 8'h7C; #100;
A = 8'h6C; B = 8'h7D; #100;
A = 8'h6C; B = 8'h7E; #100;
A = 8'h6C; B = 8'h7F; #100;
A = 8'h6C; B = 8'h80; #100;
A = 8'h6C; B = 8'h81; #100;
A = 8'h6C; B = 8'h82; #100;
A = 8'h6C; B = 8'h83; #100;
A = 8'h6C; B = 8'h84; #100;
A = 8'h6C; B = 8'h85; #100;
A = 8'h6C; B = 8'h86; #100;
A = 8'h6C; B = 8'h87; #100;
A = 8'h6C; B = 8'h88; #100;
A = 8'h6C; B = 8'h89; #100;
A = 8'h6C; B = 8'h8A; #100;
A = 8'h6C; B = 8'h8B; #100;
A = 8'h6C; B = 8'h8C; #100;
A = 8'h6C; B = 8'h8D; #100;
A = 8'h6C; B = 8'h8E; #100;
A = 8'h6C; B = 8'h8F; #100;
A = 8'h6C; B = 8'h90; #100;
A = 8'h6C; B = 8'h91; #100;
A = 8'h6C; B = 8'h92; #100;
A = 8'h6C; B = 8'h93; #100;
A = 8'h6C; B = 8'h94; #100;
A = 8'h6C; B = 8'h95; #100;
A = 8'h6C; B = 8'h96; #100;
A = 8'h6C; B = 8'h97; #100;
A = 8'h6C; B = 8'h98; #100;
A = 8'h6C; B = 8'h99; #100;
A = 8'h6C; B = 8'h9A; #100;
A = 8'h6C; B = 8'h9B; #100;
A = 8'h6C; B = 8'h9C; #100;
A = 8'h6C; B = 8'h9D; #100;
A = 8'h6C; B = 8'h9E; #100;
A = 8'h6C; B = 8'h9F; #100;
A = 8'h6C; B = 8'hA0; #100;
A = 8'h6C; B = 8'hA1; #100;
A = 8'h6C; B = 8'hA2; #100;
A = 8'h6C; B = 8'hA3; #100;
A = 8'h6C; B = 8'hA4; #100;
A = 8'h6C; B = 8'hA5; #100;
A = 8'h6C; B = 8'hA6; #100;
A = 8'h6C; B = 8'hA7; #100;
A = 8'h6C; B = 8'hA8; #100;
A = 8'h6C; B = 8'hA9; #100;
A = 8'h6C; B = 8'hAA; #100;
A = 8'h6C; B = 8'hAB; #100;
A = 8'h6C; B = 8'hAC; #100;
A = 8'h6C; B = 8'hAD; #100;
A = 8'h6C; B = 8'hAE; #100;
A = 8'h6C; B = 8'hAF; #100;
A = 8'h6C; B = 8'hB0; #100;
A = 8'h6C; B = 8'hB1; #100;
A = 8'h6C; B = 8'hB2; #100;
A = 8'h6C; B = 8'hB3; #100;
A = 8'h6C; B = 8'hB4; #100;
A = 8'h6C; B = 8'hB5; #100;
A = 8'h6C; B = 8'hB6; #100;
A = 8'h6C; B = 8'hB7; #100;
A = 8'h6C; B = 8'hB8; #100;
A = 8'h6C; B = 8'hB9; #100;
A = 8'h6C; B = 8'hBA; #100;
A = 8'h6C; B = 8'hBB; #100;
A = 8'h6C; B = 8'hBC; #100;
A = 8'h6C; B = 8'hBD; #100;
A = 8'h6C; B = 8'hBE; #100;
A = 8'h6C; B = 8'hBF; #100;
A = 8'h6C; B = 8'hC0; #100;
A = 8'h6C; B = 8'hC1; #100;
A = 8'h6C; B = 8'hC2; #100;
A = 8'h6C; B = 8'hC3; #100;
A = 8'h6C; B = 8'hC4; #100;
A = 8'h6C; B = 8'hC5; #100;
A = 8'h6C; B = 8'hC6; #100;
A = 8'h6C; B = 8'hC7; #100;
A = 8'h6C; B = 8'hC8; #100;
A = 8'h6C; B = 8'hC9; #100;
A = 8'h6C; B = 8'hCA; #100;
A = 8'h6C; B = 8'hCB; #100;
A = 8'h6C; B = 8'hCC; #100;
A = 8'h6C; B = 8'hCD; #100;
A = 8'h6C; B = 8'hCE; #100;
A = 8'h6C; B = 8'hCF; #100;
A = 8'h6C; B = 8'hD0; #100;
A = 8'h6C; B = 8'hD1; #100;
A = 8'h6C; B = 8'hD2; #100;
A = 8'h6C; B = 8'hD3; #100;
A = 8'h6C; B = 8'hD4; #100;
A = 8'h6C; B = 8'hD5; #100;
A = 8'h6C; B = 8'hD6; #100;
A = 8'h6C; B = 8'hD7; #100;
A = 8'h6C; B = 8'hD8; #100;
A = 8'h6C; B = 8'hD9; #100;
A = 8'h6C; B = 8'hDA; #100;
A = 8'h6C; B = 8'hDB; #100;
A = 8'h6C; B = 8'hDC; #100;
A = 8'h6C; B = 8'hDD; #100;
A = 8'h6C; B = 8'hDE; #100;
A = 8'h6C; B = 8'hDF; #100;
A = 8'h6C; B = 8'hE0; #100;
A = 8'h6C; B = 8'hE1; #100;
A = 8'h6C; B = 8'hE2; #100;
A = 8'h6C; B = 8'hE3; #100;
A = 8'h6C; B = 8'hE4; #100;
A = 8'h6C; B = 8'hE5; #100;
A = 8'h6C; B = 8'hE6; #100;
A = 8'h6C; B = 8'hE7; #100;
A = 8'h6C; B = 8'hE8; #100;
A = 8'h6C; B = 8'hE9; #100;
A = 8'h6C; B = 8'hEA; #100;
A = 8'h6C; B = 8'hEB; #100;
A = 8'h6C; B = 8'hEC; #100;
A = 8'h6C; B = 8'hED; #100;
A = 8'h6C; B = 8'hEE; #100;
A = 8'h6C; B = 8'hEF; #100;
A = 8'h6C; B = 8'hF0; #100;
A = 8'h6C; B = 8'hF1; #100;
A = 8'h6C; B = 8'hF2; #100;
A = 8'h6C; B = 8'hF3; #100;
A = 8'h6C; B = 8'hF4; #100;
A = 8'h6C; B = 8'hF5; #100;
A = 8'h6C; B = 8'hF6; #100;
A = 8'h6C; B = 8'hF7; #100;
A = 8'h6C; B = 8'hF8; #100;
A = 8'h6C; B = 8'hF9; #100;
A = 8'h6C; B = 8'hFA; #100;
A = 8'h6C; B = 8'hFB; #100;
A = 8'h6C; B = 8'hFC; #100;
A = 8'h6C; B = 8'hFD; #100;
A = 8'h6C; B = 8'hFE; #100;
A = 8'h6C; B = 8'hFF; #100;
A = 8'h6D; B = 8'h0; #100;
A = 8'h6D; B = 8'h1; #100;
A = 8'h6D; B = 8'h2; #100;
A = 8'h6D; B = 8'h3; #100;
A = 8'h6D; B = 8'h4; #100;
A = 8'h6D; B = 8'h5; #100;
A = 8'h6D; B = 8'h6; #100;
A = 8'h6D; B = 8'h7; #100;
A = 8'h6D; B = 8'h8; #100;
A = 8'h6D; B = 8'h9; #100;
A = 8'h6D; B = 8'hA; #100;
A = 8'h6D; B = 8'hB; #100;
A = 8'h6D; B = 8'hC; #100;
A = 8'h6D; B = 8'hD; #100;
A = 8'h6D; B = 8'hE; #100;
A = 8'h6D; B = 8'hF; #100;
A = 8'h6D; B = 8'h10; #100;
A = 8'h6D; B = 8'h11; #100;
A = 8'h6D; B = 8'h12; #100;
A = 8'h6D; B = 8'h13; #100;
A = 8'h6D; B = 8'h14; #100;
A = 8'h6D; B = 8'h15; #100;
A = 8'h6D; B = 8'h16; #100;
A = 8'h6D; B = 8'h17; #100;
A = 8'h6D; B = 8'h18; #100;
A = 8'h6D; B = 8'h19; #100;
A = 8'h6D; B = 8'h1A; #100;
A = 8'h6D; B = 8'h1B; #100;
A = 8'h6D; B = 8'h1C; #100;
A = 8'h6D; B = 8'h1D; #100;
A = 8'h6D; B = 8'h1E; #100;
A = 8'h6D; B = 8'h1F; #100;
A = 8'h6D; B = 8'h20; #100;
A = 8'h6D; B = 8'h21; #100;
A = 8'h6D; B = 8'h22; #100;
A = 8'h6D; B = 8'h23; #100;
A = 8'h6D; B = 8'h24; #100;
A = 8'h6D; B = 8'h25; #100;
A = 8'h6D; B = 8'h26; #100;
A = 8'h6D; B = 8'h27; #100;
A = 8'h6D; B = 8'h28; #100;
A = 8'h6D; B = 8'h29; #100;
A = 8'h6D; B = 8'h2A; #100;
A = 8'h6D; B = 8'h2B; #100;
A = 8'h6D; B = 8'h2C; #100;
A = 8'h6D; B = 8'h2D; #100;
A = 8'h6D; B = 8'h2E; #100;
A = 8'h6D; B = 8'h2F; #100;
A = 8'h6D; B = 8'h30; #100;
A = 8'h6D; B = 8'h31; #100;
A = 8'h6D; B = 8'h32; #100;
A = 8'h6D; B = 8'h33; #100;
A = 8'h6D; B = 8'h34; #100;
A = 8'h6D; B = 8'h35; #100;
A = 8'h6D; B = 8'h36; #100;
A = 8'h6D; B = 8'h37; #100;
A = 8'h6D; B = 8'h38; #100;
A = 8'h6D; B = 8'h39; #100;
A = 8'h6D; B = 8'h3A; #100;
A = 8'h6D; B = 8'h3B; #100;
A = 8'h6D; B = 8'h3C; #100;
A = 8'h6D; B = 8'h3D; #100;
A = 8'h6D; B = 8'h3E; #100;
A = 8'h6D; B = 8'h3F; #100;
A = 8'h6D; B = 8'h40; #100;
A = 8'h6D; B = 8'h41; #100;
A = 8'h6D; B = 8'h42; #100;
A = 8'h6D; B = 8'h43; #100;
A = 8'h6D; B = 8'h44; #100;
A = 8'h6D; B = 8'h45; #100;
A = 8'h6D; B = 8'h46; #100;
A = 8'h6D; B = 8'h47; #100;
A = 8'h6D; B = 8'h48; #100;
A = 8'h6D; B = 8'h49; #100;
A = 8'h6D; B = 8'h4A; #100;
A = 8'h6D; B = 8'h4B; #100;
A = 8'h6D; B = 8'h4C; #100;
A = 8'h6D; B = 8'h4D; #100;
A = 8'h6D; B = 8'h4E; #100;
A = 8'h6D; B = 8'h4F; #100;
A = 8'h6D; B = 8'h50; #100;
A = 8'h6D; B = 8'h51; #100;
A = 8'h6D; B = 8'h52; #100;
A = 8'h6D; B = 8'h53; #100;
A = 8'h6D; B = 8'h54; #100;
A = 8'h6D; B = 8'h55; #100;
A = 8'h6D; B = 8'h56; #100;
A = 8'h6D; B = 8'h57; #100;
A = 8'h6D; B = 8'h58; #100;
A = 8'h6D; B = 8'h59; #100;
A = 8'h6D; B = 8'h5A; #100;
A = 8'h6D; B = 8'h5B; #100;
A = 8'h6D; B = 8'h5C; #100;
A = 8'h6D; B = 8'h5D; #100;
A = 8'h6D; B = 8'h5E; #100;
A = 8'h6D; B = 8'h5F; #100;
A = 8'h6D; B = 8'h60; #100;
A = 8'h6D; B = 8'h61; #100;
A = 8'h6D; B = 8'h62; #100;
A = 8'h6D; B = 8'h63; #100;
A = 8'h6D; B = 8'h64; #100;
A = 8'h6D; B = 8'h65; #100;
A = 8'h6D; B = 8'h66; #100;
A = 8'h6D; B = 8'h67; #100;
A = 8'h6D; B = 8'h68; #100;
A = 8'h6D; B = 8'h69; #100;
A = 8'h6D; B = 8'h6A; #100;
A = 8'h6D; B = 8'h6B; #100;
A = 8'h6D; B = 8'h6C; #100;
A = 8'h6D; B = 8'h6D; #100;
A = 8'h6D; B = 8'h6E; #100;
A = 8'h6D; B = 8'h6F; #100;
A = 8'h6D; B = 8'h70; #100;
A = 8'h6D; B = 8'h71; #100;
A = 8'h6D; B = 8'h72; #100;
A = 8'h6D; B = 8'h73; #100;
A = 8'h6D; B = 8'h74; #100;
A = 8'h6D; B = 8'h75; #100;
A = 8'h6D; B = 8'h76; #100;
A = 8'h6D; B = 8'h77; #100;
A = 8'h6D; B = 8'h78; #100;
A = 8'h6D; B = 8'h79; #100;
A = 8'h6D; B = 8'h7A; #100;
A = 8'h6D; B = 8'h7B; #100;
A = 8'h6D; B = 8'h7C; #100;
A = 8'h6D; B = 8'h7D; #100;
A = 8'h6D; B = 8'h7E; #100;
A = 8'h6D; B = 8'h7F; #100;
A = 8'h6D; B = 8'h80; #100;
A = 8'h6D; B = 8'h81; #100;
A = 8'h6D; B = 8'h82; #100;
A = 8'h6D; B = 8'h83; #100;
A = 8'h6D; B = 8'h84; #100;
A = 8'h6D; B = 8'h85; #100;
A = 8'h6D; B = 8'h86; #100;
A = 8'h6D; B = 8'h87; #100;
A = 8'h6D; B = 8'h88; #100;
A = 8'h6D; B = 8'h89; #100;
A = 8'h6D; B = 8'h8A; #100;
A = 8'h6D; B = 8'h8B; #100;
A = 8'h6D; B = 8'h8C; #100;
A = 8'h6D; B = 8'h8D; #100;
A = 8'h6D; B = 8'h8E; #100;
A = 8'h6D; B = 8'h8F; #100;
A = 8'h6D; B = 8'h90; #100;
A = 8'h6D; B = 8'h91; #100;
A = 8'h6D; B = 8'h92; #100;
A = 8'h6D; B = 8'h93; #100;
A = 8'h6D; B = 8'h94; #100;
A = 8'h6D; B = 8'h95; #100;
A = 8'h6D; B = 8'h96; #100;
A = 8'h6D; B = 8'h97; #100;
A = 8'h6D; B = 8'h98; #100;
A = 8'h6D; B = 8'h99; #100;
A = 8'h6D; B = 8'h9A; #100;
A = 8'h6D; B = 8'h9B; #100;
A = 8'h6D; B = 8'h9C; #100;
A = 8'h6D; B = 8'h9D; #100;
A = 8'h6D; B = 8'h9E; #100;
A = 8'h6D; B = 8'h9F; #100;
A = 8'h6D; B = 8'hA0; #100;
A = 8'h6D; B = 8'hA1; #100;
A = 8'h6D; B = 8'hA2; #100;
A = 8'h6D; B = 8'hA3; #100;
A = 8'h6D; B = 8'hA4; #100;
A = 8'h6D; B = 8'hA5; #100;
A = 8'h6D; B = 8'hA6; #100;
A = 8'h6D; B = 8'hA7; #100;
A = 8'h6D; B = 8'hA8; #100;
A = 8'h6D; B = 8'hA9; #100;
A = 8'h6D; B = 8'hAA; #100;
A = 8'h6D; B = 8'hAB; #100;
A = 8'h6D; B = 8'hAC; #100;
A = 8'h6D; B = 8'hAD; #100;
A = 8'h6D; B = 8'hAE; #100;
A = 8'h6D; B = 8'hAF; #100;
A = 8'h6D; B = 8'hB0; #100;
A = 8'h6D; B = 8'hB1; #100;
A = 8'h6D; B = 8'hB2; #100;
A = 8'h6D; B = 8'hB3; #100;
A = 8'h6D; B = 8'hB4; #100;
A = 8'h6D; B = 8'hB5; #100;
A = 8'h6D; B = 8'hB6; #100;
A = 8'h6D; B = 8'hB7; #100;
A = 8'h6D; B = 8'hB8; #100;
A = 8'h6D; B = 8'hB9; #100;
A = 8'h6D; B = 8'hBA; #100;
A = 8'h6D; B = 8'hBB; #100;
A = 8'h6D; B = 8'hBC; #100;
A = 8'h6D; B = 8'hBD; #100;
A = 8'h6D; B = 8'hBE; #100;
A = 8'h6D; B = 8'hBF; #100;
A = 8'h6D; B = 8'hC0; #100;
A = 8'h6D; B = 8'hC1; #100;
A = 8'h6D; B = 8'hC2; #100;
A = 8'h6D; B = 8'hC3; #100;
A = 8'h6D; B = 8'hC4; #100;
A = 8'h6D; B = 8'hC5; #100;
A = 8'h6D; B = 8'hC6; #100;
A = 8'h6D; B = 8'hC7; #100;
A = 8'h6D; B = 8'hC8; #100;
A = 8'h6D; B = 8'hC9; #100;
A = 8'h6D; B = 8'hCA; #100;
A = 8'h6D; B = 8'hCB; #100;
A = 8'h6D; B = 8'hCC; #100;
A = 8'h6D; B = 8'hCD; #100;
A = 8'h6D; B = 8'hCE; #100;
A = 8'h6D; B = 8'hCF; #100;
A = 8'h6D; B = 8'hD0; #100;
A = 8'h6D; B = 8'hD1; #100;
A = 8'h6D; B = 8'hD2; #100;
A = 8'h6D; B = 8'hD3; #100;
A = 8'h6D; B = 8'hD4; #100;
A = 8'h6D; B = 8'hD5; #100;
A = 8'h6D; B = 8'hD6; #100;
A = 8'h6D; B = 8'hD7; #100;
A = 8'h6D; B = 8'hD8; #100;
A = 8'h6D; B = 8'hD9; #100;
A = 8'h6D; B = 8'hDA; #100;
A = 8'h6D; B = 8'hDB; #100;
A = 8'h6D; B = 8'hDC; #100;
A = 8'h6D; B = 8'hDD; #100;
A = 8'h6D; B = 8'hDE; #100;
A = 8'h6D; B = 8'hDF; #100;
A = 8'h6D; B = 8'hE0; #100;
A = 8'h6D; B = 8'hE1; #100;
A = 8'h6D; B = 8'hE2; #100;
A = 8'h6D; B = 8'hE3; #100;
A = 8'h6D; B = 8'hE4; #100;
A = 8'h6D; B = 8'hE5; #100;
A = 8'h6D; B = 8'hE6; #100;
A = 8'h6D; B = 8'hE7; #100;
A = 8'h6D; B = 8'hE8; #100;
A = 8'h6D; B = 8'hE9; #100;
A = 8'h6D; B = 8'hEA; #100;
A = 8'h6D; B = 8'hEB; #100;
A = 8'h6D; B = 8'hEC; #100;
A = 8'h6D; B = 8'hED; #100;
A = 8'h6D; B = 8'hEE; #100;
A = 8'h6D; B = 8'hEF; #100;
A = 8'h6D; B = 8'hF0; #100;
A = 8'h6D; B = 8'hF1; #100;
A = 8'h6D; B = 8'hF2; #100;
A = 8'h6D; B = 8'hF3; #100;
A = 8'h6D; B = 8'hF4; #100;
A = 8'h6D; B = 8'hF5; #100;
A = 8'h6D; B = 8'hF6; #100;
A = 8'h6D; B = 8'hF7; #100;
A = 8'h6D; B = 8'hF8; #100;
A = 8'h6D; B = 8'hF9; #100;
A = 8'h6D; B = 8'hFA; #100;
A = 8'h6D; B = 8'hFB; #100;
A = 8'h6D; B = 8'hFC; #100;
A = 8'h6D; B = 8'hFD; #100;
A = 8'h6D; B = 8'hFE; #100;
A = 8'h6D; B = 8'hFF; #100;
A = 8'h6E; B = 8'h0; #100;
A = 8'h6E; B = 8'h1; #100;
A = 8'h6E; B = 8'h2; #100;
A = 8'h6E; B = 8'h3; #100;
A = 8'h6E; B = 8'h4; #100;
A = 8'h6E; B = 8'h5; #100;
A = 8'h6E; B = 8'h6; #100;
A = 8'h6E; B = 8'h7; #100;
A = 8'h6E; B = 8'h8; #100;
A = 8'h6E; B = 8'h9; #100;
A = 8'h6E; B = 8'hA; #100;
A = 8'h6E; B = 8'hB; #100;
A = 8'h6E; B = 8'hC; #100;
A = 8'h6E; B = 8'hD; #100;
A = 8'h6E; B = 8'hE; #100;
A = 8'h6E; B = 8'hF; #100;
A = 8'h6E; B = 8'h10; #100;
A = 8'h6E; B = 8'h11; #100;
A = 8'h6E; B = 8'h12; #100;
A = 8'h6E; B = 8'h13; #100;
A = 8'h6E; B = 8'h14; #100;
A = 8'h6E; B = 8'h15; #100;
A = 8'h6E; B = 8'h16; #100;
A = 8'h6E; B = 8'h17; #100;
A = 8'h6E; B = 8'h18; #100;
A = 8'h6E; B = 8'h19; #100;
A = 8'h6E; B = 8'h1A; #100;
A = 8'h6E; B = 8'h1B; #100;
A = 8'h6E; B = 8'h1C; #100;
A = 8'h6E; B = 8'h1D; #100;
A = 8'h6E; B = 8'h1E; #100;
A = 8'h6E; B = 8'h1F; #100;
A = 8'h6E; B = 8'h20; #100;
A = 8'h6E; B = 8'h21; #100;
A = 8'h6E; B = 8'h22; #100;
A = 8'h6E; B = 8'h23; #100;
A = 8'h6E; B = 8'h24; #100;
A = 8'h6E; B = 8'h25; #100;
A = 8'h6E; B = 8'h26; #100;
A = 8'h6E; B = 8'h27; #100;
A = 8'h6E; B = 8'h28; #100;
A = 8'h6E; B = 8'h29; #100;
A = 8'h6E; B = 8'h2A; #100;
A = 8'h6E; B = 8'h2B; #100;
A = 8'h6E; B = 8'h2C; #100;
A = 8'h6E; B = 8'h2D; #100;
A = 8'h6E; B = 8'h2E; #100;
A = 8'h6E; B = 8'h2F; #100;
A = 8'h6E; B = 8'h30; #100;
A = 8'h6E; B = 8'h31; #100;
A = 8'h6E; B = 8'h32; #100;
A = 8'h6E; B = 8'h33; #100;
A = 8'h6E; B = 8'h34; #100;
A = 8'h6E; B = 8'h35; #100;
A = 8'h6E; B = 8'h36; #100;
A = 8'h6E; B = 8'h37; #100;
A = 8'h6E; B = 8'h38; #100;
A = 8'h6E; B = 8'h39; #100;
A = 8'h6E; B = 8'h3A; #100;
A = 8'h6E; B = 8'h3B; #100;
A = 8'h6E; B = 8'h3C; #100;
A = 8'h6E; B = 8'h3D; #100;
A = 8'h6E; B = 8'h3E; #100;
A = 8'h6E; B = 8'h3F; #100;
A = 8'h6E; B = 8'h40; #100;
A = 8'h6E; B = 8'h41; #100;
A = 8'h6E; B = 8'h42; #100;
A = 8'h6E; B = 8'h43; #100;
A = 8'h6E; B = 8'h44; #100;
A = 8'h6E; B = 8'h45; #100;
A = 8'h6E; B = 8'h46; #100;
A = 8'h6E; B = 8'h47; #100;
A = 8'h6E; B = 8'h48; #100;
A = 8'h6E; B = 8'h49; #100;
A = 8'h6E; B = 8'h4A; #100;
A = 8'h6E; B = 8'h4B; #100;
A = 8'h6E; B = 8'h4C; #100;
A = 8'h6E; B = 8'h4D; #100;
A = 8'h6E; B = 8'h4E; #100;
A = 8'h6E; B = 8'h4F; #100;
A = 8'h6E; B = 8'h50; #100;
A = 8'h6E; B = 8'h51; #100;
A = 8'h6E; B = 8'h52; #100;
A = 8'h6E; B = 8'h53; #100;
A = 8'h6E; B = 8'h54; #100;
A = 8'h6E; B = 8'h55; #100;
A = 8'h6E; B = 8'h56; #100;
A = 8'h6E; B = 8'h57; #100;
A = 8'h6E; B = 8'h58; #100;
A = 8'h6E; B = 8'h59; #100;
A = 8'h6E; B = 8'h5A; #100;
A = 8'h6E; B = 8'h5B; #100;
A = 8'h6E; B = 8'h5C; #100;
A = 8'h6E; B = 8'h5D; #100;
A = 8'h6E; B = 8'h5E; #100;
A = 8'h6E; B = 8'h5F; #100;
A = 8'h6E; B = 8'h60; #100;
A = 8'h6E; B = 8'h61; #100;
A = 8'h6E; B = 8'h62; #100;
A = 8'h6E; B = 8'h63; #100;
A = 8'h6E; B = 8'h64; #100;
A = 8'h6E; B = 8'h65; #100;
A = 8'h6E; B = 8'h66; #100;
A = 8'h6E; B = 8'h67; #100;
A = 8'h6E; B = 8'h68; #100;
A = 8'h6E; B = 8'h69; #100;
A = 8'h6E; B = 8'h6A; #100;
A = 8'h6E; B = 8'h6B; #100;
A = 8'h6E; B = 8'h6C; #100;
A = 8'h6E; B = 8'h6D; #100;
A = 8'h6E; B = 8'h6E; #100;
A = 8'h6E; B = 8'h6F; #100;
A = 8'h6E; B = 8'h70; #100;
A = 8'h6E; B = 8'h71; #100;
A = 8'h6E; B = 8'h72; #100;
A = 8'h6E; B = 8'h73; #100;
A = 8'h6E; B = 8'h74; #100;
A = 8'h6E; B = 8'h75; #100;
A = 8'h6E; B = 8'h76; #100;
A = 8'h6E; B = 8'h77; #100;
A = 8'h6E; B = 8'h78; #100;
A = 8'h6E; B = 8'h79; #100;
A = 8'h6E; B = 8'h7A; #100;
A = 8'h6E; B = 8'h7B; #100;
A = 8'h6E; B = 8'h7C; #100;
A = 8'h6E; B = 8'h7D; #100;
A = 8'h6E; B = 8'h7E; #100;
A = 8'h6E; B = 8'h7F; #100;
A = 8'h6E; B = 8'h80; #100;
A = 8'h6E; B = 8'h81; #100;
A = 8'h6E; B = 8'h82; #100;
A = 8'h6E; B = 8'h83; #100;
A = 8'h6E; B = 8'h84; #100;
A = 8'h6E; B = 8'h85; #100;
A = 8'h6E; B = 8'h86; #100;
A = 8'h6E; B = 8'h87; #100;
A = 8'h6E; B = 8'h88; #100;
A = 8'h6E; B = 8'h89; #100;
A = 8'h6E; B = 8'h8A; #100;
A = 8'h6E; B = 8'h8B; #100;
A = 8'h6E; B = 8'h8C; #100;
A = 8'h6E; B = 8'h8D; #100;
A = 8'h6E; B = 8'h8E; #100;
A = 8'h6E; B = 8'h8F; #100;
A = 8'h6E; B = 8'h90; #100;
A = 8'h6E; B = 8'h91; #100;
A = 8'h6E; B = 8'h92; #100;
A = 8'h6E; B = 8'h93; #100;
A = 8'h6E; B = 8'h94; #100;
A = 8'h6E; B = 8'h95; #100;
A = 8'h6E; B = 8'h96; #100;
A = 8'h6E; B = 8'h97; #100;
A = 8'h6E; B = 8'h98; #100;
A = 8'h6E; B = 8'h99; #100;
A = 8'h6E; B = 8'h9A; #100;
A = 8'h6E; B = 8'h9B; #100;
A = 8'h6E; B = 8'h9C; #100;
A = 8'h6E; B = 8'h9D; #100;
A = 8'h6E; B = 8'h9E; #100;
A = 8'h6E; B = 8'h9F; #100;
A = 8'h6E; B = 8'hA0; #100;
A = 8'h6E; B = 8'hA1; #100;
A = 8'h6E; B = 8'hA2; #100;
A = 8'h6E; B = 8'hA3; #100;
A = 8'h6E; B = 8'hA4; #100;
A = 8'h6E; B = 8'hA5; #100;
A = 8'h6E; B = 8'hA6; #100;
A = 8'h6E; B = 8'hA7; #100;
A = 8'h6E; B = 8'hA8; #100;
A = 8'h6E; B = 8'hA9; #100;
A = 8'h6E; B = 8'hAA; #100;
A = 8'h6E; B = 8'hAB; #100;
A = 8'h6E; B = 8'hAC; #100;
A = 8'h6E; B = 8'hAD; #100;
A = 8'h6E; B = 8'hAE; #100;
A = 8'h6E; B = 8'hAF; #100;
A = 8'h6E; B = 8'hB0; #100;
A = 8'h6E; B = 8'hB1; #100;
A = 8'h6E; B = 8'hB2; #100;
A = 8'h6E; B = 8'hB3; #100;
A = 8'h6E; B = 8'hB4; #100;
A = 8'h6E; B = 8'hB5; #100;
A = 8'h6E; B = 8'hB6; #100;
A = 8'h6E; B = 8'hB7; #100;
A = 8'h6E; B = 8'hB8; #100;
A = 8'h6E; B = 8'hB9; #100;
A = 8'h6E; B = 8'hBA; #100;
A = 8'h6E; B = 8'hBB; #100;
A = 8'h6E; B = 8'hBC; #100;
A = 8'h6E; B = 8'hBD; #100;
A = 8'h6E; B = 8'hBE; #100;
A = 8'h6E; B = 8'hBF; #100;
A = 8'h6E; B = 8'hC0; #100;
A = 8'h6E; B = 8'hC1; #100;
A = 8'h6E; B = 8'hC2; #100;
A = 8'h6E; B = 8'hC3; #100;
A = 8'h6E; B = 8'hC4; #100;
A = 8'h6E; B = 8'hC5; #100;
A = 8'h6E; B = 8'hC6; #100;
A = 8'h6E; B = 8'hC7; #100;
A = 8'h6E; B = 8'hC8; #100;
A = 8'h6E; B = 8'hC9; #100;
A = 8'h6E; B = 8'hCA; #100;
A = 8'h6E; B = 8'hCB; #100;
A = 8'h6E; B = 8'hCC; #100;
A = 8'h6E; B = 8'hCD; #100;
A = 8'h6E; B = 8'hCE; #100;
A = 8'h6E; B = 8'hCF; #100;
A = 8'h6E; B = 8'hD0; #100;
A = 8'h6E; B = 8'hD1; #100;
A = 8'h6E; B = 8'hD2; #100;
A = 8'h6E; B = 8'hD3; #100;
A = 8'h6E; B = 8'hD4; #100;
A = 8'h6E; B = 8'hD5; #100;
A = 8'h6E; B = 8'hD6; #100;
A = 8'h6E; B = 8'hD7; #100;
A = 8'h6E; B = 8'hD8; #100;
A = 8'h6E; B = 8'hD9; #100;
A = 8'h6E; B = 8'hDA; #100;
A = 8'h6E; B = 8'hDB; #100;
A = 8'h6E; B = 8'hDC; #100;
A = 8'h6E; B = 8'hDD; #100;
A = 8'h6E; B = 8'hDE; #100;
A = 8'h6E; B = 8'hDF; #100;
A = 8'h6E; B = 8'hE0; #100;
A = 8'h6E; B = 8'hE1; #100;
A = 8'h6E; B = 8'hE2; #100;
A = 8'h6E; B = 8'hE3; #100;
A = 8'h6E; B = 8'hE4; #100;
A = 8'h6E; B = 8'hE5; #100;
A = 8'h6E; B = 8'hE6; #100;
A = 8'h6E; B = 8'hE7; #100;
A = 8'h6E; B = 8'hE8; #100;
A = 8'h6E; B = 8'hE9; #100;
A = 8'h6E; B = 8'hEA; #100;
A = 8'h6E; B = 8'hEB; #100;
A = 8'h6E; B = 8'hEC; #100;
A = 8'h6E; B = 8'hED; #100;
A = 8'h6E; B = 8'hEE; #100;
A = 8'h6E; B = 8'hEF; #100;
A = 8'h6E; B = 8'hF0; #100;
A = 8'h6E; B = 8'hF1; #100;
A = 8'h6E; B = 8'hF2; #100;
A = 8'h6E; B = 8'hF3; #100;
A = 8'h6E; B = 8'hF4; #100;
A = 8'h6E; B = 8'hF5; #100;
A = 8'h6E; B = 8'hF6; #100;
A = 8'h6E; B = 8'hF7; #100;
A = 8'h6E; B = 8'hF8; #100;
A = 8'h6E; B = 8'hF9; #100;
A = 8'h6E; B = 8'hFA; #100;
A = 8'h6E; B = 8'hFB; #100;
A = 8'h6E; B = 8'hFC; #100;
A = 8'h6E; B = 8'hFD; #100;
A = 8'h6E; B = 8'hFE; #100;
A = 8'h6E; B = 8'hFF; #100;
A = 8'h6F; B = 8'h0; #100;
A = 8'h6F; B = 8'h1; #100;
A = 8'h6F; B = 8'h2; #100;
A = 8'h6F; B = 8'h3; #100;
A = 8'h6F; B = 8'h4; #100;
A = 8'h6F; B = 8'h5; #100;
A = 8'h6F; B = 8'h6; #100;
A = 8'h6F; B = 8'h7; #100;
A = 8'h6F; B = 8'h8; #100;
A = 8'h6F; B = 8'h9; #100;
A = 8'h6F; B = 8'hA; #100;
A = 8'h6F; B = 8'hB; #100;
A = 8'h6F; B = 8'hC; #100;
A = 8'h6F; B = 8'hD; #100;
A = 8'h6F; B = 8'hE; #100;
A = 8'h6F; B = 8'hF; #100;
A = 8'h6F; B = 8'h10; #100;
A = 8'h6F; B = 8'h11; #100;
A = 8'h6F; B = 8'h12; #100;
A = 8'h6F; B = 8'h13; #100;
A = 8'h6F; B = 8'h14; #100;
A = 8'h6F; B = 8'h15; #100;
A = 8'h6F; B = 8'h16; #100;
A = 8'h6F; B = 8'h17; #100;
A = 8'h6F; B = 8'h18; #100;
A = 8'h6F; B = 8'h19; #100;
A = 8'h6F; B = 8'h1A; #100;
A = 8'h6F; B = 8'h1B; #100;
A = 8'h6F; B = 8'h1C; #100;
A = 8'h6F; B = 8'h1D; #100;
A = 8'h6F; B = 8'h1E; #100;
A = 8'h6F; B = 8'h1F; #100;
A = 8'h6F; B = 8'h20; #100;
A = 8'h6F; B = 8'h21; #100;
A = 8'h6F; B = 8'h22; #100;
A = 8'h6F; B = 8'h23; #100;
A = 8'h6F; B = 8'h24; #100;
A = 8'h6F; B = 8'h25; #100;
A = 8'h6F; B = 8'h26; #100;
A = 8'h6F; B = 8'h27; #100;
A = 8'h6F; B = 8'h28; #100;
A = 8'h6F; B = 8'h29; #100;
A = 8'h6F; B = 8'h2A; #100;
A = 8'h6F; B = 8'h2B; #100;
A = 8'h6F; B = 8'h2C; #100;
A = 8'h6F; B = 8'h2D; #100;
A = 8'h6F; B = 8'h2E; #100;
A = 8'h6F; B = 8'h2F; #100;
A = 8'h6F; B = 8'h30; #100;
A = 8'h6F; B = 8'h31; #100;
A = 8'h6F; B = 8'h32; #100;
A = 8'h6F; B = 8'h33; #100;
A = 8'h6F; B = 8'h34; #100;
A = 8'h6F; B = 8'h35; #100;
A = 8'h6F; B = 8'h36; #100;
A = 8'h6F; B = 8'h37; #100;
A = 8'h6F; B = 8'h38; #100;
A = 8'h6F; B = 8'h39; #100;
A = 8'h6F; B = 8'h3A; #100;
A = 8'h6F; B = 8'h3B; #100;
A = 8'h6F; B = 8'h3C; #100;
A = 8'h6F; B = 8'h3D; #100;
A = 8'h6F; B = 8'h3E; #100;
A = 8'h6F; B = 8'h3F; #100;
A = 8'h6F; B = 8'h40; #100;
A = 8'h6F; B = 8'h41; #100;
A = 8'h6F; B = 8'h42; #100;
A = 8'h6F; B = 8'h43; #100;
A = 8'h6F; B = 8'h44; #100;
A = 8'h6F; B = 8'h45; #100;
A = 8'h6F; B = 8'h46; #100;
A = 8'h6F; B = 8'h47; #100;
A = 8'h6F; B = 8'h48; #100;
A = 8'h6F; B = 8'h49; #100;
A = 8'h6F; B = 8'h4A; #100;
A = 8'h6F; B = 8'h4B; #100;
A = 8'h6F; B = 8'h4C; #100;
A = 8'h6F; B = 8'h4D; #100;
A = 8'h6F; B = 8'h4E; #100;
A = 8'h6F; B = 8'h4F; #100;
A = 8'h6F; B = 8'h50; #100;
A = 8'h6F; B = 8'h51; #100;
A = 8'h6F; B = 8'h52; #100;
A = 8'h6F; B = 8'h53; #100;
A = 8'h6F; B = 8'h54; #100;
A = 8'h6F; B = 8'h55; #100;
A = 8'h6F; B = 8'h56; #100;
A = 8'h6F; B = 8'h57; #100;
A = 8'h6F; B = 8'h58; #100;
A = 8'h6F; B = 8'h59; #100;
A = 8'h6F; B = 8'h5A; #100;
A = 8'h6F; B = 8'h5B; #100;
A = 8'h6F; B = 8'h5C; #100;
A = 8'h6F; B = 8'h5D; #100;
A = 8'h6F; B = 8'h5E; #100;
A = 8'h6F; B = 8'h5F; #100;
A = 8'h6F; B = 8'h60; #100;
A = 8'h6F; B = 8'h61; #100;
A = 8'h6F; B = 8'h62; #100;
A = 8'h6F; B = 8'h63; #100;
A = 8'h6F; B = 8'h64; #100;
A = 8'h6F; B = 8'h65; #100;
A = 8'h6F; B = 8'h66; #100;
A = 8'h6F; B = 8'h67; #100;
A = 8'h6F; B = 8'h68; #100;
A = 8'h6F; B = 8'h69; #100;
A = 8'h6F; B = 8'h6A; #100;
A = 8'h6F; B = 8'h6B; #100;
A = 8'h6F; B = 8'h6C; #100;
A = 8'h6F; B = 8'h6D; #100;
A = 8'h6F; B = 8'h6E; #100;
A = 8'h6F; B = 8'h6F; #100;
A = 8'h6F; B = 8'h70; #100;
A = 8'h6F; B = 8'h71; #100;
A = 8'h6F; B = 8'h72; #100;
A = 8'h6F; B = 8'h73; #100;
A = 8'h6F; B = 8'h74; #100;
A = 8'h6F; B = 8'h75; #100;
A = 8'h6F; B = 8'h76; #100;
A = 8'h6F; B = 8'h77; #100;
A = 8'h6F; B = 8'h78; #100;
A = 8'h6F; B = 8'h79; #100;
A = 8'h6F; B = 8'h7A; #100;
A = 8'h6F; B = 8'h7B; #100;
A = 8'h6F; B = 8'h7C; #100;
A = 8'h6F; B = 8'h7D; #100;
A = 8'h6F; B = 8'h7E; #100;
A = 8'h6F; B = 8'h7F; #100;
A = 8'h6F; B = 8'h80; #100;
A = 8'h6F; B = 8'h81; #100;
A = 8'h6F; B = 8'h82; #100;
A = 8'h6F; B = 8'h83; #100;
A = 8'h6F; B = 8'h84; #100;
A = 8'h6F; B = 8'h85; #100;
A = 8'h6F; B = 8'h86; #100;
A = 8'h6F; B = 8'h87; #100;
A = 8'h6F; B = 8'h88; #100;
A = 8'h6F; B = 8'h89; #100;
A = 8'h6F; B = 8'h8A; #100;
A = 8'h6F; B = 8'h8B; #100;
A = 8'h6F; B = 8'h8C; #100;
A = 8'h6F; B = 8'h8D; #100;
A = 8'h6F; B = 8'h8E; #100;
A = 8'h6F; B = 8'h8F; #100;
A = 8'h6F; B = 8'h90; #100;
A = 8'h6F; B = 8'h91; #100;
A = 8'h6F; B = 8'h92; #100;
A = 8'h6F; B = 8'h93; #100;
A = 8'h6F; B = 8'h94; #100;
A = 8'h6F; B = 8'h95; #100;
A = 8'h6F; B = 8'h96; #100;
A = 8'h6F; B = 8'h97; #100;
A = 8'h6F; B = 8'h98; #100;
A = 8'h6F; B = 8'h99; #100;
A = 8'h6F; B = 8'h9A; #100;
A = 8'h6F; B = 8'h9B; #100;
A = 8'h6F; B = 8'h9C; #100;
A = 8'h6F; B = 8'h9D; #100;
A = 8'h6F; B = 8'h9E; #100;
A = 8'h6F; B = 8'h9F; #100;
A = 8'h6F; B = 8'hA0; #100;
A = 8'h6F; B = 8'hA1; #100;
A = 8'h6F; B = 8'hA2; #100;
A = 8'h6F; B = 8'hA3; #100;
A = 8'h6F; B = 8'hA4; #100;
A = 8'h6F; B = 8'hA5; #100;
A = 8'h6F; B = 8'hA6; #100;
A = 8'h6F; B = 8'hA7; #100;
A = 8'h6F; B = 8'hA8; #100;
A = 8'h6F; B = 8'hA9; #100;
A = 8'h6F; B = 8'hAA; #100;
A = 8'h6F; B = 8'hAB; #100;
A = 8'h6F; B = 8'hAC; #100;
A = 8'h6F; B = 8'hAD; #100;
A = 8'h6F; B = 8'hAE; #100;
A = 8'h6F; B = 8'hAF; #100;
A = 8'h6F; B = 8'hB0; #100;
A = 8'h6F; B = 8'hB1; #100;
A = 8'h6F; B = 8'hB2; #100;
A = 8'h6F; B = 8'hB3; #100;
A = 8'h6F; B = 8'hB4; #100;
A = 8'h6F; B = 8'hB5; #100;
A = 8'h6F; B = 8'hB6; #100;
A = 8'h6F; B = 8'hB7; #100;
A = 8'h6F; B = 8'hB8; #100;
A = 8'h6F; B = 8'hB9; #100;
A = 8'h6F; B = 8'hBA; #100;
A = 8'h6F; B = 8'hBB; #100;
A = 8'h6F; B = 8'hBC; #100;
A = 8'h6F; B = 8'hBD; #100;
A = 8'h6F; B = 8'hBE; #100;
A = 8'h6F; B = 8'hBF; #100;
A = 8'h6F; B = 8'hC0; #100;
A = 8'h6F; B = 8'hC1; #100;
A = 8'h6F; B = 8'hC2; #100;
A = 8'h6F; B = 8'hC3; #100;
A = 8'h6F; B = 8'hC4; #100;
A = 8'h6F; B = 8'hC5; #100;
A = 8'h6F; B = 8'hC6; #100;
A = 8'h6F; B = 8'hC7; #100;
A = 8'h6F; B = 8'hC8; #100;
A = 8'h6F; B = 8'hC9; #100;
A = 8'h6F; B = 8'hCA; #100;
A = 8'h6F; B = 8'hCB; #100;
A = 8'h6F; B = 8'hCC; #100;
A = 8'h6F; B = 8'hCD; #100;
A = 8'h6F; B = 8'hCE; #100;
A = 8'h6F; B = 8'hCF; #100;
A = 8'h6F; B = 8'hD0; #100;
A = 8'h6F; B = 8'hD1; #100;
A = 8'h6F; B = 8'hD2; #100;
A = 8'h6F; B = 8'hD3; #100;
A = 8'h6F; B = 8'hD4; #100;
A = 8'h6F; B = 8'hD5; #100;
A = 8'h6F; B = 8'hD6; #100;
A = 8'h6F; B = 8'hD7; #100;
A = 8'h6F; B = 8'hD8; #100;
A = 8'h6F; B = 8'hD9; #100;
A = 8'h6F; B = 8'hDA; #100;
A = 8'h6F; B = 8'hDB; #100;
A = 8'h6F; B = 8'hDC; #100;
A = 8'h6F; B = 8'hDD; #100;
A = 8'h6F; B = 8'hDE; #100;
A = 8'h6F; B = 8'hDF; #100;
A = 8'h6F; B = 8'hE0; #100;
A = 8'h6F; B = 8'hE1; #100;
A = 8'h6F; B = 8'hE2; #100;
A = 8'h6F; B = 8'hE3; #100;
A = 8'h6F; B = 8'hE4; #100;
A = 8'h6F; B = 8'hE5; #100;
A = 8'h6F; B = 8'hE6; #100;
A = 8'h6F; B = 8'hE7; #100;
A = 8'h6F; B = 8'hE8; #100;
A = 8'h6F; B = 8'hE9; #100;
A = 8'h6F; B = 8'hEA; #100;
A = 8'h6F; B = 8'hEB; #100;
A = 8'h6F; B = 8'hEC; #100;
A = 8'h6F; B = 8'hED; #100;
A = 8'h6F; B = 8'hEE; #100;
A = 8'h6F; B = 8'hEF; #100;
A = 8'h6F; B = 8'hF0; #100;
A = 8'h6F; B = 8'hF1; #100;
A = 8'h6F; B = 8'hF2; #100;
A = 8'h6F; B = 8'hF3; #100;
A = 8'h6F; B = 8'hF4; #100;
A = 8'h6F; B = 8'hF5; #100;
A = 8'h6F; B = 8'hF6; #100;
A = 8'h6F; B = 8'hF7; #100;
A = 8'h6F; B = 8'hF8; #100;
A = 8'h6F; B = 8'hF9; #100;
A = 8'h6F; B = 8'hFA; #100;
A = 8'h6F; B = 8'hFB; #100;
A = 8'h6F; B = 8'hFC; #100;
A = 8'h6F; B = 8'hFD; #100;
A = 8'h6F; B = 8'hFE; #100;
A = 8'h6F; B = 8'hFF; #100;
A = 8'h70; B = 8'h0; #100;
A = 8'h70; B = 8'h1; #100;
A = 8'h70; B = 8'h2; #100;
A = 8'h70; B = 8'h3; #100;
A = 8'h70; B = 8'h4; #100;
A = 8'h70; B = 8'h5; #100;
A = 8'h70; B = 8'h6; #100;
A = 8'h70; B = 8'h7; #100;
A = 8'h70; B = 8'h8; #100;
A = 8'h70; B = 8'h9; #100;
A = 8'h70; B = 8'hA; #100;
A = 8'h70; B = 8'hB; #100;
A = 8'h70; B = 8'hC; #100;
A = 8'h70; B = 8'hD; #100;
A = 8'h70; B = 8'hE; #100;
A = 8'h70; B = 8'hF; #100;
A = 8'h70; B = 8'h10; #100;
A = 8'h70; B = 8'h11; #100;
A = 8'h70; B = 8'h12; #100;
A = 8'h70; B = 8'h13; #100;
A = 8'h70; B = 8'h14; #100;
A = 8'h70; B = 8'h15; #100;
A = 8'h70; B = 8'h16; #100;
A = 8'h70; B = 8'h17; #100;
A = 8'h70; B = 8'h18; #100;
A = 8'h70; B = 8'h19; #100;
A = 8'h70; B = 8'h1A; #100;
A = 8'h70; B = 8'h1B; #100;
A = 8'h70; B = 8'h1C; #100;
A = 8'h70; B = 8'h1D; #100;
A = 8'h70; B = 8'h1E; #100;
A = 8'h70; B = 8'h1F; #100;
A = 8'h70; B = 8'h20; #100;
A = 8'h70; B = 8'h21; #100;
A = 8'h70; B = 8'h22; #100;
A = 8'h70; B = 8'h23; #100;
A = 8'h70; B = 8'h24; #100;
A = 8'h70; B = 8'h25; #100;
A = 8'h70; B = 8'h26; #100;
A = 8'h70; B = 8'h27; #100;
A = 8'h70; B = 8'h28; #100;
A = 8'h70; B = 8'h29; #100;
A = 8'h70; B = 8'h2A; #100;
A = 8'h70; B = 8'h2B; #100;
A = 8'h70; B = 8'h2C; #100;
A = 8'h70; B = 8'h2D; #100;
A = 8'h70; B = 8'h2E; #100;
A = 8'h70; B = 8'h2F; #100;
A = 8'h70; B = 8'h30; #100;
A = 8'h70; B = 8'h31; #100;
A = 8'h70; B = 8'h32; #100;
A = 8'h70; B = 8'h33; #100;
A = 8'h70; B = 8'h34; #100;
A = 8'h70; B = 8'h35; #100;
A = 8'h70; B = 8'h36; #100;
A = 8'h70; B = 8'h37; #100;
A = 8'h70; B = 8'h38; #100;
A = 8'h70; B = 8'h39; #100;
A = 8'h70; B = 8'h3A; #100;
A = 8'h70; B = 8'h3B; #100;
A = 8'h70; B = 8'h3C; #100;
A = 8'h70; B = 8'h3D; #100;
A = 8'h70; B = 8'h3E; #100;
A = 8'h70; B = 8'h3F; #100;
A = 8'h70; B = 8'h40; #100;
A = 8'h70; B = 8'h41; #100;
A = 8'h70; B = 8'h42; #100;
A = 8'h70; B = 8'h43; #100;
A = 8'h70; B = 8'h44; #100;
A = 8'h70; B = 8'h45; #100;
A = 8'h70; B = 8'h46; #100;
A = 8'h70; B = 8'h47; #100;
A = 8'h70; B = 8'h48; #100;
A = 8'h70; B = 8'h49; #100;
A = 8'h70; B = 8'h4A; #100;
A = 8'h70; B = 8'h4B; #100;
A = 8'h70; B = 8'h4C; #100;
A = 8'h70; B = 8'h4D; #100;
A = 8'h70; B = 8'h4E; #100;
A = 8'h70; B = 8'h4F; #100;
A = 8'h70; B = 8'h50; #100;
A = 8'h70; B = 8'h51; #100;
A = 8'h70; B = 8'h52; #100;
A = 8'h70; B = 8'h53; #100;
A = 8'h70; B = 8'h54; #100;
A = 8'h70; B = 8'h55; #100;
A = 8'h70; B = 8'h56; #100;
A = 8'h70; B = 8'h57; #100;
A = 8'h70; B = 8'h58; #100;
A = 8'h70; B = 8'h59; #100;
A = 8'h70; B = 8'h5A; #100;
A = 8'h70; B = 8'h5B; #100;
A = 8'h70; B = 8'h5C; #100;
A = 8'h70; B = 8'h5D; #100;
A = 8'h70; B = 8'h5E; #100;
A = 8'h70; B = 8'h5F; #100;
A = 8'h70; B = 8'h60; #100;
A = 8'h70; B = 8'h61; #100;
A = 8'h70; B = 8'h62; #100;
A = 8'h70; B = 8'h63; #100;
A = 8'h70; B = 8'h64; #100;
A = 8'h70; B = 8'h65; #100;
A = 8'h70; B = 8'h66; #100;
A = 8'h70; B = 8'h67; #100;
A = 8'h70; B = 8'h68; #100;
A = 8'h70; B = 8'h69; #100;
A = 8'h70; B = 8'h6A; #100;
A = 8'h70; B = 8'h6B; #100;
A = 8'h70; B = 8'h6C; #100;
A = 8'h70; B = 8'h6D; #100;
A = 8'h70; B = 8'h6E; #100;
A = 8'h70; B = 8'h6F; #100;
A = 8'h70; B = 8'h70; #100;
A = 8'h70; B = 8'h71; #100;
A = 8'h70; B = 8'h72; #100;
A = 8'h70; B = 8'h73; #100;
A = 8'h70; B = 8'h74; #100;
A = 8'h70; B = 8'h75; #100;
A = 8'h70; B = 8'h76; #100;
A = 8'h70; B = 8'h77; #100;
A = 8'h70; B = 8'h78; #100;
A = 8'h70; B = 8'h79; #100;
A = 8'h70; B = 8'h7A; #100;
A = 8'h70; B = 8'h7B; #100;
A = 8'h70; B = 8'h7C; #100;
A = 8'h70; B = 8'h7D; #100;
A = 8'h70; B = 8'h7E; #100;
A = 8'h70; B = 8'h7F; #100;
A = 8'h70; B = 8'h80; #100;
A = 8'h70; B = 8'h81; #100;
A = 8'h70; B = 8'h82; #100;
A = 8'h70; B = 8'h83; #100;
A = 8'h70; B = 8'h84; #100;
A = 8'h70; B = 8'h85; #100;
A = 8'h70; B = 8'h86; #100;
A = 8'h70; B = 8'h87; #100;
A = 8'h70; B = 8'h88; #100;
A = 8'h70; B = 8'h89; #100;
A = 8'h70; B = 8'h8A; #100;
A = 8'h70; B = 8'h8B; #100;
A = 8'h70; B = 8'h8C; #100;
A = 8'h70; B = 8'h8D; #100;
A = 8'h70; B = 8'h8E; #100;
A = 8'h70; B = 8'h8F; #100;
A = 8'h70; B = 8'h90; #100;
A = 8'h70; B = 8'h91; #100;
A = 8'h70; B = 8'h92; #100;
A = 8'h70; B = 8'h93; #100;
A = 8'h70; B = 8'h94; #100;
A = 8'h70; B = 8'h95; #100;
A = 8'h70; B = 8'h96; #100;
A = 8'h70; B = 8'h97; #100;
A = 8'h70; B = 8'h98; #100;
A = 8'h70; B = 8'h99; #100;
A = 8'h70; B = 8'h9A; #100;
A = 8'h70; B = 8'h9B; #100;
A = 8'h70; B = 8'h9C; #100;
A = 8'h70; B = 8'h9D; #100;
A = 8'h70; B = 8'h9E; #100;
A = 8'h70; B = 8'h9F; #100;
A = 8'h70; B = 8'hA0; #100;
A = 8'h70; B = 8'hA1; #100;
A = 8'h70; B = 8'hA2; #100;
A = 8'h70; B = 8'hA3; #100;
A = 8'h70; B = 8'hA4; #100;
A = 8'h70; B = 8'hA5; #100;
A = 8'h70; B = 8'hA6; #100;
A = 8'h70; B = 8'hA7; #100;
A = 8'h70; B = 8'hA8; #100;
A = 8'h70; B = 8'hA9; #100;
A = 8'h70; B = 8'hAA; #100;
A = 8'h70; B = 8'hAB; #100;
A = 8'h70; B = 8'hAC; #100;
A = 8'h70; B = 8'hAD; #100;
A = 8'h70; B = 8'hAE; #100;
A = 8'h70; B = 8'hAF; #100;
A = 8'h70; B = 8'hB0; #100;
A = 8'h70; B = 8'hB1; #100;
A = 8'h70; B = 8'hB2; #100;
A = 8'h70; B = 8'hB3; #100;
A = 8'h70; B = 8'hB4; #100;
A = 8'h70; B = 8'hB5; #100;
A = 8'h70; B = 8'hB6; #100;
A = 8'h70; B = 8'hB7; #100;
A = 8'h70; B = 8'hB8; #100;
A = 8'h70; B = 8'hB9; #100;
A = 8'h70; B = 8'hBA; #100;
A = 8'h70; B = 8'hBB; #100;
A = 8'h70; B = 8'hBC; #100;
A = 8'h70; B = 8'hBD; #100;
A = 8'h70; B = 8'hBE; #100;
A = 8'h70; B = 8'hBF; #100;
A = 8'h70; B = 8'hC0; #100;
A = 8'h70; B = 8'hC1; #100;
A = 8'h70; B = 8'hC2; #100;
A = 8'h70; B = 8'hC3; #100;
A = 8'h70; B = 8'hC4; #100;
A = 8'h70; B = 8'hC5; #100;
A = 8'h70; B = 8'hC6; #100;
A = 8'h70; B = 8'hC7; #100;
A = 8'h70; B = 8'hC8; #100;
A = 8'h70; B = 8'hC9; #100;
A = 8'h70; B = 8'hCA; #100;
A = 8'h70; B = 8'hCB; #100;
A = 8'h70; B = 8'hCC; #100;
A = 8'h70; B = 8'hCD; #100;
A = 8'h70; B = 8'hCE; #100;
A = 8'h70; B = 8'hCF; #100;
A = 8'h70; B = 8'hD0; #100;
A = 8'h70; B = 8'hD1; #100;
A = 8'h70; B = 8'hD2; #100;
A = 8'h70; B = 8'hD3; #100;
A = 8'h70; B = 8'hD4; #100;
A = 8'h70; B = 8'hD5; #100;
A = 8'h70; B = 8'hD6; #100;
A = 8'h70; B = 8'hD7; #100;
A = 8'h70; B = 8'hD8; #100;
A = 8'h70; B = 8'hD9; #100;
A = 8'h70; B = 8'hDA; #100;
A = 8'h70; B = 8'hDB; #100;
A = 8'h70; B = 8'hDC; #100;
A = 8'h70; B = 8'hDD; #100;
A = 8'h70; B = 8'hDE; #100;
A = 8'h70; B = 8'hDF; #100;
A = 8'h70; B = 8'hE0; #100;
A = 8'h70; B = 8'hE1; #100;
A = 8'h70; B = 8'hE2; #100;
A = 8'h70; B = 8'hE3; #100;
A = 8'h70; B = 8'hE4; #100;
A = 8'h70; B = 8'hE5; #100;
A = 8'h70; B = 8'hE6; #100;
A = 8'h70; B = 8'hE7; #100;
A = 8'h70; B = 8'hE8; #100;
A = 8'h70; B = 8'hE9; #100;
A = 8'h70; B = 8'hEA; #100;
A = 8'h70; B = 8'hEB; #100;
A = 8'h70; B = 8'hEC; #100;
A = 8'h70; B = 8'hED; #100;
A = 8'h70; B = 8'hEE; #100;
A = 8'h70; B = 8'hEF; #100;
A = 8'h70; B = 8'hF0; #100;
A = 8'h70; B = 8'hF1; #100;
A = 8'h70; B = 8'hF2; #100;
A = 8'h70; B = 8'hF3; #100;
A = 8'h70; B = 8'hF4; #100;
A = 8'h70; B = 8'hF5; #100;
A = 8'h70; B = 8'hF6; #100;
A = 8'h70; B = 8'hF7; #100;
A = 8'h70; B = 8'hF8; #100;
A = 8'h70; B = 8'hF9; #100;
A = 8'h70; B = 8'hFA; #100;
A = 8'h70; B = 8'hFB; #100;
A = 8'h70; B = 8'hFC; #100;
A = 8'h70; B = 8'hFD; #100;
A = 8'h70; B = 8'hFE; #100;
A = 8'h70; B = 8'hFF; #100;
A = 8'h71; B = 8'h0; #100;
A = 8'h71; B = 8'h1; #100;
A = 8'h71; B = 8'h2; #100;
A = 8'h71; B = 8'h3; #100;
A = 8'h71; B = 8'h4; #100;
A = 8'h71; B = 8'h5; #100;
A = 8'h71; B = 8'h6; #100;
A = 8'h71; B = 8'h7; #100;
A = 8'h71; B = 8'h8; #100;
A = 8'h71; B = 8'h9; #100;
A = 8'h71; B = 8'hA; #100;
A = 8'h71; B = 8'hB; #100;
A = 8'h71; B = 8'hC; #100;
A = 8'h71; B = 8'hD; #100;
A = 8'h71; B = 8'hE; #100;
A = 8'h71; B = 8'hF; #100;
A = 8'h71; B = 8'h10; #100;
A = 8'h71; B = 8'h11; #100;
A = 8'h71; B = 8'h12; #100;
A = 8'h71; B = 8'h13; #100;
A = 8'h71; B = 8'h14; #100;
A = 8'h71; B = 8'h15; #100;
A = 8'h71; B = 8'h16; #100;
A = 8'h71; B = 8'h17; #100;
A = 8'h71; B = 8'h18; #100;
A = 8'h71; B = 8'h19; #100;
A = 8'h71; B = 8'h1A; #100;
A = 8'h71; B = 8'h1B; #100;
A = 8'h71; B = 8'h1C; #100;
A = 8'h71; B = 8'h1D; #100;
A = 8'h71; B = 8'h1E; #100;
A = 8'h71; B = 8'h1F; #100;
A = 8'h71; B = 8'h20; #100;
A = 8'h71; B = 8'h21; #100;
A = 8'h71; B = 8'h22; #100;
A = 8'h71; B = 8'h23; #100;
A = 8'h71; B = 8'h24; #100;
A = 8'h71; B = 8'h25; #100;
A = 8'h71; B = 8'h26; #100;
A = 8'h71; B = 8'h27; #100;
A = 8'h71; B = 8'h28; #100;
A = 8'h71; B = 8'h29; #100;
A = 8'h71; B = 8'h2A; #100;
A = 8'h71; B = 8'h2B; #100;
A = 8'h71; B = 8'h2C; #100;
A = 8'h71; B = 8'h2D; #100;
A = 8'h71; B = 8'h2E; #100;
A = 8'h71; B = 8'h2F; #100;
A = 8'h71; B = 8'h30; #100;
A = 8'h71; B = 8'h31; #100;
A = 8'h71; B = 8'h32; #100;
A = 8'h71; B = 8'h33; #100;
A = 8'h71; B = 8'h34; #100;
A = 8'h71; B = 8'h35; #100;
A = 8'h71; B = 8'h36; #100;
A = 8'h71; B = 8'h37; #100;
A = 8'h71; B = 8'h38; #100;
A = 8'h71; B = 8'h39; #100;
A = 8'h71; B = 8'h3A; #100;
A = 8'h71; B = 8'h3B; #100;
A = 8'h71; B = 8'h3C; #100;
A = 8'h71; B = 8'h3D; #100;
A = 8'h71; B = 8'h3E; #100;
A = 8'h71; B = 8'h3F; #100;
A = 8'h71; B = 8'h40; #100;
A = 8'h71; B = 8'h41; #100;
A = 8'h71; B = 8'h42; #100;
A = 8'h71; B = 8'h43; #100;
A = 8'h71; B = 8'h44; #100;
A = 8'h71; B = 8'h45; #100;
A = 8'h71; B = 8'h46; #100;
A = 8'h71; B = 8'h47; #100;
A = 8'h71; B = 8'h48; #100;
A = 8'h71; B = 8'h49; #100;
A = 8'h71; B = 8'h4A; #100;
A = 8'h71; B = 8'h4B; #100;
A = 8'h71; B = 8'h4C; #100;
A = 8'h71; B = 8'h4D; #100;
A = 8'h71; B = 8'h4E; #100;
A = 8'h71; B = 8'h4F; #100;
A = 8'h71; B = 8'h50; #100;
A = 8'h71; B = 8'h51; #100;
A = 8'h71; B = 8'h52; #100;
A = 8'h71; B = 8'h53; #100;
A = 8'h71; B = 8'h54; #100;
A = 8'h71; B = 8'h55; #100;
A = 8'h71; B = 8'h56; #100;
A = 8'h71; B = 8'h57; #100;
A = 8'h71; B = 8'h58; #100;
A = 8'h71; B = 8'h59; #100;
A = 8'h71; B = 8'h5A; #100;
A = 8'h71; B = 8'h5B; #100;
A = 8'h71; B = 8'h5C; #100;
A = 8'h71; B = 8'h5D; #100;
A = 8'h71; B = 8'h5E; #100;
A = 8'h71; B = 8'h5F; #100;
A = 8'h71; B = 8'h60; #100;
A = 8'h71; B = 8'h61; #100;
A = 8'h71; B = 8'h62; #100;
A = 8'h71; B = 8'h63; #100;
A = 8'h71; B = 8'h64; #100;
A = 8'h71; B = 8'h65; #100;
A = 8'h71; B = 8'h66; #100;
A = 8'h71; B = 8'h67; #100;
A = 8'h71; B = 8'h68; #100;
A = 8'h71; B = 8'h69; #100;
A = 8'h71; B = 8'h6A; #100;
A = 8'h71; B = 8'h6B; #100;
A = 8'h71; B = 8'h6C; #100;
A = 8'h71; B = 8'h6D; #100;
A = 8'h71; B = 8'h6E; #100;
A = 8'h71; B = 8'h6F; #100;
A = 8'h71; B = 8'h70; #100;
A = 8'h71; B = 8'h71; #100;
A = 8'h71; B = 8'h72; #100;
A = 8'h71; B = 8'h73; #100;
A = 8'h71; B = 8'h74; #100;
A = 8'h71; B = 8'h75; #100;
A = 8'h71; B = 8'h76; #100;
A = 8'h71; B = 8'h77; #100;
A = 8'h71; B = 8'h78; #100;
A = 8'h71; B = 8'h79; #100;
A = 8'h71; B = 8'h7A; #100;
A = 8'h71; B = 8'h7B; #100;
A = 8'h71; B = 8'h7C; #100;
A = 8'h71; B = 8'h7D; #100;
A = 8'h71; B = 8'h7E; #100;
A = 8'h71; B = 8'h7F; #100;
A = 8'h71; B = 8'h80; #100;
A = 8'h71; B = 8'h81; #100;
A = 8'h71; B = 8'h82; #100;
A = 8'h71; B = 8'h83; #100;
A = 8'h71; B = 8'h84; #100;
A = 8'h71; B = 8'h85; #100;
A = 8'h71; B = 8'h86; #100;
A = 8'h71; B = 8'h87; #100;
A = 8'h71; B = 8'h88; #100;
A = 8'h71; B = 8'h89; #100;
A = 8'h71; B = 8'h8A; #100;
A = 8'h71; B = 8'h8B; #100;
A = 8'h71; B = 8'h8C; #100;
A = 8'h71; B = 8'h8D; #100;
A = 8'h71; B = 8'h8E; #100;
A = 8'h71; B = 8'h8F; #100;
A = 8'h71; B = 8'h90; #100;
A = 8'h71; B = 8'h91; #100;
A = 8'h71; B = 8'h92; #100;
A = 8'h71; B = 8'h93; #100;
A = 8'h71; B = 8'h94; #100;
A = 8'h71; B = 8'h95; #100;
A = 8'h71; B = 8'h96; #100;
A = 8'h71; B = 8'h97; #100;
A = 8'h71; B = 8'h98; #100;
A = 8'h71; B = 8'h99; #100;
A = 8'h71; B = 8'h9A; #100;
A = 8'h71; B = 8'h9B; #100;
A = 8'h71; B = 8'h9C; #100;
A = 8'h71; B = 8'h9D; #100;
A = 8'h71; B = 8'h9E; #100;
A = 8'h71; B = 8'h9F; #100;
A = 8'h71; B = 8'hA0; #100;
A = 8'h71; B = 8'hA1; #100;
A = 8'h71; B = 8'hA2; #100;
A = 8'h71; B = 8'hA3; #100;
A = 8'h71; B = 8'hA4; #100;
A = 8'h71; B = 8'hA5; #100;
A = 8'h71; B = 8'hA6; #100;
A = 8'h71; B = 8'hA7; #100;
A = 8'h71; B = 8'hA8; #100;
A = 8'h71; B = 8'hA9; #100;
A = 8'h71; B = 8'hAA; #100;
A = 8'h71; B = 8'hAB; #100;
A = 8'h71; B = 8'hAC; #100;
A = 8'h71; B = 8'hAD; #100;
A = 8'h71; B = 8'hAE; #100;
A = 8'h71; B = 8'hAF; #100;
A = 8'h71; B = 8'hB0; #100;
A = 8'h71; B = 8'hB1; #100;
A = 8'h71; B = 8'hB2; #100;
A = 8'h71; B = 8'hB3; #100;
A = 8'h71; B = 8'hB4; #100;
A = 8'h71; B = 8'hB5; #100;
A = 8'h71; B = 8'hB6; #100;
A = 8'h71; B = 8'hB7; #100;
A = 8'h71; B = 8'hB8; #100;
A = 8'h71; B = 8'hB9; #100;
A = 8'h71; B = 8'hBA; #100;
A = 8'h71; B = 8'hBB; #100;
A = 8'h71; B = 8'hBC; #100;
A = 8'h71; B = 8'hBD; #100;
A = 8'h71; B = 8'hBE; #100;
A = 8'h71; B = 8'hBF; #100;
A = 8'h71; B = 8'hC0; #100;
A = 8'h71; B = 8'hC1; #100;
A = 8'h71; B = 8'hC2; #100;
A = 8'h71; B = 8'hC3; #100;
A = 8'h71; B = 8'hC4; #100;
A = 8'h71; B = 8'hC5; #100;
A = 8'h71; B = 8'hC6; #100;
A = 8'h71; B = 8'hC7; #100;
A = 8'h71; B = 8'hC8; #100;
A = 8'h71; B = 8'hC9; #100;
A = 8'h71; B = 8'hCA; #100;
A = 8'h71; B = 8'hCB; #100;
A = 8'h71; B = 8'hCC; #100;
A = 8'h71; B = 8'hCD; #100;
A = 8'h71; B = 8'hCE; #100;
A = 8'h71; B = 8'hCF; #100;
A = 8'h71; B = 8'hD0; #100;
A = 8'h71; B = 8'hD1; #100;
A = 8'h71; B = 8'hD2; #100;
A = 8'h71; B = 8'hD3; #100;
A = 8'h71; B = 8'hD4; #100;
A = 8'h71; B = 8'hD5; #100;
A = 8'h71; B = 8'hD6; #100;
A = 8'h71; B = 8'hD7; #100;
A = 8'h71; B = 8'hD8; #100;
A = 8'h71; B = 8'hD9; #100;
A = 8'h71; B = 8'hDA; #100;
A = 8'h71; B = 8'hDB; #100;
A = 8'h71; B = 8'hDC; #100;
A = 8'h71; B = 8'hDD; #100;
A = 8'h71; B = 8'hDE; #100;
A = 8'h71; B = 8'hDF; #100;
A = 8'h71; B = 8'hE0; #100;
A = 8'h71; B = 8'hE1; #100;
A = 8'h71; B = 8'hE2; #100;
A = 8'h71; B = 8'hE3; #100;
A = 8'h71; B = 8'hE4; #100;
A = 8'h71; B = 8'hE5; #100;
A = 8'h71; B = 8'hE6; #100;
A = 8'h71; B = 8'hE7; #100;
A = 8'h71; B = 8'hE8; #100;
A = 8'h71; B = 8'hE9; #100;
A = 8'h71; B = 8'hEA; #100;
A = 8'h71; B = 8'hEB; #100;
A = 8'h71; B = 8'hEC; #100;
A = 8'h71; B = 8'hED; #100;
A = 8'h71; B = 8'hEE; #100;
A = 8'h71; B = 8'hEF; #100;
A = 8'h71; B = 8'hF0; #100;
A = 8'h71; B = 8'hF1; #100;
A = 8'h71; B = 8'hF2; #100;
A = 8'h71; B = 8'hF3; #100;
A = 8'h71; B = 8'hF4; #100;
A = 8'h71; B = 8'hF5; #100;
A = 8'h71; B = 8'hF6; #100;
A = 8'h71; B = 8'hF7; #100;
A = 8'h71; B = 8'hF8; #100;
A = 8'h71; B = 8'hF9; #100;
A = 8'h71; B = 8'hFA; #100;
A = 8'h71; B = 8'hFB; #100;
A = 8'h71; B = 8'hFC; #100;
A = 8'h71; B = 8'hFD; #100;
A = 8'h71; B = 8'hFE; #100;
A = 8'h71; B = 8'hFF; #100;
A = 8'h72; B = 8'h0; #100;
A = 8'h72; B = 8'h1; #100;
A = 8'h72; B = 8'h2; #100;
A = 8'h72; B = 8'h3; #100;
A = 8'h72; B = 8'h4; #100;
A = 8'h72; B = 8'h5; #100;
A = 8'h72; B = 8'h6; #100;
A = 8'h72; B = 8'h7; #100;
A = 8'h72; B = 8'h8; #100;
A = 8'h72; B = 8'h9; #100;
A = 8'h72; B = 8'hA; #100;
A = 8'h72; B = 8'hB; #100;
A = 8'h72; B = 8'hC; #100;
A = 8'h72; B = 8'hD; #100;
A = 8'h72; B = 8'hE; #100;
A = 8'h72; B = 8'hF; #100;
A = 8'h72; B = 8'h10; #100;
A = 8'h72; B = 8'h11; #100;
A = 8'h72; B = 8'h12; #100;
A = 8'h72; B = 8'h13; #100;
A = 8'h72; B = 8'h14; #100;
A = 8'h72; B = 8'h15; #100;
A = 8'h72; B = 8'h16; #100;
A = 8'h72; B = 8'h17; #100;
A = 8'h72; B = 8'h18; #100;
A = 8'h72; B = 8'h19; #100;
A = 8'h72; B = 8'h1A; #100;
A = 8'h72; B = 8'h1B; #100;
A = 8'h72; B = 8'h1C; #100;
A = 8'h72; B = 8'h1D; #100;
A = 8'h72; B = 8'h1E; #100;
A = 8'h72; B = 8'h1F; #100;
A = 8'h72; B = 8'h20; #100;
A = 8'h72; B = 8'h21; #100;
A = 8'h72; B = 8'h22; #100;
A = 8'h72; B = 8'h23; #100;
A = 8'h72; B = 8'h24; #100;
A = 8'h72; B = 8'h25; #100;
A = 8'h72; B = 8'h26; #100;
A = 8'h72; B = 8'h27; #100;
A = 8'h72; B = 8'h28; #100;
A = 8'h72; B = 8'h29; #100;
A = 8'h72; B = 8'h2A; #100;
A = 8'h72; B = 8'h2B; #100;
A = 8'h72; B = 8'h2C; #100;
A = 8'h72; B = 8'h2D; #100;
A = 8'h72; B = 8'h2E; #100;
A = 8'h72; B = 8'h2F; #100;
A = 8'h72; B = 8'h30; #100;
A = 8'h72; B = 8'h31; #100;
A = 8'h72; B = 8'h32; #100;
A = 8'h72; B = 8'h33; #100;
A = 8'h72; B = 8'h34; #100;
A = 8'h72; B = 8'h35; #100;
A = 8'h72; B = 8'h36; #100;
A = 8'h72; B = 8'h37; #100;
A = 8'h72; B = 8'h38; #100;
A = 8'h72; B = 8'h39; #100;
A = 8'h72; B = 8'h3A; #100;
A = 8'h72; B = 8'h3B; #100;
A = 8'h72; B = 8'h3C; #100;
A = 8'h72; B = 8'h3D; #100;
A = 8'h72; B = 8'h3E; #100;
A = 8'h72; B = 8'h3F; #100;
A = 8'h72; B = 8'h40; #100;
A = 8'h72; B = 8'h41; #100;
A = 8'h72; B = 8'h42; #100;
A = 8'h72; B = 8'h43; #100;
A = 8'h72; B = 8'h44; #100;
A = 8'h72; B = 8'h45; #100;
A = 8'h72; B = 8'h46; #100;
A = 8'h72; B = 8'h47; #100;
A = 8'h72; B = 8'h48; #100;
A = 8'h72; B = 8'h49; #100;
A = 8'h72; B = 8'h4A; #100;
A = 8'h72; B = 8'h4B; #100;
A = 8'h72; B = 8'h4C; #100;
A = 8'h72; B = 8'h4D; #100;
A = 8'h72; B = 8'h4E; #100;
A = 8'h72; B = 8'h4F; #100;
A = 8'h72; B = 8'h50; #100;
A = 8'h72; B = 8'h51; #100;
A = 8'h72; B = 8'h52; #100;
A = 8'h72; B = 8'h53; #100;
A = 8'h72; B = 8'h54; #100;
A = 8'h72; B = 8'h55; #100;
A = 8'h72; B = 8'h56; #100;
A = 8'h72; B = 8'h57; #100;
A = 8'h72; B = 8'h58; #100;
A = 8'h72; B = 8'h59; #100;
A = 8'h72; B = 8'h5A; #100;
A = 8'h72; B = 8'h5B; #100;
A = 8'h72; B = 8'h5C; #100;
A = 8'h72; B = 8'h5D; #100;
A = 8'h72; B = 8'h5E; #100;
A = 8'h72; B = 8'h5F; #100;
A = 8'h72; B = 8'h60; #100;
A = 8'h72; B = 8'h61; #100;
A = 8'h72; B = 8'h62; #100;
A = 8'h72; B = 8'h63; #100;
A = 8'h72; B = 8'h64; #100;
A = 8'h72; B = 8'h65; #100;
A = 8'h72; B = 8'h66; #100;
A = 8'h72; B = 8'h67; #100;
A = 8'h72; B = 8'h68; #100;
A = 8'h72; B = 8'h69; #100;
A = 8'h72; B = 8'h6A; #100;
A = 8'h72; B = 8'h6B; #100;
A = 8'h72; B = 8'h6C; #100;
A = 8'h72; B = 8'h6D; #100;
A = 8'h72; B = 8'h6E; #100;
A = 8'h72; B = 8'h6F; #100;
A = 8'h72; B = 8'h70; #100;
A = 8'h72; B = 8'h71; #100;
A = 8'h72; B = 8'h72; #100;
A = 8'h72; B = 8'h73; #100;
A = 8'h72; B = 8'h74; #100;
A = 8'h72; B = 8'h75; #100;
A = 8'h72; B = 8'h76; #100;
A = 8'h72; B = 8'h77; #100;
A = 8'h72; B = 8'h78; #100;
A = 8'h72; B = 8'h79; #100;
A = 8'h72; B = 8'h7A; #100;
A = 8'h72; B = 8'h7B; #100;
A = 8'h72; B = 8'h7C; #100;
A = 8'h72; B = 8'h7D; #100;
A = 8'h72; B = 8'h7E; #100;
A = 8'h72; B = 8'h7F; #100;
A = 8'h72; B = 8'h80; #100;
A = 8'h72; B = 8'h81; #100;
A = 8'h72; B = 8'h82; #100;
A = 8'h72; B = 8'h83; #100;
A = 8'h72; B = 8'h84; #100;
A = 8'h72; B = 8'h85; #100;
A = 8'h72; B = 8'h86; #100;
A = 8'h72; B = 8'h87; #100;
A = 8'h72; B = 8'h88; #100;
A = 8'h72; B = 8'h89; #100;
A = 8'h72; B = 8'h8A; #100;
A = 8'h72; B = 8'h8B; #100;
A = 8'h72; B = 8'h8C; #100;
A = 8'h72; B = 8'h8D; #100;
A = 8'h72; B = 8'h8E; #100;
A = 8'h72; B = 8'h8F; #100;
A = 8'h72; B = 8'h90; #100;
A = 8'h72; B = 8'h91; #100;
A = 8'h72; B = 8'h92; #100;
A = 8'h72; B = 8'h93; #100;
A = 8'h72; B = 8'h94; #100;
A = 8'h72; B = 8'h95; #100;
A = 8'h72; B = 8'h96; #100;
A = 8'h72; B = 8'h97; #100;
A = 8'h72; B = 8'h98; #100;
A = 8'h72; B = 8'h99; #100;
A = 8'h72; B = 8'h9A; #100;
A = 8'h72; B = 8'h9B; #100;
A = 8'h72; B = 8'h9C; #100;
A = 8'h72; B = 8'h9D; #100;
A = 8'h72; B = 8'h9E; #100;
A = 8'h72; B = 8'h9F; #100;
A = 8'h72; B = 8'hA0; #100;
A = 8'h72; B = 8'hA1; #100;
A = 8'h72; B = 8'hA2; #100;
A = 8'h72; B = 8'hA3; #100;
A = 8'h72; B = 8'hA4; #100;
A = 8'h72; B = 8'hA5; #100;
A = 8'h72; B = 8'hA6; #100;
A = 8'h72; B = 8'hA7; #100;
A = 8'h72; B = 8'hA8; #100;
A = 8'h72; B = 8'hA9; #100;
A = 8'h72; B = 8'hAA; #100;
A = 8'h72; B = 8'hAB; #100;
A = 8'h72; B = 8'hAC; #100;
A = 8'h72; B = 8'hAD; #100;
A = 8'h72; B = 8'hAE; #100;
A = 8'h72; B = 8'hAF; #100;
A = 8'h72; B = 8'hB0; #100;
A = 8'h72; B = 8'hB1; #100;
A = 8'h72; B = 8'hB2; #100;
A = 8'h72; B = 8'hB3; #100;
A = 8'h72; B = 8'hB4; #100;
A = 8'h72; B = 8'hB5; #100;
A = 8'h72; B = 8'hB6; #100;
A = 8'h72; B = 8'hB7; #100;
A = 8'h72; B = 8'hB8; #100;
A = 8'h72; B = 8'hB9; #100;
A = 8'h72; B = 8'hBA; #100;
A = 8'h72; B = 8'hBB; #100;
A = 8'h72; B = 8'hBC; #100;
A = 8'h72; B = 8'hBD; #100;
A = 8'h72; B = 8'hBE; #100;
A = 8'h72; B = 8'hBF; #100;
A = 8'h72; B = 8'hC0; #100;
A = 8'h72; B = 8'hC1; #100;
A = 8'h72; B = 8'hC2; #100;
A = 8'h72; B = 8'hC3; #100;
A = 8'h72; B = 8'hC4; #100;
A = 8'h72; B = 8'hC5; #100;
A = 8'h72; B = 8'hC6; #100;
A = 8'h72; B = 8'hC7; #100;
A = 8'h72; B = 8'hC8; #100;
A = 8'h72; B = 8'hC9; #100;
A = 8'h72; B = 8'hCA; #100;
A = 8'h72; B = 8'hCB; #100;
A = 8'h72; B = 8'hCC; #100;
A = 8'h72; B = 8'hCD; #100;
A = 8'h72; B = 8'hCE; #100;
A = 8'h72; B = 8'hCF; #100;
A = 8'h72; B = 8'hD0; #100;
A = 8'h72; B = 8'hD1; #100;
A = 8'h72; B = 8'hD2; #100;
A = 8'h72; B = 8'hD3; #100;
A = 8'h72; B = 8'hD4; #100;
A = 8'h72; B = 8'hD5; #100;
A = 8'h72; B = 8'hD6; #100;
A = 8'h72; B = 8'hD7; #100;
A = 8'h72; B = 8'hD8; #100;
A = 8'h72; B = 8'hD9; #100;
A = 8'h72; B = 8'hDA; #100;
A = 8'h72; B = 8'hDB; #100;
A = 8'h72; B = 8'hDC; #100;
A = 8'h72; B = 8'hDD; #100;
A = 8'h72; B = 8'hDE; #100;
A = 8'h72; B = 8'hDF; #100;
A = 8'h72; B = 8'hE0; #100;
A = 8'h72; B = 8'hE1; #100;
A = 8'h72; B = 8'hE2; #100;
A = 8'h72; B = 8'hE3; #100;
A = 8'h72; B = 8'hE4; #100;
A = 8'h72; B = 8'hE5; #100;
A = 8'h72; B = 8'hE6; #100;
A = 8'h72; B = 8'hE7; #100;
A = 8'h72; B = 8'hE8; #100;
A = 8'h72; B = 8'hE9; #100;
A = 8'h72; B = 8'hEA; #100;
A = 8'h72; B = 8'hEB; #100;
A = 8'h72; B = 8'hEC; #100;
A = 8'h72; B = 8'hED; #100;
A = 8'h72; B = 8'hEE; #100;
A = 8'h72; B = 8'hEF; #100;
A = 8'h72; B = 8'hF0; #100;
A = 8'h72; B = 8'hF1; #100;
A = 8'h72; B = 8'hF2; #100;
A = 8'h72; B = 8'hF3; #100;
A = 8'h72; B = 8'hF4; #100;
A = 8'h72; B = 8'hF5; #100;
A = 8'h72; B = 8'hF6; #100;
A = 8'h72; B = 8'hF7; #100;
A = 8'h72; B = 8'hF8; #100;
A = 8'h72; B = 8'hF9; #100;
A = 8'h72; B = 8'hFA; #100;
A = 8'h72; B = 8'hFB; #100;
A = 8'h72; B = 8'hFC; #100;
A = 8'h72; B = 8'hFD; #100;
A = 8'h72; B = 8'hFE; #100;
A = 8'h72; B = 8'hFF; #100;
A = 8'h73; B = 8'h0; #100;
A = 8'h73; B = 8'h1; #100;
A = 8'h73; B = 8'h2; #100;
A = 8'h73; B = 8'h3; #100;
A = 8'h73; B = 8'h4; #100;
A = 8'h73; B = 8'h5; #100;
A = 8'h73; B = 8'h6; #100;
A = 8'h73; B = 8'h7; #100;
A = 8'h73; B = 8'h8; #100;
A = 8'h73; B = 8'h9; #100;
A = 8'h73; B = 8'hA; #100;
A = 8'h73; B = 8'hB; #100;
A = 8'h73; B = 8'hC; #100;
A = 8'h73; B = 8'hD; #100;
A = 8'h73; B = 8'hE; #100;
A = 8'h73; B = 8'hF; #100;
A = 8'h73; B = 8'h10; #100;
A = 8'h73; B = 8'h11; #100;
A = 8'h73; B = 8'h12; #100;
A = 8'h73; B = 8'h13; #100;
A = 8'h73; B = 8'h14; #100;
A = 8'h73; B = 8'h15; #100;
A = 8'h73; B = 8'h16; #100;
A = 8'h73; B = 8'h17; #100;
A = 8'h73; B = 8'h18; #100;
A = 8'h73; B = 8'h19; #100;
A = 8'h73; B = 8'h1A; #100;
A = 8'h73; B = 8'h1B; #100;
A = 8'h73; B = 8'h1C; #100;
A = 8'h73; B = 8'h1D; #100;
A = 8'h73; B = 8'h1E; #100;
A = 8'h73; B = 8'h1F; #100;
A = 8'h73; B = 8'h20; #100;
A = 8'h73; B = 8'h21; #100;
A = 8'h73; B = 8'h22; #100;
A = 8'h73; B = 8'h23; #100;
A = 8'h73; B = 8'h24; #100;
A = 8'h73; B = 8'h25; #100;
A = 8'h73; B = 8'h26; #100;
A = 8'h73; B = 8'h27; #100;
A = 8'h73; B = 8'h28; #100;
A = 8'h73; B = 8'h29; #100;
A = 8'h73; B = 8'h2A; #100;
A = 8'h73; B = 8'h2B; #100;
A = 8'h73; B = 8'h2C; #100;
A = 8'h73; B = 8'h2D; #100;
A = 8'h73; B = 8'h2E; #100;
A = 8'h73; B = 8'h2F; #100;
A = 8'h73; B = 8'h30; #100;
A = 8'h73; B = 8'h31; #100;
A = 8'h73; B = 8'h32; #100;
A = 8'h73; B = 8'h33; #100;
A = 8'h73; B = 8'h34; #100;
A = 8'h73; B = 8'h35; #100;
A = 8'h73; B = 8'h36; #100;
A = 8'h73; B = 8'h37; #100;
A = 8'h73; B = 8'h38; #100;
A = 8'h73; B = 8'h39; #100;
A = 8'h73; B = 8'h3A; #100;
A = 8'h73; B = 8'h3B; #100;
A = 8'h73; B = 8'h3C; #100;
A = 8'h73; B = 8'h3D; #100;
A = 8'h73; B = 8'h3E; #100;
A = 8'h73; B = 8'h3F; #100;
A = 8'h73; B = 8'h40; #100;
A = 8'h73; B = 8'h41; #100;
A = 8'h73; B = 8'h42; #100;
A = 8'h73; B = 8'h43; #100;
A = 8'h73; B = 8'h44; #100;
A = 8'h73; B = 8'h45; #100;
A = 8'h73; B = 8'h46; #100;
A = 8'h73; B = 8'h47; #100;
A = 8'h73; B = 8'h48; #100;
A = 8'h73; B = 8'h49; #100;
A = 8'h73; B = 8'h4A; #100;
A = 8'h73; B = 8'h4B; #100;
A = 8'h73; B = 8'h4C; #100;
A = 8'h73; B = 8'h4D; #100;
A = 8'h73; B = 8'h4E; #100;
A = 8'h73; B = 8'h4F; #100;
A = 8'h73; B = 8'h50; #100;
A = 8'h73; B = 8'h51; #100;
A = 8'h73; B = 8'h52; #100;
A = 8'h73; B = 8'h53; #100;
A = 8'h73; B = 8'h54; #100;
A = 8'h73; B = 8'h55; #100;
A = 8'h73; B = 8'h56; #100;
A = 8'h73; B = 8'h57; #100;
A = 8'h73; B = 8'h58; #100;
A = 8'h73; B = 8'h59; #100;
A = 8'h73; B = 8'h5A; #100;
A = 8'h73; B = 8'h5B; #100;
A = 8'h73; B = 8'h5C; #100;
A = 8'h73; B = 8'h5D; #100;
A = 8'h73; B = 8'h5E; #100;
A = 8'h73; B = 8'h5F; #100;
A = 8'h73; B = 8'h60; #100;
A = 8'h73; B = 8'h61; #100;
A = 8'h73; B = 8'h62; #100;
A = 8'h73; B = 8'h63; #100;
A = 8'h73; B = 8'h64; #100;
A = 8'h73; B = 8'h65; #100;
A = 8'h73; B = 8'h66; #100;
A = 8'h73; B = 8'h67; #100;
A = 8'h73; B = 8'h68; #100;
A = 8'h73; B = 8'h69; #100;
A = 8'h73; B = 8'h6A; #100;
A = 8'h73; B = 8'h6B; #100;
A = 8'h73; B = 8'h6C; #100;
A = 8'h73; B = 8'h6D; #100;
A = 8'h73; B = 8'h6E; #100;
A = 8'h73; B = 8'h6F; #100;
A = 8'h73; B = 8'h70; #100;
A = 8'h73; B = 8'h71; #100;
A = 8'h73; B = 8'h72; #100;
A = 8'h73; B = 8'h73; #100;
A = 8'h73; B = 8'h74; #100;
A = 8'h73; B = 8'h75; #100;
A = 8'h73; B = 8'h76; #100;
A = 8'h73; B = 8'h77; #100;
A = 8'h73; B = 8'h78; #100;
A = 8'h73; B = 8'h79; #100;
A = 8'h73; B = 8'h7A; #100;
A = 8'h73; B = 8'h7B; #100;
A = 8'h73; B = 8'h7C; #100;
A = 8'h73; B = 8'h7D; #100;
A = 8'h73; B = 8'h7E; #100;
A = 8'h73; B = 8'h7F; #100;
A = 8'h73; B = 8'h80; #100;
A = 8'h73; B = 8'h81; #100;
A = 8'h73; B = 8'h82; #100;
A = 8'h73; B = 8'h83; #100;
A = 8'h73; B = 8'h84; #100;
A = 8'h73; B = 8'h85; #100;
A = 8'h73; B = 8'h86; #100;
A = 8'h73; B = 8'h87; #100;
A = 8'h73; B = 8'h88; #100;
A = 8'h73; B = 8'h89; #100;
A = 8'h73; B = 8'h8A; #100;
A = 8'h73; B = 8'h8B; #100;
A = 8'h73; B = 8'h8C; #100;
A = 8'h73; B = 8'h8D; #100;
A = 8'h73; B = 8'h8E; #100;
A = 8'h73; B = 8'h8F; #100;
A = 8'h73; B = 8'h90; #100;
A = 8'h73; B = 8'h91; #100;
A = 8'h73; B = 8'h92; #100;
A = 8'h73; B = 8'h93; #100;
A = 8'h73; B = 8'h94; #100;
A = 8'h73; B = 8'h95; #100;
A = 8'h73; B = 8'h96; #100;
A = 8'h73; B = 8'h97; #100;
A = 8'h73; B = 8'h98; #100;
A = 8'h73; B = 8'h99; #100;
A = 8'h73; B = 8'h9A; #100;
A = 8'h73; B = 8'h9B; #100;
A = 8'h73; B = 8'h9C; #100;
A = 8'h73; B = 8'h9D; #100;
A = 8'h73; B = 8'h9E; #100;
A = 8'h73; B = 8'h9F; #100;
A = 8'h73; B = 8'hA0; #100;
A = 8'h73; B = 8'hA1; #100;
A = 8'h73; B = 8'hA2; #100;
A = 8'h73; B = 8'hA3; #100;
A = 8'h73; B = 8'hA4; #100;
A = 8'h73; B = 8'hA5; #100;
A = 8'h73; B = 8'hA6; #100;
A = 8'h73; B = 8'hA7; #100;
A = 8'h73; B = 8'hA8; #100;
A = 8'h73; B = 8'hA9; #100;
A = 8'h73; B = 8'hAA; #100;
A = 8'h73; B = 8'hAB; #100;
A = 8'h73; B = 8'hAC; #100;
A = 8'h73; B = 8'hAD; #100;
A = 8'h73; B = 8'hAE; #100;
A = 8'h73; B = 8'hAF; #100;
A = 8'h73; B = 8'hB0; #100;
A = 8'h73; B = 8'hB1; #100;
A = 8'h73; B = 8'hB2; #100;
A = 8'h73; B = 8'hB3; #100;
A = 8'h73; B = 8'hB4; #100;
A = 8'h73; B = 8'hB5; #100;
A = 8'h73; B = 8'hB6; #100;
A = 8'h73; B = 8'hB7; #100;
A = 8'h73; B = 8'hB8; #100;
A = 8'h73; B = 8'hB9; #100;
A = 8'h73; B = 8'hBA; #100;
A = 8'h73; B = 8'hBB; #100;
A = 8'h73; B = 8'hBC; #100;
A = 8'h73; B = 8'hBD; #100;
A = 8'h73; B = 8'hBE; #100;
A = 8'h73; B = 8'hBF; #100;
A = 8'h73; B = 8'hC0; #100;
A = 8'h73; B = 8'hC1; #100;
A = 8'h73; B = 8'hC2; #100;
A = 8'h73; B = 8'hC3; #100;
A = 8'h73; B = 8'hC4; #100;
A = 8'h73; B = 8'hC5; #100;
A = 8'h73; B = 8'hC6; #100;
A = 8'h73; B = 8'hC7; #100;
A = 8'h73; B = 8'hC8; #100;
A = 8'h73; B = 8'hC9; #100;
A = 8'h73; B = 8'hCA; #100;
A = 8'h73; B = 8'hCB; #100;
A = 8'h73; B = 8'hCC; #100;
A = 8'h73; B = 8'hCD; #100;
A = 8'h73; B = 8'hCE; #100;
A = 8'h73; B = 8'hCF; #100;
A = 8'h73; B = 8'hD0; #100;
A = 8'h73; B = 8'hD1; #100;
A = 8'h73; B = 8'hD2; #100;
A = 8'h73; B = 8'hD3; #100;
A = 8'h73; B = 8'hD4; #100;
A = 8'h73; B = 8'hD5; #100;
A = 8'h73; B = 8'hD6; #100;
A = 8'h73; B = 8'hD7; #100;
A = 8'h73; B = 8'hD8; #100;
A = 8'h73; B = 8'hD9; #100;
A = 8'h73; B = 8'hDA; #100;
A = 8'h73; B = 8'hDB; #100;
A = 8'h73; B = 8'hDC; #100;
A = 8'h73; B = 8'hDD; #100;
A = 8'h73; B = 8'hDE; #100;
A = 8'h73; B = 8'hDF; #100;
A = 8'h73; B = 8'hE0; #100;
A = 8'h73; B = 8'hE1; #100;
A = 8'h73; B = 8'hE2; #100;
A = 8'h73; B = 8'hE3; #100;
A = 8'h73; B = 8'hE4; #100;
A = 8'h73; B = 8'hE5; #100;
A = 8'h73; B = 8'hE6; #100;
A = 8'h73; B = 8'hE7; #100;
A = 8'h73; B = 8'hE8; #100;
A = 8'h73; B = 8'hE9; #100;
A = 8'h73; B = 8'hEA; #100;
A = 8'h73; B = 8'hEB; #100;
A = 8'h73; B = 8'hEC; #100;
A = 8'h73; B = 8'hED; #100;
A = 8'h73; B = 8'hEE; #100;
A = 8'h73; B = 8'hEF; #100;
A = 8'h73; B = 8'hF0; #100;
A = 8'h73; B = 8'hF1; #100;
A = 8'h73; B = 8'hF2; #100;
A = 8'h73; B = 8'hF3; #100;
A = 8'h73; B = 8'hF4; #100;
A = 8'h73; B = 8'hF5; #100;
A = 8'h73; B = 8'hF6; #100;
A = 8'h73; B = 8'hF7; #100;
A = 8'h73; B = 8'hF8; #100;
A = 8'h73; B = 8'hF9; #100;
A = 8'h73; B = 8'hFA; #100;
A = 8'h73; B = 8'hFB; #100;
A = 8'h73; B = 8'hFC; #100;
A = 8'h73; B = 8'hFD; #100;
A = 8'h73; B = 8'hFE; #100;
A = 8'h73; B = 8'hFF; #100;
A = 8'h74; B = 8'h0; #100;
A = 8'h74; B = 8'h1; #100;
A = 8'h74; B = 8'h2; #100;
A = 8'h74; B = 8'h3; #100;
A = 8'h74; B = 8'h4; #100;
A = 8'h74; B = 8'h5; #100;
A = 8'h74; B = 8'h6; #100;
A = 8'h74; B = 8'h7; #100;
A = 8'h74; B = 8'h8; #100;
A = 8'h74; B = 8'h9; #100;
A = 8'h74; B = 8'hA; #100;
A = 8'h74; B = 8'hB; #100;
A = 8'h74; B = 8'hC; #100;
A = 8'h74; B = 8'hD; #100;
A = 8'h74; B = 8'hE; #100;
A = 8'h74; B = 8'hF; #100;
A = 8'h74; B = 8'h10; #100;
A = 8'h74; B = 8'h11; #100;
A = 8'h74; B = 8'h12; #100;
A = 8'h74; B = 8'h13; #100;
A = 8'h74; B = 8'h14; #100;
A = 8'h74; B = 8'h15; #100;
A = 8'h74; B = 8'h16; #100;
A = 8'h74; B = 8'h17; #100;
A = 8'h74; B = 8'h18; #100;
A = 8'h74; B = 8'h19; #100;
A = 8'h74; B = 8'h1A; #100;
A = 8'h74; B = 8'h1B; #100;
A = 8'h74; B = 8'h1C; #100;
A = 8'h74; B = 8'h1D; #100;
A = 8'h74; B = 8'h1E; #100;
A = 8'h74; B = 8'h1F; #100;
A = 8'h74; B = 8'h20; #100;
A = 8'h74; B = 8'h21; #100;
A = 8'h74; B = 8'h22; #100;
A = 8'h74; B = 8'h23; #100;
A = 8'h74; B = 8'h24; #100;
A = 8'h74; B = 8'h25; #100;
A = 8'h74; B = 8'h26; #100;
A = 8'h74; B = 8'h27; #100;
A = 8'h74; B = 8'h28; #100;
A = 8'h74; B = 8'h29; #100;
A = 8'h74; B = 8'h2A; #100;
A = 8'h74; B = 8'h2B; #100;
A = 8'h74; B = 8'h2C; #100;
A = 8'h74; B = 8'h2D; #100;
A = 8'h74; B = 8'h2E; #100;
A = 8'h74; B = 8'h2F; #100;
A = 8'h74; B = 8'h30; #100;
A = 8'h74; B = 8'h31; #100;
A = 8'h74; B = 8'h32; #100;
A = 8'h74; B = 8'h33; #100;
A = 8'h74; B = 8'h34; #100;
A = 8'h74; B = 8'h35; #100;
A = 8'h74; B = 8'h36; #100;
A = 8'h74; B = 8'h37; #100;
A = 8'h74; B = 8'h38; #100;
A = 8'h74; B = 8'h39; #100;
A = 8'h74; B = 8'h3A; #100;
A = 8'h74; B = 8'h3B; #100;
A = 8'h74; B = 8'h3C; #100;
A = 8'h74; B = 8'h3D; #100;
A = 8'h74; B = 8'h3E; #100;
A = 8'h74; B = 8'h3F; #100;
A = 8'h74; B = 8'h40; #100;
A = 8'h74; B = 8'h41; #100;
A = 8'h74; B = 8'h42; #100;
A = 8'h74; B = 8'h43; #100;
A = 8'h74; B = 8'h44; #100;
A = 8'h74; B = 8'h45; #100;
A = 8'h74; B = 8'h46; #100;
A = 8'h74; B = 8'h47; #100;
A = 8'h74; B = 8'h48; #100;
A = 8'h74; B = 8'h49; #100;
A = 8'h74; B = 8'h4A; #100;
A = 8'h74; B = 8'h4B; #100;
A = 8'h74; B = 8'h4C; #100;
A = 8'h74; B = 8'h4D; #100;
A = 8'h74; B = 8'h4E; #100;
A = 8'h74; B = 8'h4F; #100;
A = 8'h74; B = 8'h50; #100;
A = 8'h74; B = 8'h51; #100;
A = 8'h74; B = 8'h52; #100;
A = 8'h74; B = 8'h53; #100;
A = 8'h74; B = 8'h54; #100;
A = 8'h74; B = 8'h55; #100;
A = 8'h74; B = 8'h56; #100;
A = 8'h74; B = 8'h57; #100;
A = 8'h74; B = 8'h58; #100;
A = 8'h74; B = 8'h59; #100;
A = 8'h74; B = 8'h5A; #100;
A = 8'h74; B = 8'h5B; #100;
A = 8'h74; B = 8'h5C; #100;
A = 8'h74; B = 8'h5D; #100;
A = 8'h74; B = 8'h5E; #100;
A = 8'h74; B = 8'h5F; #100;
A = 8'h74; B = 8'h60; #100;
A = 8'h74; B = 8'h61; #100;
A = 8'h74; B = 8'h62; #100;
A = 8'h74; B = 8'h63; #100;
A = 8'h74; B = 8'h64; #100;
A = 8'h74; B = 8'h65; #100;
A = 8'h74; B = 8'h66; #100;
A = 8'h74; B = 8'h67; #100;
A = 8'h74; B = 8'h68; #100;
A = 8'h74; B = 8'h69; #100;
A = 8'h74; B = 8'h6A; #100;
A = 8'h74; B = 8'h6B; #100;
A = 8'h74; B = 8'h6C; #100;
A = 8'h74; B = 8'h6D; #100;
A = 8'h74; B = 8'h6E; #100;
A = 8'h74; B = 8'h6F; #100;
A = 8'h74; B = 8'h70; #100;
A = 8'h74; B = 8'h71; #100;
A = 8'h74; B = 8'h72; #100;
A = 8'h74; B = 8'h73; #100;
A = 8'h74; B = 8'h74; #100;
A = 8'h74; B = 8'h75; #100;
A = 8'h74; B = 8'h76; #100;
A = 8'h74; B = 8'h77; #100;
A = 8'h74; B = 8'h78; #100;
A = 8'h74; B = 8'h79; #100;
A = 8'h74; B = 8'h7A; #100;
A = 8'h74; B = 8'h7B; #100;
A = 8'h74; B = 8'h7C; #100;
A = 8'h74; B = 8'h7D; #100;
A = 8'h74; B = 8'h7E; #100;
A = 8'h74; B = 8'h7F; #100;
A = 8'h74; B = 8'h80; #100;
A = 8'h74; B = 8'h81; #100;
A = 8'h74; B = 8'h82; #100;
A = 8'h74; B = 8'h83; #100;
A = 8'h74; B = 8'h84; #100;
A = 8'h74; B = 8'h85; #100;
A = 8'h74; B = 8'h86; #100;
A = 8'h74; B = 8'h87; #100;
A = 8'h74; B = 8'h88; #100;
A = 8'h74; B = 8'h89; #100;
A = 8'h74; B = 8'h8A; #100;
A = 8'h74; B = 8'h8B; #100;
A = 8'h74; B = 8'h8C; #100;
A = 8'h74; B = 8'h8D; #100;
A = 8'h74; B = 8'h8E; #100;
A = 8'h74; B = 8'h8F; #100;
A = 8'h74; B = 8'h90; #100;
A = 8'h74; B = 8'h91; #100;
A = 8'h74; B = 8'h92; #100;
A = 8'h74; B = 8'h93; #100;
A = 8'h74; B = 8'h94; #100;
A = 8'h74; B = 8'h95; #100;
A = 8'h74; B = 8'h96; #100;
A = 8'h74; B = 8'h97; #100;
A = 8'h74; B = 8'h98; #100;
A = 8'h74; B = 8'h99; #100;
A = 8'h74; B = 8'h9A; #100;
A = 8'h74; B = 8'h9B; #100;
A = 8'h74; B = 8'h9C; #100;
A = 8'h74; B = 8'h9D; #100;
A = 8'h74; B = 8'h9E; #100;
A = 8'h74; B = 8'h9F; #100;
A = 8'h74; B = 8'hA0; #100;
A = 8'h74; B = 8'hA1; #100;
A = 8'h74; B = 8'hA2; #100;
A = 8'h74; B = 8'hA3; #100;
A = 8'h74; B = 8'hA4; #100;
A = 8'h74; B = 8'hA5; #100;
A = 8'h74; B = 8'hA6; #100;
A = 8'h74; B = 8'hA7; #100;
A = 8'h74; B = 8'hA8; #100;
A = 8'h74; B = 8'hA9; #100;
A = 8'h74; B = 8'hAA; #100;
A = 8'h74; B = 8'hAB; #100;
A = 8'h74; B = 8'hAC; #100;
A = 8'h74; B = 8'hAD; #100;
A = 8'h74; B = 8'hAE; #100;
A = 8'h74; B = 8'hAF; #100;
A = 8'h74; B = 8'hB0; #100;
A = 8'h74; B = 8'hB1; #100;
A = 8'h74; B = 8'hB2; #100;
A = 8'h74; B = 8'hB3; #100;
A = 8'h74; B = 8'hB4; #100;
A = 8'h74; B = 8'hB5; #100;
A = 8'h74; B = 8'hB6; #100;
A = 8'h74; B = 8'hB7; #100;
A = 8'h74; B = 8'hB8; #100;
A = 8'h74; B = 8'hB9; #100;
A = 8'h74; B = 8'hBA; #100;
A = 8'h74; B = 8'hBB; #100;
A = 8'h74; B = 8'hBC; #100;
A = 8'h74; B = 8'hBD; #100;
A = 8'h74; B = 8'hBE; #100;
A = 8'h74; B = 8'hBF; #100;
A = 8'h74; B = 8'hC0; #100;
A = 8'h74; B = 8'hC1; #100;
A = 8'h74; B = 8'hC2; #100;
A = 8'h74; B = 8'hC3; #100;
A = 8'h74; B = 8'hC4; #100;
A = 8'h74; B = 8'hC5; #100;
A = 8'h74; B = 8'hC6; #100;
A = 8'h74; B = 8'hC7; #100;
A = 8'h74; B = 8'hC8; #100;
A = 8'h74; B = 8'hC9; #100;
A = 8'h74; B = 8'hCA; #100;
A = 8'h74; B = 8'hCB; #100;
A = 8'h74; B = 8'hCC; #100;
A = 8'h74; B = 8'hCD; #100;
A = 8'h74; B = 8'hCE; #100;
A = 8'h74; B = 8'hCF; #100;
A = 8'h74; B = 8'hD0; #100;
A = 8'h74; B = 8'hD1; #100;
A = 8'h74; B = 8'hD2; #100;
A = 8'h74; B = 8'hD3; #100;
A = 8'h74; B = 8'hD4; #100;
A = 8'h74; B = 8'hD5; #100;
A = 8'h74; B = 8'hD6; #100;
A = 8'h74; B = 8'hD7; #100;
A = 8'h74; B = 8'hD8; #100;
A = 8'h74; B = 8'hD9; #100;
A = 8'h74; B = 8'hDA; #100;
A = 8'h74; B = 8'hDB; #100;
A = 8'h74; B = 8'hDC; #100;
A = 8'h74; B = 8'hDD; #100;
A = 8'h74; B = 8'hDE; #100;
A = 8'h74; B = 8'hDF; #100;
A = 8'h74; B = 8'hE0; #100;
A = 8'h74; B = 8'hE1; #100;
A = 8'h74; B = 8'hE2; #100;
A = 8'h74; B = 8'hE3; #100;
A = 8'h74; B = 8'hE4; #100;
A = 8'h74; B = 8'hE5; #100;
A = 8'h74; B = 8'hE6; #100;
A = 8'h74; B = 8'hE7; #100;
A = 8'h74; B = 8'hE8; #100;
A = 8'h74; B = 8'hE9; #100;
A = 8'h74; B = 8'hEA; #100;
A = 8'h74; B = 8'hEB; #100;
A = 8'h74; B = 8'hEC; #100;
A = 8'h74; B = 8'hED; #100;
A = 8'h74; B = 8'hEE; #100;
A = 8'h74; B = 8'hEF; #100;
A = 8'h74; B = 8'hF0; #100;
A = 8'h74; B = 8'hF1; #100;
A = 8'h74; B = 8'hF2; #100;
A = 8'h74; B = 8'hF3; #100;
A = 8'h74; B = 8'hF4; #100;
A = 8'h74; B = 8'hF5; #100;
A = 8'h74; B = 8'hF6; #100;
A = 8'h74; B = 8'hF7; #100;
A = 8'h74; B = 8'hF8; #100;
A = 8'h74; B = 8'hF9; #100;
A = 8'h74; B = 8'hFA; #100;
A = 8'h74; B = 8'hFB; #100;
A = 8'h74; B = 8'hFC; #100;
A = 8'h74; B = 8'hFD; #100;
A = 8'h74; B = 8'hFE; #100;
A = 8'h74; B = 8'hFF; #100;
A = 8'h75; B = 8'h0; #100;
A = 8'h75; B = 8'h1; #100;
A = 8'h75; B = 8'h2; #100;
A = 8'h75; B = 8'h3; #100;
A = 8'h75; B = 8'h4; #100;
A = 8'h75; B = 8'h5; #100;
A = 8'h75; B = 8'h6; #100;
A = 8'h75; B = 8'h7; #100;
A = 8'h75; B = 8'h8; #100;
A = 8'h75; B = 8'h9; #100;
A = 8'h75; B = 8'hA; #100;
A = 8'h75; B = 8'hB; #100;
A = 8'h75; B = 8'hC; #100;
A = 8'h75; B = 8'hD; #100;
A = 8'h75; B = 8'hE; #100;
A = 8'h75; B = 8'hF; #100;
A = 8'h75; B = 8'h10; #100;
A = 8'h75; B = 8'h11; #100;
A = 8'h75; B = 8'h12; #100;
A = 8'h75; B = 8'h13; #100;
A = 8'h75; B = 8'h14; #100;
A = 8'h75; B = 8'h15; #100;
A = 8'h75; B = 8'h16; #100;
A = 8'h75; B = 8'h17; #100;
A = 8'h75; B = 8'h18; #100;
A = 8'h75; B = 8'h19; #100;
A = 8'h75; B = 8'h1A; #100;
A = 8'h75; B = 8'h1B; #100;
A = 8'h75; B = 8'h1C; #100;
A = 8'h75; B = 8'h1D; #100;
A = 8'h75; B = 8'h1E; #100;
A = 8'h75; B = 8'h1F; #100;
A = 8'h75; B = 8'h20; #100;
A = 8'h75; B = 8'h21; #100;
A = 8'h75; B = 8'h22; #100;
A = 8'h75; B = 8'h23; #100;
A = 8'h75; B = 8'h24; #100;
A = 8'h75; B = 8'h25; #100;
A = 8'h75; B = 8'h26; #100;
A = 8'h75; B = 8'h27; #100;
A = 8'h75; B = 8'h28; #100;
A = 8'h75; B = 8'h29; #100;
A = 8'h75; B = 8'h2A; #100;
A = 8'h75; B = 8'h2B; #100;
A = 8'h75; B = 8'h2C; #100;
A = 8'h75; B = 8'h2D; #100;
A = 8'h75; B = 8'h2E; #100;
A = 8'h75; B = 8'h2F; #100;
A = 8'h75; B = 8'h30; #100;
A = 8'h75; B = 8'h31; #100;
A = 8'h75; B = 8'h32; #100;
A = 8'h75; B = 8'h33; #100;
A = 8'h75; B = 8'h34; #100;
A = 8'h75; B = 8'h35; #100;
A = 8'h75; B = 8'h36; #100;
A = 8'h75; B = 8'h37; #100;
A = 8'h75; B = 8'h38; #100;
A = 8'h75; B = 8'h39; #100;
A = 8'h75; B = 8'h3A; #100;
A = 8'h75; B = 8'h3B; #100;
A = 8'h75; B = 8'h3C; #100;
A = 8'h75; B = 8'h3D; #100;
A = 8'h75; B = 8'h3E; #100;
A = 8'h75; B = 8'h3F; #100;
A = 8'h75; B = 8'h40; #100;
A = 8'h75; B = 8'h41; #100;
A = 8'h75; B = 8'h42; #100;
A = 8'h75; B = 8'h43; #100;
A = 8'h75; B = 8'h44; #100;
A = 8'h75; B = 8'h45; #100;
A = 8'h75; B = 8'h46; #100;
A = 8'h75; B = 8'h47; #100;
A = 8'h75; B = 8'h48; #100;
A = 8'h75; B = 8'h49; #100;
A = 8'h75; B = 8'h4A; #100;
A = 8'h75; B = 8'h4B; #100;
A = 8'h75; B = 8'h4C; #100;
A = 8'h75; B = 8'h4D; #100;
A = 8'h75; B = 8'h4E; #100;
A = 8'h75; B = 8'h4F; #100;
A = 8'h75; B = 8'h50; #100;
A = 8'h75; B = 8'h51; #100;
A = 8'h75; B = 8'h52; #100;
A = 8'h75; B = 8'h53; #100;
A = 8'h75; B = 8'h54; #100;
A = 8'h75; B = 8'h55; #100;
A = 8'h75; B = 8'h56; #100;
A = 8'h75; B = 8'h57; #100;
A = 8'h75; B = 8'h58; #100;
A = 8'h75; B = 8'h59; #100;
A = 8'h75; B = 8'h5A; #100;
A = 8'h75; B = 8'h5B; #100;
A = 8'h75; B = 8'h5C; #100;
A = 8'h75; B = 8'h5D; #100;
A = 8'h75; B = 8'h5E; #100;
A = 8'h75; B = 8'h5F; #100;
A = 8'h75; B = 8'h60; #100;
A = 8'h75; B = 8'h61; #100;
A = 8'h75; B = 8'h62; #100;
A = 8'h75; B = 8'h63; #100;
A = 8'h75; B = 8'h64; #100;
A = 8'h75; B = 8'h65; #100;
A = 8'h75; B = 8'h66; #100;
A = 8'h75; B = 8'h67; #100;
A = 8'h75; B = 8'h68; #100;
A = 8'h75; B = 8'h69; #100;
A = 8'h75; B = 8'h6A; #100;
A = 8'h75; B = 8'h6B; #100;
A = 8'h75; B = 8'h6C; #100;
A = 8'h75; B = 8'h6D; #100;
A = 8'h75; B = 8'h6E; #100;
A = 8'h75; B = 8'h6F; #100;
A = 8'h75; B = 8'h70; #100;
A = 8'h75; B = 8'h71; #100;
A = 8'h75; B = 8'h72; #100;
A = 8'h75; B = 8'h73; #100;
A = 8'h75; B = 8'h74; #100;
A = 8'h75; B = 8'h75; #100;
A = 8'h75; B = 8'h76; #100;
A = 8'h75; B = 8'h77; #100;
A = 8'h75; B = 8'h78; #100;
A = 8'h75; B = 8'h79; #100;
A = 8'h75; B = 8'h7A; #100;
A = 8'h75; B = 8'h7B; #100;
A = 8'h75; B = 8'h7C; #100;
A = 8'h75; B = 8'h7D; #100;
A = 8'h75; B = 8'h7E; #100;
A = 8'h75; B = 8'h7F; #100;
A = 8'h75; B = 8'h80; #100;
A = 8'h75; B = 8'h81; #100;
A = 8'h75; B = 8'h82; #100;
A = 8'h75; B = 8'h83; #100;
A = 8'h75; B = 8'h84; #100;
A = 8'h75; B = 8'h85; #100;
A = 8'h75; B = 8'h86; #100;
A = 8'h75; B = 8'h87; #100;
A = 8'h75; B = 8'h88; #100;
A = 8'h75; B = 8'h89; #100;
A = 8'h75; B = 8'h8A; #100;
A = 8'h75; B = 8'h8B; #100;
A = 8'h75; B = 8'h8C; #100;
A = 8'h75; B = 8'h8D; #100;
A = 8'h75; B = 8'h8E; #100;
A = 8'h75; B = 8'h8F; #100;
A = 8'h75; B = 8'h90; #100;
A = 8'h75; B = 8'h91; #100;
A = 8'h75; B = 8'h92; #100;
A = 8'h75; B = 8'h93; #100;
A = 8'h75; B = 8'h94; #100;
A = 8'h75; B = 8'h95; #100;
A = 8'h75; B = 8'h96; #100;
A = 8'h75; B = 8'h97; #100;
A = 8'h75; B = 8'h98; #100;
A = 8'h75; B = 8'h99; #100;
A = 8'h75; B = 8'h9A; #100;
A = 8'h75; B = 8'h9B; #100;
A = 8'h75; B = 8'h9C; #100;
A = 8'h75; B = 8'h9D; #100;
A = 8'h75; B = 8'h9E; #100;
A = 8'h75; B = 8'h9F; #100;
A = 8'h75; B = 8'hA0; #100;
A = 8'h75; B = 8'hA1; #100;
A = 8'h75; B = 8'hA2; #100;
A = 8'h75; B = 8'hA3; #100;
A = 8'h75; B = 8'hA4; #100;
A = 8'h75; B = 8'hA5; #100;
A = 8'h75; B = 8'hA6; #100;
A = 8'h75; B = 8'hA7; #100;
A = 8'h75; B = 8'hA8; #100;
A = 8'h75; B = 8'hA9; #100;
A = 8'h75; B = 8'hAA; #100;
A = 8'h75; B = 8'hAB; #100;
A = 8'h75; B = 8'hAC; #100;
A = 8'h75; B = 8'hAD; #100;
A = 8'h75; B = 8'hAE; #100;
A = 8'h75; B = 8'hAF; #100;
A = 8'h75; B = 8'hB0; #100;
A = 8'h75; B = 8'hB1; #100;
A = 8'h75; B = 8'hB2; #100;
A = 8'h75; B = 8'hB3; #100;
A = 8'h75; B = 8'hB4; #100;
A = 8'h75; B = 8'hB5; #100;
A = 8'h75; B = 8'hB6; #100;
A = 8'h75; B = 8'hB7; #100;
A = 8'h75; B = 8'hB8; #100;
A = 8'h75; B = 8'hB9; #100;
A = 8'h75; B = 8'hBA; #100;
A = 8'h75; B = 8'hBB; #100;
A = 8'h75; B = 8'hBC; #100;
A = 8'h75; B = 8'hBD; #100;
A = 8'h75; B = 8'hBE; #100;
A = 8'h75; B = 8'hBF; #100;
A = 8'h75; B = 8'hC0; #100;
A = 8'h75; B = 8'hC1; #100;
A = 8'h75; B = 8'hC2; #100;
A = 8'h75; B = 8'hC3; #100;
A = 8'h75; B = 8'hC4; #100;
A = 8'h75; B = 8'hC5; #100;
A = 8'h75; B = 8'hC6; #100;
A = 8'h75; B = 8'hC7; #100;
A = 8'h75; B = 8'hC8; #100;
A = 8'h75; B = 8'hC9; #100;
A = 8'h75; B = 8'hCA; #100;
A = 8'h75; B = 8'hCB; #100;
A = 8'h75; B = 8'hCC; #100;
A = 8'h75; B = 8'hCD; #100;
A = 8'h75; B = 8'hCE; #100;
A = 8'h75; B = 8'hCF; #100;
A = 8'h75; B = 8'hD0; #100;
A = 8'h75; B = 8'hD1; #100;
A = 8'h75; B = 8'hD2; #100;
A = 8'h75; B = 8'hD3; #100;
A = 8'h75; B = 8'hD4; #100;
A = 8'h75; B = 8'hD5; #100;
A = 8'h75; B = 8'hD6; #100;
A = 8'h75; B = 8'hD7; #100;
A = 8'h75; B = 8'hD8; #100;
A = 8'h75; B = 8'hD9; #100;
A = 8'h75; B = 8'hDA; #100;
A = 8'h75; B = 8'hDB; #100;
A = 8'h75; B = 8'hDC; #100;
A = 8'h75; B = 8'hDD; #100;
A = 8'h75; B = 8'hDE; #100;
A = 8'h75; B = 8'hDF; #100;
A = 8'h75; B = 8'hE0; #100;
A = 8'h75; B = 8'hE1; #100;
A = 8'h75; B = 8'hE2; #100;
A = 8'h75; B = 8'hE3; #100;
A = 8'h75; B = 8'hE4; #100;
A = 8'h75; B = 8'hE5; #100;
A = 8'h75; B = 8'hE6; #100;
A = 8'h75; B = 8'hE7; #100;
A = 8'h75; B = 8'hE8; #100;
A = 8'h75; B = 8'hE9; #100;
A = 8'h75; B = 8'hEA; #100;
A = 8'h75; B = 8'hEB; #100;
A = 8'h75; B = 8'hEC; #100;
A = 8'h75; B = 8'hED; #100;
A = 8'h75; B = 8'hEE; #100;
A = 8'h75; B = 8'hEF; #100;
A = 8'h75; B = 8'hF0; #100;
A = 8'h75; B = 8'hF1; #100;
A = 8'h75; B = 8'hF2; #100;
A = 8'h75; B = 8'hF3; #100;
A = 8'h75; B = 8'hF4; #100;
A = 8'h75; B = 8'hF5; #100;
A = 8'h75; B = 8'hF6; #100;
A = 8'h75; B = 8'hF7; #100;
A = 8'h75; B = 8'hF8; #100;
A = 8'h75; B = 8'hF9; #100;
A = 8'h75; B = 8'hFA; #100;
A = 8'h75; B = 8'hFB; #100;
A = 8'h75; B = 8'hFC; #100;
A = 8'h75; B = 8'hFD; #100;
A = 8'h75; B = 8'hFE; #100;
A = 8'h75; B = 8'hFF; #100;
A = 8'h76; B = 8'h0; #100;
A = 8'h76; B = 8'h1; #100;
A = 8'h76; B = 8'h2; #100;
A = 8'h76; B = 8'h3; #100;
A = 8'h76; B = 8'h4; #100;
A = 8'h76; B = 8'h5; #100;
A = 8'h76; B = 8'h6; #100;
A = 8'h76; B = 8'h7; #100;
A = 8'h76; B = 8'h8; #100;
A = 8'h76; B = 8'h9; #100;
A = 8'h76; B = 8'hA; #100;
A = 8'h76; B = 8'hB; #100;
A = 8'h76; B = 8'hC; #100;
A = 8'h76; B = 8'hD; #100;
A = 8'h76; B = 8'hE; #100;
A = 8'h76; B = 8'hF; #100;
A = 8'h76; B = 8'h10; #100;
A = 8'h76; B = 8'h11; #100;
A = 8'h76; B = 8'h12; #100;
A = 8'h76; B = 8'h13; #100;
A = 8'h76; B = 8'h14; #100;
A = 8'h76; B = 8'h15; #100;
A = 8'h76; B = 8'h16; #100;
A = 8'h76; B = 8'h17; #100;
A = 8'h76; B = 8'h18; #100;
A = 8'h76; B = 8'h19; #100;
A = 8'h76; B = 8'h1A; #100;
A = 8'h76; B = 8'h1B; #100;
A = 8'h76; B = 8'h1C; #100;
A = 8'h76; B = 8'h1D; #100;
A = 8'h76; B = 8'h1E; #100;
A = 8'h76; B = 8'h1F; #100;
A = 8'h76; B = 8'h20; #100;
A = 8'h76; B = 8'h21; #100;
A = 8'h76; B = 8'h22; #100;
A = 8'h76; B = 8'h23; #100;
A = 8'h76; B = 8'h24; #100;
A = 8'h76; B = 8'h25; #100;
A = 8'h76; B = 8'h26; #100;
A = 8'h76; B = 8'h27; #100;
A = 8'h76; B = 8'h28; #100;
A = 8'h76; B = 8'h29; #100;
A = 8'h76; B = 8'h2A; #100;
A = 8'h76; B = 8'h2B; #100;
A = 8'h76; B = 8'h2C; #100;
A = 8'h76; B = 8'h2D; #100;
A = 8'h76; B = 8'h2E; #100;
A = 8'h76; B = 8'h2F; #100;
A = 8'h76; B = 8'h30; #100;
A = 8'h76; B = 8'h31; #100;
A = 8'h76; B = 8'h32; #100;
A = 8'h76; B = 8'h33; #100;
A = 8'h76; B = 8'h34; #100;
A = 8'h76; B = 8'h35; #100;
A = 8'h76; B = 8'h36; #100;
A = 8'h76; B = 8'h37; #100;
A = 8'h76; B = 8'h38; #100;
A = 8'h76; B = 8'h39; #100;
A = 8'h76; B = 8'h3A; #100;
A = 8'h76; B = 8'h3B; #100;
A = 8'h76; B = 8'h3C; #100;
A = 8'h76; B = 8'h3D; #100;
A = 8'h76; B = 8'h3E; #100;
A = 8'h76; B = 8'h3F; #100;
A = 8'h76; B = 8'h40; #100;
A = 8'h76; B = 8'h41; #100;
A = 8'h76; B = 8'h42; #100;
A = 8'h76; B = 8'h43; #100;
A = 8'h76; B = 8'h44; #100;
A = 8'h76; B = 8'h45; #100;
A = 8'h76; B = 8'h46; #100;
A = 8'h76; B = 8'h47; #100;
A = 8'h76; B = 8'h48; #100;
A = 8'h76; B = 8'h49; #100;
A = 8'h76; B = 8'h4A; #100;
A = 8'h76; B = 8'h4B; #100;
A = 8'h76; B = 8'h4C; #100;
A = 8'h76; B = 8'h4D; #100;
A = 8'h76; B = 8'h4E; #100;
A = 8'h76; B = 8'h4F; #100;
A = 8'h76; B = 8'h50; #100;
A = 8'h76; B = 8'h51; #100;
A = 8'h76; B = 8'h52; #100;
A = 8'h76; B = 8'h53; #100;
A = 8'h76; B = 8'h54; #100;
A = 8'h76; B = 8'h55; #100;
A = 8'h76; B = 8'h56; #100;
A = 8'h76; B = 8'h57; #100;
A = 8'h76; B = 8'h58; #100;
A = 8'h76; B = 8'h59; #100;
A = 8'h76; B = 8'h5A; #100;
A = 8'h76; B = 8'h5B; #100;
A = 8'h76; B = 8'h5C; #100;
A = 8'h76; B = 8'h5D; #100;
A = 8'h76; B = 8'h5E; #100;
A = 8'h76; B = 8'h5F; #100;
A = 8'h76; B = 8'h60; #100;
A = 8'h76; B = 8'h61; #100;
A = 8'h76; B = 8'h62; #100;
A = 8'h76; B = 8'h63; #100;
A = 8'h76; B = 8'h64; #100;
A = 8'h76; B = 8'h65; #100;
A = 8'h76; B = 8'h66; #100;
A = 8'h76; B = 8'h67; #100;
A = 8'h76; B = 8'h68; #100;
A = 8'h76; B = 8'h69; #100;
A = 8'h76; B = 8'h6A; #100;
A = 8'h76; B = 8'h6B; #100;
A = 8'h76; B = 8'h6C; #100;
A = 8'h76; B = 8'h6D; #100;
A = 8'h76; B = 8'h6E; #100;
A = 8'h76; B = 8'h6F; #100;
A = 8'h76; B = 8'h70; #100;
A = 8'h76; B = 8'h71; #100;
A = 8'h76; B = 8'h72; #100;
A = 8'h76; B = 8'h73; #100;
A = 8'h76; B = 8'h74; #100;
A = 8'h76; B = 8'h75; #100;
A = 8'h76; B = 8'h76; #100;
A = 8'h76; B = 8'h77; #100;
A = 8'h76; B = 8'h78; #100;
A = 8'h76; B = 8'h79; #100;
A = 8'h76; B = 8'h7A; #100;
A = 8'h76; B = 8'h7B; #100;
A = 8'h76; B = 8'h7C; #100;
A = 8'h76; B = 8'h7D; #100;
A = 8'h76; B = 8'h7E; #100;
A = 8'h76; B = 8'h7F; #100;
A = 8'h76; B = 8'h80; #100;
A = 8'h76; B = 8'h81; #100;
A = 8'h76; B = 8'h82; #100;
A = 8'h76; B = 8'h83; #100;
A = 8'h76; B = 8'h84; #100;
A = 8'h76; B = 8'h85; #100;
A = 8'h76; B = 8'h86; #100;
A = 8'h76; B = 8'h87; #100;
A = 8'h76; B = 8'h88; #100;
A = 8'h76; B = 8'h89; #100;
A = 8'h76; B = 8'h8A; #100;
A = 8'h76; B = 8'h8B; #100;
A = 8'h76; B = 8'h8C; #100;
A = 8'h76; B = 8'h8D; #100;
A = 8'h76; B = 8'h8E; #100;
A = 8'h76; B = 8'h8F; #100;
A = 8'h76; B = 8'h90; #100;
A = 8'h76; B = 8'h91; #100;
A = 8'h76; B = 8'h92; #100;
A = 8'h76; B = 8'h93; #100;
A = 8'h76; B = 8'h94; #100;
A = 8'h76; B = 8'h95; #100;
A = 8'h76; B = 8'h96; #100;
A = 8'h76; B = 8'h97; #100;
A = 8'h76; B = 8'h98; #100;
A = 8'h76; B = 8'h99; #100;
A = 8'h76; B = 8'h9A; #100;
A = 8'h76; B = 8'h9B; #100;
A = 8'h76; B = 8'h9C; #100;
A = 8'h76; B = 8'h9D; #100;
A = 8'h76; B = 8'h9E; #100;
A = 8'h76; B = 8'h9F; #100;
A = 8'h76; B = 8'hA0; #100;
A = 8'h76; B = 8'hA1; #100;
A = 8'h76; B = 8'hA2; #100;
A = 8'h76; B = 8'hA3; #100;
A = 8'h76; B = 8'hA4; #100;
A = 8'h76; B = 8'hA5; #100;
A = 8'h76; B = 8'hA6; #100;
A = 8'h76; B = 8'hA7; #100;
A = 8'h76; B = 8'hA8; #100;
A = 8'h76; B = 8'hA9; #100;
A = 8'h76; B = 8'hAA; #100;
A = 8'h76; B = 8'hAB; #100;
A = 8'h76; B = 8'hAC; #100;
A = 8'h76; B = 8'hAD; #100;
A = 8'h76; B = 8'hAE; #100;
A = 8'h76; B = 8'hAF; #100;
A = 8'h76; B = 8'hB0; #100;
A = 8'h76; B = 8'hB1; #100;
A = 8'h76; B = 8'hB2; #100;
A = 8'h76; B = 8'hB3; #100;
A = 8'h76; B = 8'hB4; #100;
A = 8'h76; B = 8'hB5; #100;
A = 8'h76; B = 8'hB6; #100;
A = 8'h76; B = 8'hB7; #100;
A = 8'h76; B = 8'hB8; #100;
A = 8'h76; B = 8'hB9; #100;
A = 8'h76; B = 8'hBA; #100;
A = 8'h76; B = 8'hBB; #100;
A = 8'h76; B = 8'hBC; #100;
A = 8'h76; B = 8'hBD; #100;
A = 8'h76; B = 8'hBE; #100;
A = 8'h76; B = 8'hBF; #100;
A = 8'h76; B = 8'hC0; #100;
A = 8'h76; B = 8'hC1; #100;
A = 8'h76; B = 8'hC2; #100;
A = 8'h76; B = 8'hC3; #100;
A = 8'h76; B = 8'hC4; #100;
A = 8'h76; B = 8'hC5; #100;
A = 8'h76; B = 8'hC6; #100;
A = 8'h76; B = 8'hC7; #100;
A = 8'h76; B = 8'hC8; #100;
A = 8'h76; B = 8'hC9; #100;
A = 8'h76; B = 8'hCA; #100;
A = 8'h76; B = 8'hCB; #100;
A = 8'h76; B = 8'hCC; #100;
A = 8'h76; B = 8'hCD; #100;
A = 8'h76; B = 8'hCE; #100;
A = 8'h76; B = 8'hCF; #100;
A = 8'h76; B = 8'hD0; #100;
A = 8'h76; B = 8'hD1; #100;
A = 8'h76; B = 8'hD2; #100;
A = 8'h76; B = 8'hD3; #100;
A = 8'h76; B = 8'hD4; #100;
A = 8'h76; B = 8'hD5; #100;
A = 8'h76; B = 8'hD6; #100;
A = 8'h76; B = 8'hD7; #100;
A = 8'h76; B = 8'hD8; #100;
A = 8'h76; B = 8'hD9; #100;
A = 8'h76; B = 8'hDA; #100;
A = 8'h76; B = 8'hDB; #100;
A = 8'h76; B = 8'hDC; #100;
A = 8'h76; B = 8'hDD; #100;
A = 8'h76; B = 8'hDE; #100;
A = 8'h76; B = 8'hDF; #100;
A = 8'h76; B = 8'hE0; #100;
A = 8'h76; B = 8'hE1; #100;
A = 8'h76; B = 8'hE2; #100;
A = 8'h76; B = 8'hE3; #100;
A = 8'h76; B = 8'hE4; #100;
A = 8'h76; B = 8'hE5; #100;
A = 8'h76; B = 8'hE6; #100;
A = 8'h76; B = 8'hE7; #100;
A = 8'h76; B = 8'hE8; #100;
A = 8'h76; B = 8'hE9; #100;
A = 8'h76; B = 8'hEA; #100;
A = 8'h76; B = 8'hEB; #100;
A = 8'h76; B = 8'hEC; #100;
A = 8'h76; B = 8'hED; #100;
A = 8'h76; B = 8'hEE; #100;
A = 8'h76; B = 8'hEF; #100;
A = 8'h76; B = 8'hF0; #100;
A = 8'h76; B = 8'hF1; #100;
A = 8'h76; B = 8'hF2; #100;
A = 8'h76; B = 8'hF3; #100;
A = 8'h76; B = 8'hF4; #100;
A = 8'h76; B = 8'hF5; #100;
A = 8'h76; B = 8'hF6; #100;
A = 8'h76; B = 8'hF7; #100;
A = 8'h76; B = 8'hF8; #100;
A = 8'h76; B = 8'hF9; #100;
A = 8'h76; B = 8'hFA; #100;
A = 8'h76; B = 8'hFB; #100;
A = 8'h76; B = 8'hFC; #100;
A = 8'h76; B = 8'hFD; #100;
A = 8'h76; B = 8'hFE; #100;
A = 8'h76; B = 8'hFF; #100;
A = 8'h77; B = 8'h0; #100;
A = 8'h77; B = 8'h1; #100;
A = 8'h77; B = 8'h2; #100;
A = 8'h77; B = 8'h3; #100;
A = 8'h77; B = 8'h4; #100;
A = 8'h77; B = 8'h5; #100;
A = 8'h77; B = 8'h6; #100;
A = 8'h77; B = 8'h7; #100;
A = 8'h77; B = 8'h8; #100;
A = 8'h77; B = 8'h9; #100;
A = 8'h77; B = 8'hA; #100;
A = 8'h77; B = 8'hB; #100;
A = 8'h77; B = 8'hC; #100;
A = 8'h77; B = 8'hD; #100;
A = 8'h77; B = 8'hE; #100;
A = 8'h77; B = 8'hF; #100;
A = 8'h77; B = 8'h10; #100;
A = 8'h77; B = 8'h11; #100;
A = 8'h77; B = 8'h12; #100;
A = 8'h77; B = 8'h13; #100;
A = 8'h77; B = 8'h14; #100;
A = 8'h77; B = 8'h15; #100;
A = 8'h77; B = 8'h16; #100;
A = 8'h77; B = 8'h17; #100;
A = 8'h77; B = 8'h18; #100;
A = 8'h77; B = 8'h19; #100;
A = 8'h77; B = 8'h1A; #100;
A = 8'h77; B = 8'h1B; #100;
A = 8'h77; B = 8'h1C; #100;
A = 8'h77; B = 8'h1D; #100;
A = 8'h77; B = 8'h1E; #100;
A = 8'h77; B = 8'h1F; #100;
A = 8'h77; B = 8'h20; #100;
A = 8'h77; B = 8'h21; #100;
A = 8'h77; B = 8'h22; #100;
A = 8'h77; B = 8'h23; #100;
A = 8'h77; B = 8'h24; #100;
A = 8'h77; B = 8'h25; #100;
A = 8'h77; B = 8'h26; #100;
A = 8'h77; B = 8'h27; #100;
A = 8'h77; B = 8'h28; #100;
A = 8'h77; B = 8'h29; #100;
A = 8'h77; B = 8'h2A; #100;
A = 8'h77; B = 8'h2B; #100;
A = 8'h77; B = 8'h2C; #100;
A = 8'h77; B = 8'h2D; #100;
A = 8'h77; B = 8'h2E; #100;
A = 8'h77; B = 8'h2F; #100;
A = 8'h77; B = 8'h30; #100;
A = 8'h77; B = 8'h31; #100;
A = 8'h77; B = 8'h32; #100;
A = 8'h77; B = 8'h33; #100;
A = 8'h77; B = 8'h34; #100;
A = 8'h77; B = 8'h35; #100;
A = 8'h77; B = 8'h36; #100;
A = 8'h77; B = 8'h37; #100;
A = 8'h77; B = 8'h38; #100;
A = 8'h77; B = 8'h39; #100;
A = 8'h77; B = 8'h3A; #100;
A = 8'h77; B = 8'h3B; #100;
A = 8'h77; B = 8'h3C; #100;
A = 8'h77; B = 8'h3D; #100;
A = 8'h77; B = 8'h3E; #100;
A = 8'h77; B = 8'h3F; #100;
A = 8'h77; B = 8'h40; #100;
A = 8'h77; B = 8'h41; #100;
A = 8'h77; B = 8'h42; #100;
A = 8'h77; B = 8'h43; #100;
A = 8'h77; B = 8'h44; #100;
A = 8'h77; B = 8'h45; #100;
A = 8'h77; B = 8'h46; #100;
A = 8'h77; B = 8'h47; #100;
A = 8'h77; B = 8'h48; #100;
A = 8'h77; B = 8'h49; #100;
A = 8'h77; B = 8'h4A; #100;
A = 8'h77; B = 8'h4B; #100;
A = 8'h77; B = 8'h4C; #100;
A = 8'h77; B = 8'h4D; #100;
A = 8'h77; B = 8'h4E; #100;
A = 8'h77; B = 8'h4F; #100;
A = 8'h77; B = 8'h50; #100;
A = 8'h77; B = 8'h51; #100;
A = 8'h77; B = 8'h52; #100;
A = 8'h77; B = 8'h53; #100;
A = 8'h77; B = 8'h54; #100;
A = 8'h77; B = 8'h55; #100;
A = 8'h77; B = 8'h56; #100;
A = 8'h77; B = 8'h57; #100;
A = 8'h77; B = 8'h58; #100;
A = 8'h77; B = 8'h59; #100;
A = 8'h77; B = 8'h5A; #100;
A = 8'h77; B = 8'h5B; #100;
A = 8'h77; B = 8'h5C; #100;
A = 8'h77; B = 8'h5D; #100;
A = 8'h77; B = 8'h5E; #100;
A = 8'h77; B = 8'h5F; #100;
A = 8'h77; B = 8'h60; #100;
A = 8'h77; B = 8'h61; #100;
A = 8'h77; B = 8'h62; #100;
A = 8'h77; B = 8'h63; #100;
A = 8'h77; B = 8'h64; #100;
A = 8'h77; B = 8'h65; #100;
A = 8'h77; B = 8'h66; #100;
A = 8'h77; B = 8'h67; #100;
A = 8'h77; B = 8'h68; #100;
A = 8'h77; B = 8'h69; #100;
A = 8'h77; B = 8'h6A; #100;
A = 8'h77; B = 8'h6B; #100;
A = 8'h77; B = 8'h6C; #100;
A = 8'h77; B = 8'h6D; #100;
A = 8'h77; B = 8'h6E; #100;
A = 8'h77; B = 8'h6F; #100;
A = 8'h77; B = 8'h70; #100;
A = 8'h77; B = 8'h71; #100;
A = 8'h77; B = 8'h72; #100;
A = 8'h77; B = 8'h73; #100;
A = 8'h77; B = 8'h74; #100;
A = 8'h77; B = 8'h75; #100;
A = 8'h77; B = 8'h76; #100;
A = 8'h77; B = 8'h77; #100;
A = 8'h77; B = 8'h78; #100;
A = 8'h77; B = 8'h79; #100;
A = 8'h77; B = 8'h7A; #100;
A = 8'h77; B = 8'h7B; #100;
A = 8'h77; B = 8'h7C; #100;
A = 8'h77; B = 8'h7D; #100;
A = 8'h77; B = 8'h7E; #100;
A = 8'h77; B = 8'h7F; #100;
A = 8'h77; B = 8'h80; #100;
A = 8'h77; B = 8'h81; #100;
A = 8'h77; B = 8'h82; #100;
A = 8'h77; B = 8'h83; #100;
A = 8'h77; B = 8'h84; #100;
A = 8'h77; B = 8'h85; #100;
A = 8'h77; B = 8'h86; #100;
A = 8'h77; B = 8'h87; #100;
A = 8'h77; B = 8'h88; #100;
A = 8'h77; B = 8'h89; #100;
A = 8'h77; B = 8'h8A; #100;
A = 8'h77; B = 8'h8B; #100;
A = 8'h77; B = 8'h8C; #100;
A = 8'h77; B = 8'h8D; #100;
A = 8'h77; B = 8'h8E; #100;
A = 8'h77; B = 8'h8F; #100;
A = 8'h77; B = 8'h90; #100;
A = 8'h77; B = 8'h91; #100;
A = 8'h77; B = 8'h92; #100;
A = 8'h77; B = 8'h93; #100;
A = 8'h77; B = 8'h94; #100;
A = 8'h77; B = 8'h95; #100;
A = 8'h77; B = 8'h96; #100;
A = 8'h77; B = 8'h97; #100;
A = 8'h77; B = 8'h98; #100;
A = 8'h77; B = 8'h99; #100;
A = 8'h77; B = 8'h9A; #100;
A = 8'h77; B = 8'h9B; #100;
A = 8'h77; B = 8'h9C; #100;
A = 8'h77; B = 8'h9D; #100;
A = 8'h77; B = 8'h9E; #100;
A = 8'h77; B = 8'h9F; #100;
A = 8'h77; B = 8'hA0; #100;
A = 8'h77; B = 8'hA1; #100;
A = 8'h77; B = 8'hA2; #100;
A = 8'h77; B = 8'hA3; #100;
A = 8'h77; B = 8'hA4; #100;
A = 8'h77; B = 8'hA5; #100;
A = 8'h77; B = 8'hA6; #100;
A = 8'h77; B = 8'hA7; #100;
A = 8'h77; B = 8'hA8; #100;
A = 8'h77; B = 8'hA9; #100;
A = 8'h77; B = 8'hAA; #100;
A = 8'h77; B = 8'hAB; #100;
A = 8'h77; B = 8'hAC; #100;
A = 8'h77; B = 8'hAD; #100;
A = 8'h77; B = 8'hAE; #100;
A = 8'h77; B = 8'hAF; #100;
A = 8'h77; B = 8'hB0; #100;
A = 8'h77; B = 8'hB1; #100;
A = 8'h77; B = 8'hB2; #100;
A = 8'h77; B = 8'hB3; #100;
A = 8'h77; B = 8'hB4; #100;
A = 8'h77; B = 8'hB5; #100;
A = 8'h77; B = 8'hB6; #100;
A = 8'h77; B = 8'hB7; #100;
A = 8'h77; B = 8'hB8; #100;
A = 8'h77; B = 8'hB9; #100;
A = 8'h77; B = 8'hBA; #100;
A = 8'h77; B = 8'hBB; #100;
A = 8'h77; B = 8'hBC; #100;
A = 8'h77; B = 8'hBD; #100;
A = 8'h77; B = 8'hBE; #100;
A = 8'h77; B = 8'hBF; #100;
A = 8'h77; B = 8'hC0; #100;
A = 8'h77; B = 8'hC1; #100;
A = 8'h77; B = 8'hC2; #100;
A = 8'h77; B = 8'hC3; #100;
A = 8'h77; B = 8'hC4; #100;
A = 8'h77; B = 8'hC5; #100;
A = 8'h77; B = 8'hC6; #100;
A = 8'h77; B = 8'hC7; #100;
A = 8'h77; B = 8'hC8; #100;
A = 8'h77; B = 8'hC9; #100;
A = 8'h77; B = 8'hCA; #100;
A = 8'h77; B = 8'hCB; #100;
A = 8'h77; B = 8'hCC; #100;
A = 8'h77; B = 8'hCD; #100;
A = 8'h77; B = 8'hCE; #100;
A = 8'h77; B = 8'hCF; #100;
A = 8'h77; B = 8'hD0; #100;
A = 8'h77; B = 8'hD1; #100;
A = 8'h77; B = 8'hD2; #100;
A = 8'h77; B = 8'hD3; #100;
A = 8'h77; B = 8'hD4; #100;
A = 8'h77; B = 8'hD5; #100;
A = 8'h77; B = 8'hD6; #100;
A = 8'h77; B = 8'hD7; #100;
A = 8'h77; B = 8'hD8; #100;
A = 8'h77; B = 8'hD9; #100;
A = 8'h77; B = 8'hDA; #100;
A = 8'h77; B = 8'hDB; #100;
A = 8'h77; B = 8'hDC; #100;
A = 8'h77; B = 8'hDD; #100;
A = 8'h77; B = 8'hDE; #100;
A = 8'h77; B = 8'hDF; #100;
A = 8'h77; B = 8'hE0; #100;
A = 8'h77; B = 8'hE1; #100;
A = 8'h77; B = 8'hE2; #100;
A = 8'h77; B = 8'hE3; #100;
A = 8'h77; B = 8'hE4; #100;
A = 8'h77; B = 8'hE5; #100;
A = 8'h77; B = 8'hE6; #100;
A = 8'h77; B = 8'hE7; #100;
A = 8'h77; B = 8'hE8; #100;
A = 8'h77; B = 8'hE9; #100;
A = 8'h77; B = 8'hEA; #100;
A = 8'h77; B = 8'hEB; #100;
A = 8'h77; B = 8'hEC; #100;
A = 8'h77; B = 8'hED; #100;
A = 8'h77; B = 8'hEE; #100;
A = 8'h77; B = 8'hEF; #100;
A = 8'h77; B = 8'hF0; #100;
A = 8'h77; B = 8'hF1; #100;
A = 8'h77; B = 8'hF2; #100;
A = 8'h77; B = 8'hF3; #100;
A = 8'h77; B = 8'hF4; #100;
A = 8'h77; B = 8'hF5; #100;
A = 8'h77; B = 8'hF6; #100;
A = 8'h77; B = 8'hF7; #100;
A = 8'h77; B = 8'hF8; #100;
A = 8'h77; B = 8'hF9; #100;
A = 8'h77; B = 8'hFA; #100;
A = 8'h77; B = 8'hFB; #100;
A = 8'h77; B = 8'hFC; #100;
A = 8'h77; B = 8'hFD; #100;
A = 8'h77; B = 8'hFE; #100;
A = 8'h77; B = 8'hFF; #100;
A = 8'h78; B = 8'h0; #100;
A = 8'h78; B = 8'h1; #100;
A = 8'h78; B = 8'h2; #100;
A = 8'h78; B = 8'h3; #100;
A = 8'h78; B = 8'h4; #100;
A = 8'h78; B = 8'h5; #100;
A = 8'h78; B = 8'h6; #100;
A = 8'h78; B = 8'h7; #100;
A = 8'h78; B = 8'h8; #100;
A = 8'h78; B = 8'h9; #100;
A = 8'h78; B = 8'hA; #100;
A = 8'h78; B = 8'hB; #100;
A = 8'h78; B = 8'hC; #100;
A = 8'h78; B = 8'hD; #100;
A = 8'h78; B = 8'hE; #100;
A = 8'h78; B = 8'hF; #100;
A = 8'h78; B = 8'h10; #100;
A = 8'h78; B = 8'h11; #100;
A = 8'h78; B = 8'h12; #100;
A = 8'h78; B = 8'h13; #100;
A = 8'h78; B = 8'h14; #100;
A = 8'h78; B = 8'h15; #100;
A = 8'h78; B = 8'h16; #100;
A = 8'h78; B = 8'h17; #100;
A = 8'h78; B = 8'h18; #100;
A = 8'h78; B = 8'h19; #100;
A = 8'h78; B = 8'h1A; #100;
A = 8'h78; B = 8'h1B; #100;
A = 8'h78; B = 8'h1C; #100;
A = 8'h78; B = 8'h1D; #100;
A = 8'h78; B = 8'h1E; #100;
A = 8'h78; B = 8'h1F; #100;
A = 8'h78; B = 8'h20; #100;
A = 8'h78; B = 8'h21; #100;
A = 8'h78; B = 8'h22; #100;
A = 8'h78; B = 8'h23; #100;
A = 8'h78; B = 8'h24; #100;
A = 8'h78; B = 8'h25; #100;
A = 8'h78; B = 8'h26; #100;
A = 8'h78; B = 8'h27; #100;
A = 8'h78; B = 8'h28; #100;
A = 8'h78; B = 8'h29; #100;
A = 8'h78; B = 8'h2A; #100;
A = 8'h78; B = 8'h2B; #100;
A = 8'h78; B = 8'h2C; #100;
A = 8'h78; B = 8'h2D; #100;
A = 8'h78; B = 8'h2E; #100;
A = 8'h78; B = 8'h2F; #100;
A = 8'h78; B = 8'h30; #100;
A = 8'h78; B = 8'h31; #100;
A = 8'h78; B = 8'h32; #100;
A = 8'h78; B = 8'h33; #100;
A = 8'h78; B = 8'h34; #100;
A = 8'h78; B = 8'h35; #100;
A = 8'h78; B = 8'h36; #100;
A = 8'h78; B = 8'h37; #100;
A = 8'h78; B = 8'h38; #100;
A = 8'h78; B = 8'h39; #100;
A = 8'h78; B = 8'h3A; #100;
A = 8'h78; B = 8'h3B; #100;
A = 8'h78; B = 8'h3C; #100;
A = 8'h78; B = 8'h3D; #100;
A = 8'h78; B = 8'h3E; #100;
A = 8'h78; B = 8'h3F; #100;
A = 8'h78; B = 8'h40; #100;
A = 8'h78; B = 8'h41; #100;
A = 8'h78; B = 8'h42; #100;
A = 8'h78; B = 8'h43; #100;
A = 8'h78; B = 8'h44; #100;
A = 8'h78; B = 8'h45; #100;
A = 8'h78; B = 8'h46; #100;
A = 8'h78; B = 8'h47; #100;
A = 8'h78; B = 8'h48; #100;
A = 8'h78; B = 8'h49; #100;
A = 8'h78; B = 8'h4A; #100;
A = 8'h78; B = 8'h4B; #100;
A = 8'h78; B = 8'h4C; #100;
A = 8'h78; B = 8'h4D; #100;
A = 8'h78; B = 8'h4E; #100;
A = 8'h78; B = 8'h4F; #100;
A = 8'h78; B = 8'h50; #100;
A = 8'h78; B = 8'h51; #100;
A = 8'h78; B = 8'h52; #100;
A = 8'h78; B = 8'h53; #100;
A = 8'h78; B = 8'h54; #100;
A = 8'h78; B = 8'h55; #100;
A = 8'h78; B = 8'h56; #100;
A = 8'h78; B = 8'h57; #100;
A = 8'h78; B = 8'h58; #100;
A = 8'h78; B = 8'h59; #100;
A = 8'h78; B = 8'h5A; #100;
A = 8'h78; B = 8'h5B; #100;
A = 8'h78; B = 8'h5C; #100;
A = 8'h78; B = 8'h5D; #100;
A = 8'h78; B = 8'h5E; #100;
A = 8'h78; B = 8'h5F; #100;
A = 8'h78; B = 8'h60; #100;
A = 8'h78; B = 8'h61; #100;
A = 8'h78; B = 8'h62; #100;
A = 8'h78; B = 8'h63; #100;
A = 8'h78; B = 8'h64; #100;
A = 8'h78; B = 8'h65; #100;
A = 8'h78; B = 8'h66; #100;
A = 8'h78; B = 8'h67; #100;
A = 8'h78; B = 8'h68; #100;
A = 8'h78; B = 8'h69; #100;
A = 8'h78; B = 8'h6A; #100;
A = 8'h78; B = 8'h6B; #100;
A = 8'h78; B = 8'h6C; #100;
A = 8'h78; B = 8'h6D; #100;
A = 8'h78; B = 8'h6E; #100;
A = 8'h78; B = 8'h6F; #100;
A = 8'h78; B = 8'h70; #100;
A = 8'h78; B = 8'h71; #100;
A = 8'h78; B = 8'h72; #100;
A = 8'h78; B = 8'h73; #100;
A = 8'h78; B = 8'h74; #100;
A = 8'h78; B = 8'h75; #100;
A = 8'h78; B = 8'h76; #100;
A = 8'h78; B = 8'h77; #100;
A = 8'h78; B = 8'h78; #100;
A = 8'h78; B = 8'h79; #100;
A = 8'h78; B = 8'h7A; #100;
A = 8'h78; B = 8'h7B; #100;
A = 8'h78; B = 8'h7C; #100;
A = 8'h78; B = 8'h7D; #100;
A = 8'h78; B = 8'h7E; #100;
A = 8'h78; B = 8'h7F; #100;
A = 8'h78; B = 8'h80; #100;
A = 8'h78; B = 8'h81; #100;
A = 8'h78; B = 8'h82; #100;
A = 8'h78; B = 8'h83; #100;
A = 8'h78; B = 8'h84; #100;
A = 8'h78; B = 8'h85; #100;
A = 8'h78; B = 8'h86; #100;
A = 8'h78; B = 8'h87; #100;
A = 8'h78; B = 8'h88; #100;
A = 8'h78; B = 8'h89; #100;
A = 8'h78; B = 8'h8A; #100;
A = 8'h78; B = 8'h8B; #100;
A = 8'h78; B = 8'h8C; #100;
A = 8'h78; B = 8'h8D; #100;
A = 8'h78; B = 8'h8E; #100;
A = 8'h78; B = 8'h8F; #100;
A = 8'h78; B = 8'h90; #100;
A = 8'h78; B = 8'h91; #100;
A = 8'h78; B = 8'h92; #100;
A = 8'h78; B = 8'h93; #100;
A = 8'h78; B = 8'h94; #100;
A = 8'h78; B = 8'h95; #100;
A = 8'h78; B = 8'h96; #100;
A = 8'h78; B = 8'h97; #100;
A = 8'h78; B = 8'h98; #100;
A = 8'h78; B = 8'h99; #100;
A = 8'h78; B = 8'h9A; #100;
A = 8'h78; B = 8'h9B; #100;
A = 8'h78; B = 8'h9C; #100;
A = 8'h78; B = 8'h9D; #100;
A = 8'h78; B = 8'h9E; #100;
A = 8'h78; B = 8'h9F; #100;
A = 8'h78; B = 8'hA0; #100;
A = 8'h78; B = 8'hA1; #100;
A = 8'h78; B = 8'hA2; #100;
A = 8'h78; B = 8'hA3; #100;
A = 8'h78; B = 8'hA4; #100;
A = 8'h78; B = 8'hA5; #100;
A = 8'h78; B = 8'hA6; #100;
A = 8'h78; B = 8'hA7; #100;
A = 8'h78; B = 8'hA8; #100;
A = 8'h78; B = 8'hA9; #100;
A = 8'h78; B = 8'hAA; #100;
A = 8'h78; B = 8'hAB; #100;
A = 8'h78; B = 8'hAC; #100;
A = 8'h78; B = 8'hAD; #100;
A = 8'h78; B = 8'hAE; #100;
A = 8'h78; B = 8'hAF; #100;
A = 8'h78; B = 8'hB0; #100;
A = 8'h78; B = 8'hB1; #100;
A = 8'h78; B = 8'hB2; #100;
A = 8'h78; B = 8'hB3; #100;
A = 8'h78; B = 8'hB4; #100;
A = 8'h78; B = 8'hB5; #100;
A = 8'h78; B = 8'hB6; #100;
A = 8'h78; B = 8'hB7; #100;
A = 8'h78; B = 8'hB8; #100;
A = 8'h78; B = 8'hB9; #100;
A = 8'h78; B = 8'hBA; #100;
A = 8'h78; B = 8'hBB; #100;
A = 8'h78; B = 8'hBC; #100;
A = 8'h78; B = 8'hBD; #100;
A = 8'h78; B = 8'hBE; #100;
A = 8'h78; B = 8'hBF; #100;
A = 8'h78; B = 8'hC0; #100;
A = 8'h78; B = 8'hC1; #100;
A = 8'h78; B = 8'hC2; #100;
A = 8'h78; B = 8'hC3; #100;
A = 8'h78; B = 8'hC4; #100;
A = 8'h78; B = 8'hC5; #100;
A = 8'h78; B = 8'hC6; #100;
A = 8'h78; B = 8'hC7; #100;
A = 8'h78; B = 8'hC8; #100;
A = 8'h78; B = 8'hC9; #100;
A = 8'h78; B = 8'hCA; #100;
A = 8'h78; B = 8'hCB; #100;
A = 8'h78; B = 8'hCC; #100;
A = 8'h78; B = 8'hCD; #100;
A = 8'h78; B = 8'hCE; #100;
A = 8'h78; B = 8'hCF; #100;
A = 8'h78; B = 8'hD0; #100;
A = 8'h78; B = 8'hD1; #100;
A = 8'h78; B = 8'hD2; #100;
A = 8'h78; B = 8'hD3; #100;
A = 8'h78; B = 8'hD4; #100;
A = 8'h78; B = 8'hD5; #100;
A = 8'h78; B = 8'hD6; #100;
A = 8'h78; B = 8'hD7; #100;
A = 8'h78; B = 8'hD8; #100;
A = 8'h78; B = 8'hD9; #100;
A = 8'h78; B = 8'hDA; #100;
A = 8'h78; B = 8'hDB; #100;
A = 8'h78; B = 8'hDC; #100;
A = 8'h78; B = 8'hDD; #100;
A = 8'h78; B = 8'hDE; #100;
A = 8'h78; B = 8'hDF; #100;
A = 8'h78; B = 8'hE0; #100;
A = 8'h78; B = 8'hE1; #100;
A = 8'h78; B = 8'hE2; #100;
A = 8'h78; B = 8'hE3; #100;
A = 8'h78; B = 8'hE4; #100;
A = 8'h78; B = 8'hE5; #100;
A = 8'h78; B = 8'hE6; #100;
A = 8'h78; B = 8'hE7; #100;
A = 8'h78; B = 8'hE8; #100;
A = 8'h78; B = 8'hE9; #100;
A = 8'h78; B = 8'hEA; #100;
A = 8'h78; B = 8'hEB; #100;
A = 8'h78; B = 8'hEC; #100;
A = 8'h78; B = 8'hED; #100;
A = 8'h78; B = 8'hEE; #100;
A = 8'h78; B = 8'hEF; #100;
A = 8'h78; B = 8'hF0; #100;
A = 8'h78; B = 8'hF1; #100;
A = 8'h78; B = 8'hF2; #100;
A = 8'h78; B = 8'hF3; #100;
A = 8'h78; B = 8'hF4; #100;
A = 8'h78; B = 8'hF5; #100;
A = 8'h78; B = 8'hF6; #100;
A = 8'h78; B = 8'hF7; #100;
A = 8'h78; B = 8'hF8; #100;
A = 8'h78; B = 8'hF9; #100;
A = 8'h78; B = 8'hFA; #100;
A = 8'h78; B = 8'hFB; #100;
A = 8'h78; B = 8'hFC; #100;
A = 8'h78; B = 8'hFD; #100;
A = 8'h78; B = 8'hFE; #100;
A = 8'h78; B = 8'hFF; #100;
A = 8'h79; B = 8'h0; #100;
A = 8'h79; B = 8'h1; #100;
A = 8'h79; B = 8'h2; #100;
A = 8'h79; B = 8'h3; #100;
A = 8'h79; B = 8'h4; #100;
A = 8'h79; B = 8'h5; #100;
A = 8'h79; B = 8'h6; #100;
A = 8'h79; B = 8'h7; #100;
A = 8'h79; B = 8'h8; #100;
A = 8'h79; B = 8'h9; #100;
A = 8'h79; B = 8'hA; #100;
A = 8'h79; B = 8'hB; #100;
A = 8'h79; B = 8'hC; #100;
A = 8'h79; B = 8'hD; #100;
A = 8'h79; B = 8'hE; #100;
A = 8'h79; B = 8'hF; #100;
A = 8'h79; B = 8'h10; #100;
A = 8'h79; B = 8'h11; #100;
A = 8'h79; B = 8'h12; #100;
A = 8'h79; B = 8'h13; #100;
A = 8'h79; B = 8'h14; #100;
A = 8'h79; B = 8'h15; #100;
A = 8'h79; B = 8'h16; #100;
A = 8'h79; B = 8'h17; #100;
A = 8'h79; B = 8'h18; #100;
A = 8'h79; B = 8'h19; #100;
A = 8'h79; B = 8'h1A; #100;
A = 8'h79; B = 8'h1B; #100;
A = 8'h79; B = 8'h1C; #100;
A = 8'h79; B = 8'h1D; #100;
A = 8'h79; B = 8'h1E; #100;
A = 8'h79; B = 8'h1F; #100;
A = 8'h79; B = 8'h20; #100;
A = 8'h79; B = 8'h21; #100;
A = 8'h79; B = 8'h22; #100;
A = 8'h79; B = 8'h23; #100;
A = 8'h79; B = 8'h24; #100;
A = 8'h79; B = 8'h25; #100;
A = 8'h79; B = 8'h26; #100;
A = 8'h79; B = 8'h27; #100;
A = 8'h79; B = 8'h28; #100;
A = 8'h79; B = 8'h29; #100;
A = 8'h79; B = 8'h2A; #100;
A = 8'h79; B = 8'h2B; #100;
A = 8'h79; B = 8'h2C; #100;
A = 8'h79; B = 8'h2D; #100;
A = 8'h79; B = 8'h2E; #100;
A = 8'h79; B = 8'h2F; #100;
A = 8'h79; B = 8'h30; #100;
A = 8'h79; B = 8'h31; #100;
A = 8'h79; B = 8'h32; #100;
A = 8'h79; B = 8'h33; #100;
A = 8'h79; B = 8'h34; #100;
A = 8'h79; B = 8'h35; #100;
A = 8'h79; B = 8'h36; #100;
A = 8'h79; B = 8'h37; #100;
A = 8'h79; B = 8'h38; #100;
A = 8'h79; B = 8'h39; #100;
A = 8'h79; B = 8'h3A; #100;
A = 8'h79; B = 8'h3B; #100;
A = 8'h79; B = 8'h3C; #100;
A = 8'h79; B = 8'h3D; #100;
A = 8'h79; B = 8'h3E; #100;
A = 8'h79; B = 8'h3F; #100;
A = 8'h79; B = 8'h40; #100;
A = 8'h79; B = 8'h41; #100;
A = 8'h79; B = 8'h42; #100;
A = 8'h79; B = 8'h43; #100;
A = 8'h79; B = 8'h44; #100;
A = 8'h79; B = 8'h45; #100;
A = 8'h79; B = 8'h46; #100;
A = 8'h79; B = 8'h47; #100;
A = 8'h79; B = 8'h48; #100;
A = 8'h79; B = 8'h49; #100;
A = 8'h79; B = 8'h4A; #100;
A = 8'h79; B = 8'h4B; #100;
A = 8'h79; B = 8'h4C; #100;
A = 8'h79; B = 8'h4D; #100;
A = 8'h79; B = 8'h4E; #100;
A = 8'h79; B = 8'h4F; #100;
A = 8'h79; B = 8'h50; #100;
A = 8'h79; B = 8'h51; #100;
A = 8'h79; B = 8'h52; #100;
A = 8'h79; B = 8'h53; #100;
A = 8'h79; B = 8'h54; #100;
A = 8'h79; B = 8'h55; #100;
A = 8'h79; B = 8'h56; #100;
A = 8'h79; B = 8'h57; #100;
A = 8'h79; B = 8'h58; #100;
A = 8'h79; B = 8'h59; #100;
A = 8'h79; B = 8'h5A; #100;
A = 8'h79; B = 8'h5B; #100;
A = 8'h79; B = 8'h5C; #100;
A = 8'h79; B = 8'h5D; #100;
A = 8'h79; B = 8'h5E; #100;
A = 8'h79; B = 8'h5F; #100;
A = 8'h79; B = 8'h60; #100;
A = 8'h79; B = 8'h61; #100;
A = 8'h79; B = 8'h62; #100;
A = 8'h79; B = 8'h63; #100;
A = 8'h79; B = 8'h64; #100;
A = 8'h79; B = 8'h65; #100;
A = 8'h79; B = 8'h66; #100;
A = 8'h79; B = 8'h67; #100;
A = 8'h79; B = 8'h68; #100;
A = 8'h79; B = 8'h69; #100;
A = 8'h79; B = 8'h6A; #100;
A = 8'h79; B = 8'h6B; #100;
A = 8'h79; B = 8'h6C; #100;
A = 8'h79; B = 8'h6D; #100;
A = 8'h79; B = 8'h6E; #100;
A = 8'h79; B = 8'h6F; #100;
A = 8'h79; B = 8'h70; #100;
A = 8'h79; B = 8'h71; #100;
A = 8'h79; B = 8'h72; #100;
A = 8'h79; B = 8'h73; #100;
A = 8'h79; B = 8'h74; #100;
A = 8'h79; B = 8'h75; #100;
A = 8'h79; B = 8'h76; #100;
A = 8'h79; B = 8'h77; #100;
A = 8'h79; B = 8'h78; #100;
A = 8'h79; B = 8'h79; #100;
A = 8'h79; B = 8'h7A; #100;
A = 8'h79; B = 8'h7B; #100;
A = 8'h79; B = 8'h7C; #100;
A = 8'h79; B = 8'h7D; #100;
A = 8'h79; B = 8'h7E; #100;
A = 8'h79; B = 8'h7F; #100;
A = 8'h79; B = 8'h80; #100;
A = 8'h79; B = 8'h81; #100;
A = 8'h79; B = 8'h82; #100;
A = 8'h79; B = 8'h83; #100;
A = 8'h79; B = 8'h84; #100;
A = 8'h79; B = 8'h85; #100;
A = 8'h79; B = 8'h86; #100;
A = 8'h79; B = 8'h87; #100;
A = 8'h79; B = 8'h88; #100;
A = 8'h79; B = 8'h89; #100;
A = 8'h79; B = 8'h8A; #100;
A = 8'h79; B = 8'h8B; #100;
A = 8'h79; B = 8'h8C; #100;
A = 8'h79; B = 8'h8D; #100;
A = 8'h79; B = 8'h8E; #100;
A = 8'h79; B = 8'h8F; #100;
A = 8'h79; B = 8'h90; #100;
A = 8'h79; B = 8'h91; #100;
A = 8'h79; B = 8'h92; #100;
A = 8'h79; B = 8'h93; #100;
A = 8'h79; B = 8'h94; #100;
A = 8'h79; B = 8'h95; #100;
A = 8'h79; B = 8'h96; #100;
A = 8'h79; B = 8'h97; #100;
A = 8'h79; B = 8'h98; #100;
A = 8'h79; B = 8'h99; #100;
A = 8'h79; B = 8'h9A; #100;
A = 8'h79; B = 8'h9B; #100;
A = 8'h79; B = 8'h9C; #100;
A = 8'h79; B = 8'h9D; #100;
A = 8'h79; B = 8'h9E; #100;
A = 8'h79; B = 8'h9F; #100;
A = 8'h79; B = 8'hA0; #100;
A = 8'h79; B = 8'hA1; #100;
A = 8'h79; B = 8'hA2; #100;
A = 8'h79; B = 8'hA3; #100;
A = 8'h79; B = 8'hA4; #100;
A = 8'h79; B = 8'hA5; #100;
A = 8'h79; B = 8'hA6; #100;
A = 8'h79; B = 8'hA7; #100;
A = 8'h79; B = 8'hA8; #100;
A = 8'h79; B = 8'hA9; #100;
A = 8'h79; B = 8'hAA; #100;
A = 8'h79; B = 8'hAB; #100;
A = 8'h79; B = 8'hAC; #100;
A = 8'h79; B = 8'hAD; #100;
A = 8'h79; B = 8'hAE; #100;
A = 8'h79; B = 8'hAF; #100;
A = 8'h79; B = 8'hB0; #100;
A = 8'h79; B = 8'hB1; #100;
A = 8'h79; B = 8'hB2; #100;
A = 8'h79; B = 8'hB3; #100;
A = 8'h79; B = 8'hB4; #100;
A = 8'h79; B = 8'hB5; #100;
A = 8'h79; B = 8'hB6; #100;
A = 8'h79; B = 8'hB7; #100;
A = 8'h79; B = 8'hB8; #100;
A = 8'h79; B = 8'hB9; #100;
A = 8'h79; B = 8'hBA; #100;
A = 8'h79; B = 8'hBB; #100;
A = 8'h79; B = 8'hBC; #100;
A = 8'h79; B = 8'hBD; #100;
A = 8'h79; B = 8'hBE; #100;
A = 8'h79; B = 8'hBF; #100;
A = 8'h79; B = 8'hC0; #100;
A = 8'h79; B = 8'hC1; #100;
A = 8'h79; B = 8'hC2; #100;
A = 8'h79; B = 8'hC3; #100;
A = 8'h79; B = 8'hC4; #100;
A = 8'h79; B = 8'hC5; #100;
A = 8'h79; B = 8'hC6; #100;
A = 8'h79; B = 8'hC7; #100;
A = 8'h79; B = 8'hC8; #100;
A = 8'h79; B = 8'hC9; #100;
A = 8'h79; B = 8'hCA; #100;
A = 8'h79; B = 8'hCB; #100;
A = 8'h79; B = 8'hCC; #100;
A = 8'h79; B = 8'hCD; #100;
A = 8'h79; B = 8'hCE; #100;
A = 8'h79; B = 8'hCF; #100;
A = 8'h79; B = 8'hD0; #100;
A = 8'h79; B = 8'hD1; #100;
A = 8'h79; B = 8'hD2; #100;
A = 8'h79; B = 8'hD3; #100;
A = 8'h79; B = 8'hD4; #100;
A = 8'h79; B = 8'hD5; #100;
A = 8'h79; B = 8'hD6; #100;
A = 8'h79; B = 8'hD7; #100;
A = 8'h79; B = 8'hD8; #100;
A = 8'h79; B = 8'hD9; #100;
A = 8'h79; B = 8'hDA; #100;
A = 8'h79; B = 8'hDB; #100;
A = 8'h79; B = 8'hDC; #100;
A = 8'h79; B = 8'hDD; #100;
A = 8'h79; B = 8'hDE; #100;
A = 8'h79; B = 8'hDF; #100;
A = 8'h79; B = 8'hE0; #100;
A = 8'h79; B = 8'hE1; #100;
A = 8'h79; B = 8'hE2; #100;
A = 8'h79; B = 8'hE3; #100;
A = 8'h79; B = 8'hE4; #100;
A = 8'h79; B = 8'hE5; #100;
A = 8'h79; B = 8'hE6; #100;
A = 8'h79; B = 8'hE7; #100;
A = 8'h79; B = 8'hE8; #100;
A = 8'h79; B = 8'hE9; #100;
A = 8'h79; B = 8'hEA; #100;
A = 8'h79; B = 8'hEB; #100;
A = 8'h79; B = 8'hEC; #100;
A = 8'h79; B = 8'hED; #100;
A = 8'h79; B = 8'hEE; #100;
A = 8'h79; B = 8'hEF; #100;
A = 8'h79; B = 8'hF0; #100;
A = 8'h79; B = 8'hF1; #100;
A = 8'h79; B = 8'hF2; #100;
A = 8'h79; B = 8'hF3; #100;
A = 8'h79; B = 8'hF4; #100;
A = 8'h79; B = 8'hF5; #100;
A = 8'h79; B = 8'hF6; #100;
A = 8'h79; B = 8'hF7; #100;
A = 8'h79; B = 8'hF8; #100;
A = 8'h79; B = 8'hF9; #100;
A = 8'h79; B = 8'hFA; #100;
A = 8'h79; B = 8'hFB; #100;
A = 8'h79; B = 8'hFC; #100;
A = 8'h79; B = 8'hFD; #100;
A = 8'h79; B = 8'hFE; #100;
A = 8'h79; B = 8'hFF; #100;
A = 8'h7A; B = 8'h0; #100;
A = 8'h7A; B = 8'h1; #100;
A = 8'h7A; B = 8'h2; #100;
A = 8'h7A; B = 8'h3; #100;
A = 8'h7A; B = 8'h4; #100;
A = 8'h7A; B = 8'h5; #100;
A = 8'h7A; B = 8'h6; #100;
A = 8'h7A; B = 8'h7; #100;
A = 8'h7A; B = 8'h8; #100;
A = 8'h7A; B = 8'h9; #100;
A = 8'h7A; B = 8'hA; #100;
A = 8'h7A; B = 8'hB; #100;
A = 8'h7A; B = 8'hC; #100;
A = 8'h7A; B = 8'hD; #100;
A = 8'h7A; B = 8'hE; #100;
A = 8'h7A; B = 8'hF; #100;
A = 8'h7A; B = 8'h10; #100;
A = 8'h7A; B = 8'h11; #100;
A = 8'h7A; B = 8'h12; #100;
A = 8'h7A; B = 8'h13; #100;
A = 8'h7A; B = 8'h14; #100;
A = 8'h7A; B = 8'h15; #100;
A = 8'h7A; B = 8'h16; #100;
A = 8'h7A; B = 8'h17; #100;
A = 8'h7A; B = 8'h18; #100;
A = 8'h7A; B = 8'h19; #100;
A = 8'h7A; B = 8'h1A; #100;
A = 8'h7A; B = 8'h1B; #100;
A = 8'h7A; B = 8'h1C; #100;
A = 8'h7A; B = 8'h1D; #100;
A = 8'h7A; B = 8'h1E; #100;
A = 8'h7A; B = 8'h1F; #100;
A = 8'h7A; B = 8'h20; #100;
A = 8'h7A; B = 8'h21; #100;
A = 8'h7A; B = 8'h22; #100;
A = 8'h7A; B = 8'h23; #100;
A = 8'h7A; B = 8'h24; #100;
A = 8'h7A; B = 8'h25; #100;
A = 8'h7A; B = 8'h26; #100;
A = 8'h7A; B = 8'h27; #100;
A = 8'h7A; B = 8'h28; #100;
A = 8'h7A; B = 8'h29; #100;
A = 8'h7A; B = 8'h2A; #100;
A = 8'h7A; B = 8'h2B; #100;
A = 8'h7A; B = 8'h2C; #100;
A = 8'h7A; B = 8'h2D; #100;
A = 8'h7A; B = 8'h2E; #100;
A = 8'h7A; B = 8'h2F; #100;
A = 8'h7A; B = 8'h30; #100;
A = 8'h7A; B = 8'h31; #100;
A = 8'h7A; B = 8'h32; #100;
A = 8'h7A; B = 8'h33; #100;
A = 8'h7A; B = 8'h34; #100;
A = 8'h7A; B = 8'h35; #100;
A = 8'h7A; B = 8'h36; #100;
A = 8'h7A; B = 8'h37; #100;
A = 8'h7A; B = 8'h38; #100;
A = 8'h7A; B = 8'h39; #100;
A = 8'h7A; B = 8'h3A; #100;
A = 8'h7A; B = 8'h3B; #100;
A = 8'h7A; B = 8'h3C; #100;
A = 8'h7A; B = 8'h3D; #100;
A = 8'h7A; B = 8'h3E; #100;
A = 8'h7A; B = 8'h3F; #100;
A = 8'h7A; B = 8'h40; #100;
A = 8'h7A; B = 8'h41; #100;
A = 8'h7A; B = 8'h42; #100;
A = 8'h7A; B = 8'h43; #100;
A = 8'h7A; B = 8'h44; #100;
A = 8'h7A; B = 8'h45; #100;
A = 8'h7A; B = 8'h46; #100;
A = 8'h7A; B = 8'h47; #100;
A = 8'h7A; B = 8'h48; #100;
A = 8'h7A; B = 8'h49; #100;
A = 8'h7A; B = 8'h4A; #100;
A = 8'h7A; B = 8'h4B; #100;
A = 8'h7A; B = 8'h4C; #100;
A = 8'h7A; B = 8'h4D; #100;
A = 8'h7A; B = 8'h4E; #100;
A = 8'h7A; B = 8'h4F; #100;
A = 8'h7A; B = 8'h50; #100;
A = 8'h7A; B = 8'h51; #100;
A = 8'h7A; B = 8'h52; #100;
A = 8'h7A; B = 8'h53; #100;
A = 8'h7A; B = 8'h54; #100;
A = 8'h7A; B = 8'h55; #100;
A = 8'h7A; B = 8'h56; #100;
A = 8'h7A; B = 8'h57; #100;
A = 8'h7A; B = 8'h58; #100;
A = 8'h7A; B = 8'h59; #100;
A = 8'h7A; B = 8'h5A; #100;
A = 8'h7A; B = 8'h5B; #100;
A = 8'h7A; B = 8'h5C; #100;
A = 8'h7A; B = 8'h5D; #100;
A = 8'h7A; B = 8'h5E; #100;
A = 8'h7A; B = 8'h5F; #100;
A = 8'h7A; B = 8'h60; #100;
A = 8'h7A; B = 8'h61; #100;
A = 8'h7A; B = 8'h62; #100;
A = 8'h7A; B = 8'h63; #100;
A = 8'h7A; B = 8'h64; #100;
A = 8'h7A; B = 8'h65; #100;
A = 8'h7A; B = 8'h66; #100;
A = 8'h7A; B = 8'h67; #100;
A = 8'h7A; B = 8'h68; #100;
A = 8'h7A; B = 8'h69; #100;
A = 8'h7A; B = 8'h6A; #100;
A = 8'h7A; B = 8'h6B; #100;
A = 8'h7A; B = 8'h6C; #100;
A = 8'h7A; B = 8'h6D; #100;
A = 8'h7A; B = 8'h6E; #100;
A = 8'h7A; B = 8'h6F; #100;
A = 8'h7A; B = 8'h70; #100;
A = 8'h7A; B = 8'h71; #100;
A = 8'h7A; B = 8'h72; #100;
A = 8'h7A; B = 8'h73; #100;
A = 8'h7A; B = 8'h74; #100;
A = 8'h7A; B = 8'h75; #100;
A = 8'h7A; B = 8'h76; #100;
A = 8'h7A; B = 8'h77; #100;
A = 8'h7A; B = 8'h78; #100;
A = 8'h7A; B = 8'h79; #100;
A = 8'h7A; B = 8'h7A; #100;
A = 8'h7A; B = 8'h7B; #100;
A = 8'h7A; B = 8'h7C; #100;
A = 8'h7A; B = 8'h7D; #100;
A = 8'h7A; B = 8'h7E; #100;
A = 8'h7A; B = 8'h7F; #100;
A = 8'h7A; B = 8'h80; #100;
A = 8'h7A; B = 8'h81; #100;
A = 8'h7A; B = 8'h82; #100;
A = 8'h7A; B = 8'h83; #100;
A = 8'h7A; B = 8'h84; #100;
A = 8'h7A; B = 8'h85; #100;
A = 8'h7A; B = 8'h86; #100;
A = 8'h7A; B = 8'h87; #100;
A = 8'h7A; B = 8'h88; #100;
A = 8'h7A; B = 8'h89; #100;
A = 8'h7A; B = 8'h8A; #100;
A = 8'h7A; B = 8'h8B; #100;
A = 8'h7A; B = 8'h8C; #100;
A = 8'h7A; B = 8'h8D; #100;
A = 8'h7A; B = 8'h8E; #100;
A = 8'h7A; B = 8'h8F; #100;
A = 8'h7A; B = 8'h90; #100;
A = 8'h7A; B = 8'h91; #100;
A = 8'h7A; B = 8'h92; #100;
A = 8'h7A; B = 8'h93; #100;
A = 8'h7A; B = 8'h94; #100;
A = 8'h7A; B = 8'h95; #100;
A = 8'h7A; B = 8'h96; #100;
A = 8'h7A; B = 8'h97; #100;
A = 8'h7A; B = 8'h98; #100;
A = 8'h7A; B = 8'h99; #100;
A = 8'h7A; B = 8'h9A; #100;
A = 8'h7A; B = 8'h9B; #100;
A = 8'h7A; B = 8'h9C; #100;
A = 8'h7A; B = 8'h9D; #100;
A = 8'h7A; B = 8'h9E; #100;
A = 8'h7A; B = 8'h9F; #100;
A = 8'h7A; B = 8'hA0; #100;
A = 8'h7A; B = 8'hA1; #100;
A = 8'h7A; B = 8'hA2; #100;
A = 8'h7A; B = 8'hA3; #100;
A = 8'h7A; B = 8'hA4; #100;
A = 8'h7A; B = 8'hA5; #100;
A = 8'h7A; B = 8'hA6; #100;
A = 8'h7A; B = 8'hA7; #100;
A = 8'h7A; B = 8'hA8; #100;
A = 8'h7A; B = 8'hA9; #100;
A = 8'h7A; B = 8'hAA; #100;
A = 8'h7A; B = 8'hAB; #100;
A = 8'h7A; B = 8'hAC; #100;
A = 8'h7A; B = 8'hAD; #100;
A = 8'h7A; B = 8'hAE; #100;
A = 8'h7A; B = 8'hAF; #100;
A = 8'h7A; B = 8'hB0; #100;
A = 8'h7A; B = 8'hB1; #100;
A = 8'h7A; B = 8'hB2; #100;
A = 8'h7A; B = 8'hB3; #100;
A = 8'h7A; B = 8'hB4; #100;
A = 8'h7A; B = 8'hB5; #100;
A = 8'h7A; B = 8'hB6; #100;
A = 8'h7A; B = 8'hB7; #100;
A = 8'h7A; B = 8'hB8; #100;
A = 8'h7A; B = 8'hB9; #100;
A = 8'h7A; B = 8'hBA; #100;
A = 8'h7A; B = 8'hBB; #100;
A = 8'h7A; B = 8'hBC; #100;
A = 8'h7A; B = 8'hBD; #100;
A = 8'h7A; B = 8'hBE; #100;
A = 8'h7A; B = 8'hBF; #100;
A = 8'h7A; B = 8'hC0; #100;
A = 8'h7A; B = 8'hC1; #100;
A = 8'h7A; B = 8'hC2; #100;
A = 8'h7A; B = 8'hC3; #100;
A = 8'h7A; B = 8'hC4; #100;
A = 8'h7A; B = 8'hC5; #100;
A = 8'h7A; B = 8'hC6; #100;
A = 8'h7A; B = 8'hC7; #100;
A = 8'h7A; B = 8'hC8; #100;
A = 8'h7A; B = 8'hC9; #100;
A = 8'h7A; B = 8'hCA; #100;
A = 8'h7A; B = 8'hCB; #100;
A = 8'h7A; B = 8'hCC; #100;
A = 8'h7A; B = 8'hCD; #100;
A = 8'h7A; B = 8'hCE; #100;
A = 8'h7A; B = 8'hCF; #100;
A = 8'h7A; B = 8'hD0; #100;
A = 8'h7A; B = 8'hD1; #100;
A = 8'h7A; B = 8'hD2; #100;
A = 8'h7A; B = 8'hD3; #100;
A = 8'h7A; B = 8'hD4; #100;
A = 8'h7A; B = 8'hD5; #100;
A = 8'h7A; B = 8'hD6; #100;
A = 8'h7A; B = 8'hD7; #100;
A = 8'h7A; B = 8'hD8; #100;
A = 8'h7A; B = 8'hD9; #100;
A = 8'h7A; B = 8'hDA; #100;
A = 8'h7A; B = 8'hDB; #100;
A = 8'h7A; B = 8'hDC; #100;
A = 8'h7A; B = 8'hDD; #100;
A = 8'h7A; B = 8'hDE; #100;
A = 8'h7A; B = 8'hDF; #100;
A = 8'h7A; B = 8'hE0; #100;
A = 8'h7A; B = 8'hE1; #100;
A = 8'h7A; B = 8'hE2; #100;
A = 8'h7A; B = 8'hE3; #100;
A = 8'h7A; B = 8'hE4; #100;
A = 8'h7A; B = 8'hE5; #100;
A = 8'h7A; B = 8'hE6; #100;
A = 8'h7A; B = 8'hE7; #100;
A = 8'h7A; B = 8'hE8; #100;
A = 8'h7A; B = 8'hE9; #100;
A = 8'h7A; B = 8'hEA; #100;
A = 8'h7A; B = 8'hEB; #100;
A = 8'h7A; B = 8'hEC; #100;
A = 8'h7A; B = 8'hED; #100;
A = 8'h7A; B = 8'hEE; #100;
A = 8'h7A; B = 8'hEF; #100;
A = 8'h7A; B = 8'hF0; #100;
A = 8'h7A; B = 8'hF1; #100;
A = 8'h7A; B = 8'hF2; #100;
A = 8'h7A; B = 8'hF3; #100;
A = 8'h7A; B = 8'hF4; #100;
A = 8'h7A; B = 8'hF5; #100;
A = 8'h7A; B = 8'hF6; #100;
A = 8'h7A; B = 8'hF7; #100;
A = 8'h7A; B = 8'hF8; #100;
A = 8'h7A; B = 8'hF9; #100;
A = 8'h7A; B = 8'hFA; #100;
A = 8'h7A; B = 8'hFB; #100;
A = 8'h7A; B = 8'hFC; #100;
A = 8'h7A; B = 8'hFD; #100;
A = 8'h7A; B = 8'hFE; #100;
A = 8'h7A; B = 8'hFF; #100;
A = 8'h7B; B = 8'h0; #100;
A = 8'h7B; B = 8'h1; #100;
A = 8'h7B; B = 8'h2; #100;
A = 8'h7B; B = 8'h3; #100;
A = 8'h7B; B = 8'h4; #100;
A = 8'h7B; B = 8'h5; #100;
A = 8'h7B; B = 8'h6; #100;
A = 8'h7B; B = 8'h7; #100;
A = 8'h7B; B = 8'h8; #100;
A = 8'h7B; B = 8'h9; #100;
A = 8'h7B; B = 8'hA; #100;
A = 8'h7B; B = 8'hB; #100;
A = 8'h7B; B = 8'hC; #100;
A = 8'h7B; B = 8'hD; #100;
A = 8'h7B; B = 8'hE; #100;
A = 8'h7B; B = 8'hF; #100;
A = 8'h7B; B = 8'h10; #100;
A = 8'h7B; B = 8'h11; #100;
A = 8'h7B; B = 8'h12; #100;
A = 8'h7B; B = 8'h13; #100;
A = 8'h7B; B = 8'h14; #100;
A = 8'h7B; B = 8'h15; #100;
A = 8'h7B; B = 8'h16; #100;
A = 8'h7B; B = 8'h17; #100;
A = 8'h7B; B = 8'h18; #100;
A = 8'h7B; B = 8'h19; #100;
A = 8'h7B; B = 8'h1A; #100;
A = 8'h7B; B = 8'h1B; #100;
A = 8'h7B; B = 8'h1C; #100;
A = 8'h7B; B = 8'h1D; #100;
A = 8'h7B; B = 8'h1E; #100;
A = 8'h7B; B = 8'h1F; #100;
A = 8'h7B; B = 8'h20; #100;
A = 8'h7B; B = 8'h21; #100;
A = 8'h7B; B = 8'h22; #100;
A = 8'h7B; B = 8'h23; #100;
A = 8'h7B; B = 8'h24; #100;
A = 8'h7B; B = 8'h25; #100;
A = 8'h7B; B = 8'h26; #100;
A = 8'h7B; B = 8'h27; #100;
A = 8'h7B; B = 8'h28; #100;
A = 8'h7B; B = 8'h29; #100;
A = 8'h7B; B = 8'h2A; #100;
A = 8'h7B; B = 8'h2B; #100;
A = 8'h7B; B = 8'h2C; #100;
A = 8'h7B; B = 8'h2D; #100;
A = 8'h7B; B = 8'h2E; #100;
A = 8'h7B; B = 8'h2F; #100;
A = 8'h7B; B = 8'h30; #100;
A = 8'h7B; B = 8'h31; #100;
A = 8'h7B; B = 8'h32; #100;
A = 8'h7B; B = 8'h33; #100;
A = 8'h7B; B = 8'h34; #100;
A = 8'h7B; B = 8'h35; #100;
A = 8'h7B; B = 8'h36; #100;
A = 8'h7B; B = 8'h37; #100;
A = 8'h7B; B = 8'h38; #100;
A = 8'h7B; B = 8'h39; #100;
A = 8'h7B; B = 8'h3A; #100;
A = 8'h7B; B = 8'h3B; #100;
A = 8'h7B; B = 8'h3C; #100;
A = 8'h7B; B = 8'h3D; #100;
A = 8'h7B; B = 8'h3E; #100;
A = 8'h7B; B = 8'h3F; #100;
A = 8'h7B; B = 8'h40; #100;
A = 8'h7B; B = 8'h41; #100;
A = 8'h7B; B = 8'h42; #100;
A = 8'h7B; B = 8'h43; #100;
A = 8'h7B; B = 8'h44; #100;
A = 8'h7B; B = 8'h45; #100;
A = 8'h7B; B = 8'h46; #100;
A = 8'h7B; B = 8'h47; #100;
A = 8'h7B; B = 8'h48; #100;
A = 8'h7B; B = 8'h49; #100;
A = 8'h7B; B = 8'h4A; #100;
A = 8'h7B; B = 8'h4B; #100;
A = 8'h7B; B = 8'h4C; #100;
A = 8'h7B; B = 8'h4D; #100;
A = 8'h7B; B = 8'h4E; #100;
A = 8'h7B; B = 8'h4F; #100;
A = 8'h7B; B = 8'h50; #100;
A = 8'h7B; B = 8'h51; #100;
A = 8'h7B; B = 8'h52; #100;
A = 8'h7B; B = 8'h53; #100;
A = 8'h7B; B = 8'h54; #100;
A = 8'h7B; B = 8'h55; #100;
A = 8'h7B; B = 8'h56; #100;
A = 8'h7B; B = 8'h57; #100;
A = 8'h7B; B = 8'h58; #100;
A = 8'h7B; B = 8'h59; #100;
A = 8'h7B; B = 8'h5A; #100;
A = 8'h7B; B = 8'h5B; #100;
A = 8'h7B; B = 8'h5C; #100;
A = 8'h7B; B = 8'h5D; #100;
A = 8'h7B; B = 8'h5E; #100;
A = 8'h7B; B = 8'h5F; #100;
A = 8'h7B; B = 8'h60; #100;
A = 8'h7B; B = 8'h61; #100;
A = 8'h7B; B = 8'h62; #100;
A = 8'h7B; B = 8'h63; #100;
A = 8'h7B; B = 8'h64; #100;
A = 8'h7B; B = 8'h65; #100;
A = 8'h7B; B = 8'h66; #100;
A = 8'h7B; B = 8'h67; #100;
A = 8'h7B; B = 8'h68; #100;
A = 8'h7B; B = 8'h69; #100;
A = 8'h7B; B = 8'h6A; #100;
A = 8'h7B; B = 8'h6B; #100;
A = 8'h7B; B = 8'h6C; #100;
A = 8'h7B; B = 8'h6D; #100;
A = 8'h7B; B = 8'h6E; #100;
A = 8'h7B; B = 8'h6F; #100;
A = 8'h7B; B = 8'h70; #100;
A = 8'h7B; B = 8'h71; #100;
A = 8'h7B; B = 8'h72; #100;
A = 8'h7B; B = 8'h73; #100;
A = 8'h7B; B = 8'h74; #100;
A = 8'h7B; B = 8'h75; #100;
A = 8'h7B; B = 8'h76; #100;
A = 8'h7B; B = 8'h77; #100;
A = 8'h7B; B = 8'h78; #100;
A = 8'h7B; B = 8'h79; #100;
A = 8'h7B; B = 8'h7A; #100;
A = 8'h7B; B = 8'h7B; #100;
A = 8'h7B; B = 8'h7C; #100;
A = 8'h7B; B = 8'h7D; #100;
A = 8'h7B; B = 8'h7E; #100;
A = 8'h7B; B = 8'h7F; #100;
A = 8'h7B; B = 8'h80; #100;
A = 8'h7B; B = 8'h81; #100;
A = 8'h7B; B = 8'h82; #100;
A = 8'h7B; B = 8'h83; #100;
A = 8'h7B; B = 8'h84; #100;
A = 8'h7B; B = 8'h85; #100;
A = 8'h7B; B = 8'h86; #100;
A = 8'h7B; B = 8'h87; #100;
A = 8'h7B; B = 8'h88; #100;
A = 8'h7B; B = 8'h89; #100;
A = 8'h7B; B = 8'h8A; #100;
A = 8'h7B; B = 8'h8B; #100;
A = 8'h7B; B = 8'h8C; #100;
A = 8'h7B; B = 8'h8D; #100;
A = 8'h7B; B = 8'h8E; #100;
A = 8'h7B; B = 8'h8F; #100;
A = 8'h7B; B = 8'h90; #100;
A = 8'h7B; B = 8'h91; #100;
A = 8'h7B; B = 8'h92; #100;
A = 8'h7B; B = 8'h93; #100;
A = 8'h7B; B = 8'h94; #100;
A = 8'h7B; B = 8'h95; #100;
A = 8'h7B; B = 8'h96; #100;
A = 8'h7B; B = 8'h97; #100;
A = 8'h7B; B = 8'h98; #100;
A = 8'h7B; B = 8'h99; #100;
A = 8'h7B; B = 8'h9A; #100;
A = 8'h7B; B = 8'h9B; #100;
A = 8'h7B; B = 8'h9C; #100;
A = 8'h7B; B = 8'h9D; #100;
A = 8'h7B; B = 8'h9E; #100;
A = 8'h7B; B = 8'h9F; #100;
A = 8'h7B; B = 8'hA0; #100;
A = 8'h7B; B = 8'hA1; #100;
A = 8'h7B; B = 8'hA2; #100;
A = 8'h7B; B = 8'hA3; #100;
A = 8'h7B; B = 8'hA4; #100;
A = 8'h7B; B = 8'hA5; #100;
A = 8'h7B; B = 8'hA6; #100;
A = 8'h7B; B = 8'hA7; #100;
A = 8'h7B; B = 8'hA8; #100;
A = 8'h7B; B = 8'hA9; #100;
A = 8'h7B; B = 8'hAA; #100;
A = 8'h7B; B = 8'hAB; #100;
A = 8'h7B; B = 8'hAC; #100;
A = 8'h7B; B = 8'hAD; #100;
A = 8'h7B; B = 8'hAE; #100;
A = 8'h7B; B = 8'hAF; #100;
A = 8'h7B; B = 8'hB0; #100;
A = 8'h7B; B = 8'hB1; #100;
A = 8'h7B; B = 8'hB2; #100;
A = 8'h7B; B = 8'hB3; #100;
A = 8'h7B; B = 8'hB4; #100;
A = 8'h7B; B = 8'hB5; #100;
A = 8'h7B; B = 8'hB6; #100;
A = 8'h7B; B = 8'hB7; #100;
A = 8'h7B; B = 8'hB8; #100;
A = 8'h7B; B = 8'hB9; #100;
A = 8'h7B; B = 8'hBA; #100;
A = 8'h7B; B = 8'hBB; #100;
A = 8'h7B; B = 8'hBC; #100;
A = 8'h7B; B = 8'hBD; #100;
A = 8'h7B; B = 8'hBE; #100;
A = 8'h7B; B = 8'hBF; #100;
A = 8'h7B; B = 8'hC0; #100;
A = 8'h7B; B = 8'hC1; #100;
A = 8'h7B; B = 8'hC2; #100;
A = 8'h7B; B = 8'hC3; #100;
A = 8'h7B; B = 8'hC4; #100;
A = 8'h7B; B = 8'hC5; #100;
A = 8'h7B; B = 8'hC6; #100;
A = 8'h7B; B = 8'hC7; #100;
A = 8'h7B; B = 8'hC8; #100;
A = 8'h7B; B = 8'hC9; #100;
A = 8'h7B; B = 8'hCA; #100;
A = 8'h7B; B = 8'hCB; #100;
A = 8'h7B; B = 8'hCC; #100;
A = 8'h7B; B = 8'hCD; #100;
A = 8'h7B; B = 8'hCE; #100;
A = 8'h7B; B = 8'hCF; #100;
A = 8'h7B; B = 8'hD0; #100;
A = 8'h7B; B = 8'hD1; #100;
A = 8'h7B; B = 8'hD2; #100;
A = 8'h7B; B = 8'hD3; #100;
A = 8'h7B; B = 8'hD4; #100;
A = 8'h7B; B = 8'hD5; #100;
A = 8'h7B; B = 8'hD6; #100;
A = 8'h7B; B = 8'hD7; #100;
A = 8'h7B; B = 8'hD8; #100;
A = 8'h7B; B = 8'hD9; #100;
A = 8'h7B; B = 8'hDA; #100;
A = 8'h7B; B = 8'hDB; #100;
A = 8'h7B; B = 8'hDC; #100;
A = 8'h7B; B = 8'hDD; #100;
A = 8'h7B; B = 8'hDE; #100;
A = 8'h7B; B = 8'hDF; #100;
A = 8'h7B; B = 8'hE0; #100;
A = 8'h7B; B = 8'hE1; #100;
A = 8'h7B; B = 8'hE2; #100;
A = 8'h7B; B = 8'hE3; #100;
A = 8'h7B; B = 8'hE4; #100;
A = 8'h7B; B = 8'hE5; #100;
A = 8'h7B; B = 8'hE6; #100;
A = 8'h7B; B = 8'hE7; #100;
A = 8'h7B; B = 8'hE8; #100;
A = 8'h7B; B = 8'hE9; #100;
A = 8'h7B; B = 8'hEA; #100;
A = 8'h7B; B = 8'hEB; #100;
A = 8'h7B; B = 8'hEC; #100;
A = 8'h7B; B = 8'hED; #100;
A = 8'h7B; B = 8'hEE; #100;
A = 8'h7B; B = 8'hEF; #100;
A = 8'h7B; B = 8'hF0; #100;
A = 8'h7B; B = 8'hF1; #100;
A = 8'h7B; B = 8'hF2; #100;
A = 8'h7B; B = 8'hF3; #100;
A = 8'h7B; B = 8'hF4; #100;
A = 8'h7B; B = 8'hF5; #100;
A = 8'h7B; B = 8'hF6; #100;
A = 8'h7B; B = 8'hF7; #100;
A = 8'h7B; B = 8'hF8; #100;
A = 8'h7B; B = 8'hF9; #100;
A = 8'h7B; B = 8'hFA; #100;
A = 8'h7B; B = 8'hFB; #100;
A = 8'h7B; B = 8'hFC; #100;
A = 8'h7B; B = 8'hFD; #100;
A = 8'h7B; B = 8'hFE; #100;
A = 8'h7B; B = 8'hFF; #100;
A = 8'h7C; B = 8'h0; #100;
A = 8'h7C; B = 8'h1; #100;
A = 8'h7C; B = 8'h2; #100;
A = 8'h7C; B = 8'h3; #100;
A = 8'h7C; B = 8'h4; #100;
A = 8'h7C; B = 8'h5; #100;
A = 8'h7C; B = 8'h6; #100;
A = 8'h7C; B = 8'h7; #100;
A = 8'h7C; B = 8'h8; #100;
A = 8'h7C; B = 8'h9; #100;
A = 8'h7C; B = 8'hA; #100;
A = 8'h7C; B = 8'hB; #100;
A = 8'h7C; B = 8'hC; #100;
A = 8'h7C; B = 8'hD; #100;
A = 8'h7C; B = 8'hE; #100;
A = 8'h7C; B = 8'hF; #100;
A = 8'h7C; B = 8'h10; #100;
A = 8'h7C; B = 8'h11; #100;
A = 8'h7C; B = 8'h12; #100;
A = 8'h7C; B = 8'h13; #100;
A = 8'h7C; B = 8'h14; #100;
A = 8'h7C; B = 8'h15; #100;
A = 8'h7C; B = 8'h16; #100;
A = 8'h7C; B = 8'h17; #100;
A = 8'h7C; B = 8'h18; #100;
A = 8'h7C; B = 8'h19; #100;
A = 8'h7C; B = 8'h1A; #100;
A = 8'h7C; B = 8'h1B; #100;
A = 8'h7C; B = 8'h1C; #100;
A = 8'h7C; B = 8'h1D; #100;
A = 8'h7C; B = 8'h1E; #100;
A = 8'h7C; B = 8'h1F; #100;
A = 8'h7C; B = 8'h20; #100;
A = 8'h7C; B = 8'h21; #100;
A = 8'h7C; B = 8'h22; #100;
A = 8'h7C; B = 8'h23; #100;
A = 8'h7C; B = 8'h24; #100;
A = 8'h7C; B = 8'h25; #100;
A = 8'h7C; B = 8'h26; #100;
A = 8'h7C; B = 8'h27; #100;
A = 8'h7C; B = 8'h28; #100;
A = 8'h7C; B = 8'h29; #100;
A = 8'h7C; B = 8'h2A; #100;
A = 8'h7C; B = 8'h2B; #100;
A = 8'h7C; B = 8'h2C; #100;
A = 8'h7C; B = 8'h2D; #100;
A = 8'h7C; B = 8'h2E; #100;
A = 8'h7C; B = 8'h2F; #100;
A = 8'h7C; B = 8'h30; #100;
A = 8'h7C; B = 8'h31; #100;
A = 8'h7C; B = 8'h32; #100;
A = 8'h7C; B = 8'h33; #100;
A = 8'h7C; B = 8'h34; #100;
A = 8'h7C; B = 8'h35; #100;
A = 8'h7C; B = 8'h36; #100;
A = 8'h7C; B = 8'h37; #100;
A = 8'h7C; B = 8'h38; #100;
A = 8'h7C; B = 8'h39; #100;
A = 8'h7C; B = 8'h3A; #100;
A = 8'h7C; B = 8'h3B; #100;
A = 8'h7C; B = 8'h3C; #100;
A = 8'h7C; B = 8'h3D; #100;
A = 8'h7C; B = 8'h3E; #100;
A = 8'h7C; B = 8'h3F; #100;
A = 8'h7C; B = 8'h40; #100;
A = 8'h7C; B = 8'h41; #100;
A = 8'h7C; B = 8'h42; #100;
A = 8'h7C; B = 8'h43; #100;
A = 8'h7C; B = 8'h44; #100;
A = 8'h7C; B = 8'h45; #100;
A = 8'h7C; B = 8'h46; #100;
A = 8'h7C; B = 8'h47; #100;
A = 8'h7C; B = 8'h48; #100;
A = 8'h7C; B = 8'h49; #100;
A = 8'h7C; B = 8'h4A; #100;
A = 8'h7C; B = 8'h4B; #100;
A = 8'h7C; B = 8'h4C; #100;
A = 8'h7C; B = 8'h4D; #100;
A = 8'h7C; B = 8'h4E; #100;
A = 8'h7C; B = 8'h4F; #100;
A = 8'h7C; B = 8'h50; #100;
A = 8'h7C; B = 8'h51; #100;
A = 8'h7C; B = 8'h52; #100;
A = 8'h7C; B = 8'h53; #100;
A = 8'h7C; B = 8'h54; #100;
A = 8'h7C; B = 8'h55; #100;
A = 8'h7C; B = 8'h56; #100;
A = 8'h7C; B = 8'h57; #100;
A = 8'h7C; B = 8'h58; #100;
A = 8'h7C; B = 8'h59; #100;
A = 8'h7C; B = 8'h5A; #100;
A = 8'h7C; B = 8'h5B; #100;
A = 8'h7C; B = 8'h5C; #100;
A = 8'h7C; B = 8'h5D; #100;
A = 8'h7C; B = 8'h5E; #100;
A = 8'h7C; B = 8'h5F; #100;
A = 8'h7C; B = 8'h60; #100;
A = 8'h7C; B = 8'h61; #100;
A = 8'h7C; B = 8'h62; #100;
A = 8'h7C; B = 8'h63; #100;
A = 8'h7C; B = 8'h64; #100;
A = 8'h7C; B = 8'h65; #100;
A = 8'h7C; B = 8'h66; #100;
A = 8'h7C; B = 8'h67; #100;
A = 8'h7C; B = 8'h68; #100;
A = 8'h7C; B = 8'h69; #100;
A = 8'h7C; B = 8'h6A; #100;
A = 8'h7C; B = 8'h6B; #100;
A = 8'h7C; B = 8'h6C; #100;
A = 8'h7C; B = 8'h6D; #100;
A = 8'h7C; B = 8'h6E; #100;
A = 8'h7C; B = 8'h6F; #100;
A = 8'h7C; B = 8'h70; #100;
A = 8'h7C; B = 8'h71; #100;
A = 8'h7C; B = 8'h72; #100;
A = 8'h7C; B = 8'h73; #100;
A = 8'h7C; B = 8'h74; #100;
A = 8'h7C; B = 8'h75; #100;
A = 8'h7C; B = 8'h76; #100;
A = 8'h7C; B = 8'h77; #100;
A = 8'h7C; B = 8'h78; #100;
A = 8'h7C; B = 8'h79; #100;
A = 8'h7C; B = 8'h7A; #100;
A = 8'h7C; B = 8'h7B; #100;
A = 8'h7C; B = 8'h7C; #100;
A = 8'h7C; B = 8'h7D; #100;
A = 8'h7C; B = 8'h7E; #100;
A = 8'h7C; B = 8'h7F; #100;
A = 8'h7C; B = 8'h80; #100;
A = 8'h7C; B = 8'h81; #100;
A = 8'h7C; B = 8'h82; #100;
A = 8'h7C; B = 8'h83; #100;
A = 8'h7C; B = 8'h84; #100;
A = 8'h7C; B = 8'h85; #100;
A = 8'h7C; B = 8'h86; #100;
A = 8'h7C; B = 8'h87; #100;
A = 8'h7C; B = 8'h88; #100;
A = 8'h7C; B = 8'h89; #100;
A = 8'h7C; B = 8'h8A; #100;
A = 8'h7C; B = 8'h8B; #100;
A = 8'h7C; B = 8'h8C; #100;
A = 8'h7C; B = 8'h8D; #100;
A = 8'h7C; B = 8'h8E; #100;
A = 8'h7C; B = 8'h8F; #100;
A = 8'h7C; B = 8'h90; #100;
A = 8'h7C; B = 8'h91; #100;
A = 8'h7C; B = 8'h92; #100;
A = 8'h7C; B = 8'h93; #100;
A = 8'h7C; B = 8'h94; #100;
A = 8'h7C; B = 8'h95; #100;
A = 8'h7C; B = 8'h96; #100;
A = 8'h7C; B = 8'h97; #100;
A = 8'h7C; B = 8'h98; #100;
A = 8'h7C; B = 8'h99; #100;
A = 8'h7C; B = 8'h9A; #100;
A = 8'h7C; B = 8'h9B; #100;
A = 8'h7C; B = 8'h9C; #100;
A = 8'h7C; B = 8'h9D; #100;
A = 8'h7C; B = 8'h9E; #100;
A = 8'h7C; B = 8'h9F; #100;
A = 8'h7C; B = 8'hA0; #100;
A = 8'h7C; B = 8'hA1; #100;
A = 8'h7C; B = 8'hA2; #100;
A = 8'h7C; B = 8'hA3; #100;
A = 8'h7C; B = 8'hA4; #100;
A = 8'h7C; B = 8'hA5; #100;
A = 8'h7C; B = 8'hA6; #100;
A = 8'h7C; B = 8'hA7; #100;
A = 8'h7C; B = 8'hA8; #100;
A = 8'h7C; B = 8'hA9; #100;
A = 8'h7C; B = 8'hAA; #100;
A = 8'h7C; B = 8'hAB; #100;
A = 8'h7C; B = 8'hAC; #100;
A = 8'h7C; B = 8'hAD; #100;
A = 8'h7C; B = 8'hAE; #100;
A = 8'h7C; B = 8'hAF; #100;
A = 8'h7C; B = 8'hB0; #100;
A = 8'h7C; B = 8'hB1; #100;
A = 8'h7C; B = 8'hB2; #100;
A = 8'h7C; B = 8'hB3; #100;
A = 8'h7C; B = 8'hB4; #100;
A = 8'h7C; B = 8'hB5; #100;
A = 8'h7C; B = 8'hB6; #100;
A = 8'h7C; B = 8'hB7; #100;
A = 8'h7C; B = 8'hB8; #100;
A = 8'h7C; B = 8'hB9; #100;
A = 8'h7C; B = 8'hBA; #100;
A = 8'h7C; B = 8'hBB; #100;
A = 8'h7C; B = 8'hBC; #100;
A = 8'h7C; B = 8'hBD; #100;
A = 8'h7C; B = 8'hBE; #100;
A = 8'h7C; B = 8'hBF; #100;
A = 8'h7C; B = 8'hC0; #100;
A = 8'h7C; B = 8'hC1; #100;
A = 8'h7C; B = 8'hC2; #100;
A = 8'h7C; B = 8'hC3; #100;
A = 8'h7C; B = 8'hC4; #100;
A = 8'h7C; B = 8'hC5; #100;
A = 8'h7C; B = 8'hC6; #100;
A = 8'h7C; B = 8'hC7; #100;
A = 8'h7C; B = 8'hC8; #100;
A = 8'h7C; B = 8'hC9; #100;
A = 8'h7C; B = 8'hCA; #100;
A = 8'h7C; B = 8'hCB; #100;
A = 8'h7C; B = 8'hCC; #100;
A = 8'h7C; B = 8'hCD; #100;
A = 8'h7C; B = 8'hCE; #100;
A = 8'h7C; B = 8'hCF; #100;
A = 8'h7C; B = 8'hD0; #100;
A = 8'h7C; B = 8'hD1; #100;
A = 8'h7C; B = 8'hD2; #100;
A = 8'h7C; B = 8'hD3; #100;
A = 8'h7C; B = 8'hD4; #100;
A = 8'h7C; B = 8'hD5; #100;
A = 8'h7C; B = 8'hD6; #100;
A = 8'h7C; B = 8'hD7; #100;
A = 8'h7C; B = 8'hD8; #100;
A = 8'h7C; B = 8'hD9; #100;
A = 8'h7C; B = 8'hDA; #100;
A = 8'h7C; B = 8'hDB; #100;
A = 8'h7C; B = 8'hDC; #100;
A = 8'h7C; B = 8'hDD; #100;
A = 8'h7C; B = 8'hDE; #100;
A = 8'h7C; B = 8'hDF; #100;
A = 8'h7C; B = 8'hE0; #100;
A = 8'h7C; B = 8'hE1; #100;
A = 8'h7C; B = 8'hE2; #100;
A = 8'h7C; B = 8'hE3; #100;
A = 8'h7C; B = 8'hE4; #100;
A = 8'h7C; B = 8'hE5; #100;
A = 8'h7C; B = 8'hE6; #100;
A = 8'h7C; B = 8'hE7; #100;
A = 8'h7C; B = 8'hE8; #100;
A = 8'h7C; B = 8'hE9; #100;
A = 8'h7C; B = 8'hEA; #100;
A = 8'h7C; B = 8'hEB; #100;
A = 8'h7C; B = 8'hEC; #100;
A = 8'h7C; B = 8'hED; #100;
A = 8'h7C; B = 8'hEE; #100;
A = 8'h7C; B = 8'hEF; #100;
A = 8'h7C; B = 8'hF0; #100;
A = 8'h7C; B = 8'hF1; #100;
A = 8'h7C; B = 8'hF2; #100;
A = 8'h7C; B = 8'hF3; #100;
A = 8'h7C; B = 8'hF4; #100;
A = 8'h7C; B = 8'hF5; #100;
A = 8'h7C; B = 8'hF6; #100;
A = 8'h7C; B = 8'hF7; #100;
A = 8'h7C; B = 8'hF8; #100;
A = 8'h7C; B = 8'hF9; #100;
A = 8'h7C; B = 8'hFA; #100;
A = 8'h7C; B = 8'hFB; #100;
A = 8'h7C; B = 8'hFC; #100;
A = 8'h7C; B = 8'hFD; #100;
A = 8'h7C; B = 8'hFE; #100;
A = 8'h7C; B = 8'hFF; #100;
A = 8'h7D; B = 8'h0; #100;
A = 8'h7D; B = 8'h1; #100;
A = 8'h7D; B = 8'h2; #100;
A = 8'h7D; B = 8'h3; #100;
A = 8'h7D; B = 8'h4; #100;
A = 8'h7D; B = 8'h5; #100;
A = 8'h7D; B = 8'h6; #100;
A = 8'h7D; B = 8'h7; #100;
A = 8'h7D; B = 8'h8; #100;
A = 8'h7D; B = 8'h9; #100;
A = 8'h7D; B = 8'hA; #100;
A = 8'h7D; B = 8'hB; #100;
A = 8'h7D; B = 8'hC; #100;
A = 8'h7D; B = 8'hD; #100;
A = 8'h7D; B = 8'hE; #100;
A = 8'h7D; B = 8'hF; #100;
A = 8'h7D; B = 8'h10; #100;
A = 8'h7D; B = 8'h11; #100;
A = 8'h7D; B = 8'h12; #100;
A = 8'h7D; B = 8'h13; #100;
A = 8'h7D; B = 8'h14; #100;
A = 8'h7D; B = 8'h15; #100;
A = 8'h7D; B = 8'h16; #100;
A = 8'h7D; B = 8'h17; #100;
A = 8'h7D; B = 8'h18; #100;
A = 8'h7D; B = 8'h19; #100;
A = 8'h7D; B = 8'h1A; #100;
A = 8'h7D; B = 8'h1B; #100;
A = 8'h7D; B = 8'h1C; #100;
A = 8'h7D; B = 8'h1D; #100;
A = 8'h7D; B = 8'h1E; #100;
A = 8'h7D; B = 8'h1F; #100;
A = 8'h7D; B = 8'h20; #100;
A = 8'h7D; B = 8'h21; #100;
A = 8'h7D; B = 8'h22; #100;
A = 8'h7D; B = 8'h23; #100;
A = 8'h7D; B = 8'h24; #100;
A = 8'h7D; B = 8'h25; #100;
A = 8'h7D; B = 8'h26; #100;
A = 8'h7D; B = 8'h27; #100;
A = 8'h7D; B = 8'h28; #100;
A = 8'h7D; B = 8'h29; #100;
A = 8'h7D; B = 8'h2A; #100;
A = 8'h7D; B = 8'h2B; #100;
A = 8'h7D; B = 8'h2C; #100;
A = 8'h7D; B = 8'h2D; #100;
A = 8'h7D; B = 8'h2E; #100;
A = 8'h7D; B = 8'h2F; #100;
A = 8'h7D; B = 8'h30; #100;
A = 8'h7D; B = 8'h31; #100;
A = 8'h7D; B = 8'h32; #100;
A = 8'h7D; B = 8'h33; #100;
A = 8'h7D; B = 8'h34; #100;
A = 8'h7D; B = 8'h35; #100;
A = 8'h7D; B = 8'h36; #100;
A = 8'h7D; B = 8'h37; #100;
A = 8'h7D; B = 8'h38; #100;
A = 8'h7D; B = 8'h39; #100;
A = 8'h7D; B = 8'h3A; #100;
A = 8'h7D; B = 8'h3B; #100;
A = 8'h7D; B = 8'h3C; #100;
A = 8'h7D; B = 8'h3D; #100;
A = 8'h7D; B = 8'h3E; #100;
A = 8'h7D; B = 8'h3F; #100;
A = 8'h7D; B = 8'h40; #100;
A = 8'h7D; B = 8'h41; #100;
A = 8'h7D; B = 8'h42; #100;
A = 8'h7D; B = 8'h43; #100;
A = 8'h7D; B = 8'h44; #100;
A = 8'h7D; B = 8'h45; #100;
A = 8'h7D; B = 8'h46; #100;
A = 8'h7D; B = 8'h47; #100;
A = 8'h7D; B = 8'h48; #100;
A = 8'h7D; B = 8'h49; #100;
A = 8'h7D; B = 8'h4A; #100;
A = 8'h7D; B = 8'h4B; #100;
A = 8'h7D; B = 8'h4C; #100;
A = 8'h7D; B = 8'h4D; #100;
A = 8'h7D; B = 8'h4E; #100;
A = 8'h7D; B = 8'h4F; #100;
A = 8'h7D; B = 8'h50; #100;
A = 8'h7D; B = 8'h51; #100;
A = 8'h7D; B = 8'h52; #100;
A = 8'h7D; B = 8'h53; #100;
A = 8'h7D; B = 8'h54; #100;
A = 8'h7D; B = 8'h55; #100;
A = 8'h7D; B = 8'h56; #100;
A = 8'h7D; B = 8'h57; #100;
A = 8'h7D; B = 8'h58; #100;
A = 8'h7D; B = 8'h59; #100;
A = 8'h7D; B = 8'h5A; #100;
A = 8'h7D; B = 8'h5B; #100;
A = 8'h7D; B = 8'h5C; #100;
A = 8'h7D; B = 8'h5D; #100;
A = 8'h7D; B = 8'h5E; #100;
A = 8'h7D; B = 8'h5F; #100;
A = 8'h7D; B = 8'h60; #100;
A = 8'h7D; B = 8'h61; #100;
A = 8'h7D; B = 8'h62; #100;
A = 8'h7D; B = 8'h63; #100;
A = 8'h7D; B = 8'h64; #100;
A = 8'h7D; B = 8'h65; #100;
A = 8'h7D; B = 8'h66; #100;
A = 8'h7D; B = 8'h67; #100;
A = 8'h7D; B = 8'h68; #100;
A = 8'h7D; B = 8'h69; #100;
A = 8'h7D; B = 8'h6A; #100;
A = 8'h7D; B = 8'h6B; #100;
A = 8'h7D; B = 8'h6C; #100;
A = 8'h7D; B = 8'h6D; #100;
A = 8'h7D; B = 8'h6E; #100;
A = 8'h7D; B = 8'h6F; #100;
A = 8'h7D; B = 8'h70; #100;
A = 8'h7D; B = 8'h71; #100;
A = 8'h7D; B = 8'h72; #100;
A = 8'h7D; B = 8'h73; #100;
A = 8'h7D; B = 8'h74; #100;
A = 8'h7D; B = 8'h75; #100;
A = 8'h7D; B = 8'h76; #100;
A = 8'h7D; B = 8'h77; #100;
A = 8'h7D; B = 8'h78; #100;
A = 8'h7D; B = 8'h79; #100;
A = 8'h7D; B = 8'h7A; #100;
A = 8'h7D; B = 8'h7B; #100;
A = 8'h7D; B = 8'h7C; #100;
A = 8'h7D; B = 8'h7D; #100;
A = 8'h7D; B = 8'h7E; #100;
A = 8'h7D; B = 8'h7F; #100;
A = 8'h7D; B = 8'h80; #100;
A = 8'h7D; B = 8'h81; #100;
A = 8'h7D; B = 8'h82; #100;
A = 8'h7D; B = 8'h83; #100;
A = 8'h7D; B = 8'h84; #100;
A = 8'h7D; B = 8'h85; #100;
A = 8'h7D; B = 8'h86; #100;
A = 8'h7D; B = 8'h87; #100;
A = 8'h7D; B = 8'h88; #100;
A = 8'h7D; B = 8'h89; #100;
A = 8'h7D; B = 8'h8A; #100;
A = 8'h7D; B = 8'h8B; #100;
A = 8'h7D; B = 8'h8C; #100;
A = 8'h7D; B = 8'h8D; #100;
A = 8'h7D; B = 8'h8E; #100;
A = 8'h7D; B = 8'h8F; #100;
A = 8'h7D; B = 8'h90; #100;
A = 8'h7D; B = 8'h91; #100;
A = 8'h7D; B = 8'h92; #100;
A = 8'h7D; B = 8'h93; #100;
A = 8'h7D; B = 8'h94; #100;
A = 8'h7D; B = 8'h95; #100;
A = 8'h7D; B = 8'h96; #100;
A = 8'h7D; B = 8'h97; #100;
A = 8'h7D; B = 8'h98; #100;
A = 8'h7D; B = 8'h99; #100;
A = 8'h7D; B = 8'h9A; #100;
A = 8'h7D; B = 8'h9B; #100;
A = 8'h7D; B = 8'h9C; #100;
A = 8'h7D; B = 8'h9D; #100;
A = 8'h7D; B = 8'h9E; #100;
A = 8'h7D; B = 8'h9F; #100;
A = 8'h7D; B = 8'hA0; #100;
A = 8'h7D; B = 8'hA1; #100;
A = 8'h7D; B = 8'hA2; #100;
A = 8'h7D; B = 8'hA3; #100;
A = 8'h7D; B = 8'hA4; #100;
A = 8'h7D; B = 8'hA5; #100;
A = 8'h7D; B = 8'hA6; #100;
A = 8'h7D; B = 8'hA7; #100;
A = 8'h7D; B = 8'hA8; #100;
A = 8'h7D; B = 8'hA9; #100;
A = 8'h7D; B = 8'hAA; #100;
A = 8'h7D; B = 8'hAB; #100;
A = 8'h7D; B = 8'hAC; #100;
A = 8'h7D; B = 8'hAD; #100;
A = 8'h7D; B = 8'hAE; #100;
A = 8'h7D; B = 8'hAF; #100;
A = 8'h7D; B = 8'hB0; #100;
A = 8'h7D; B = 8'hB1; #100;
A = 8'h7D; B = 8'hB2; #100;
A = 8'h7D; B = 8'hB3; #100;
A = 8'h7D; B = 8'hB4; #100;
A = 8'h7D; B = 8'hB5; #100;
A = 8'h7D; B = 8'hB6; #100;
A = 8'h7D; B = 8'hB7; #100;
A = 8'h7D; B = 8'hB8; #100;
A = 8'h7D; B = 8'hB9; #100;
A = 8'h7D; B = 8'hBA; #100;
A = 8'h7D; B = 8'hBB; #100;
A = 8'h7D; B = 8'hBC; #100;
A = 8'h7D; B = 8'hBD; #100;
A = 8'h7D; B = 8'hBE; #100;
A = 8'h7D; B = 8'hBF; #100;
A = 8'h7D; B = 8'hC0; #100;
A = 8'h7D; B = 8'hC1; #100;
A = 8'h7D; B = 8'hC2; #100;
A = 8'h7D; B = 8'hC3; #100;
A = 8'h7D; B = 8'hC4; #100;
A = 8'h7D; B = 8'hC5; #100;
A = 8'h7D; B = 8'hC6; #100;
A = 8'h7D; B = 8'hC7; #100;
A = 8'h7D; B = 8'hC8; #100;
A = 8'h7D; B = 8'hC9; #100;
A = 8'h7D; B = 8'hCA; #100;
A = 8'h7D; B = 8'hCB; #100;
A = 8'h7D; B = 8'hCC; #100;
A = 8'h7D; B = 8'hCD; #100;
A = 8'h7D; B = 8'hCE; #100;
A = 8'h7D; B = 8'hCF; #100;
A = 8'h7D; B = 8'hD0; #100;
A = 8'h7D; B = 8'hD1; #100;
A = 8'h7D; B = 8'hD2; #100;
A = 8'h7D; B = 8'hD3; #100;
A = 8'h7D; B = 8'hD4; #100;
A = 8'h7D; B = 8'hD5; #100;
A = 8'h7D; B = 8'hD6; #100;
A = 8'h7D; B = 8'hD7; #100;
A = 8'h7D; B = 8'hD8; #100;
A = 8'h7D; B = 8'hD9; #100;
A = 8'h7D; B = 8'hDA; #100;
A = 8'h7D; B = 8'hDB; #100;
A = 8'h7D; B = 8'hDC; #100;
A = 8'h7D; B = 8'hDD; #100;
A = 8'h7D; B = 8'hDE; #100;
A = 8'h7D; B = 8'hDF; #100;
A = 8'h7D; B = 8'hE0; #100;
A = 8'h7D; B = 8'hE1; #100;
A = 8'h7D; B = 8'hE2; #100;
A = 8'h7D; B = 8'hE3; #100;
A = 8'h7D; B = 8'hE4; #100;
A = 8'h7D; B = 8'hE5; #100;
A = 8'h7D; B = 8'hE6; #100;
A = 8'h7D; B = 8'hE7; #100;
A = 8'h7D; B = 8'hE8; #100;
A = 8'h7D; B = 8'hE9; #100;
A = 8'h7D; B = 8'hEA; #100;
A = 8'h7D; B = 8'hEB; #100;
A = 8'h7D; B = 8'hEC; #100;
A = 8'h7D; B = 8'hED; #100;
A = 8'h7D; B = 8'hEE; #100;
A = 8'h7D; B = 8'hEF; #100;
A = 8'h7D; B = 8'hF0; #100;
A = 8'h7D; B = 8'hF1; #100;
A = 8'h7D; B = 8'hF2; #100;
A = 8'h7D; B = 8'hF3; #100;
A = 8'h7D; B = 8'hF4; #100;
A = 8'h7D; B = 8'hF5; #100;
A = 8'h7D; B = 8'hF6; #100;
A = 8'h7D; B = 8'hF7; #100;
A = 8'h7D; B = 8'hF8; #100;
A = 8'h7D; B = 8'hF9; #100;
A = 8'h7D; B = 8'hFA; #100;
A = 8'h7D; B = 8'hFB; #100;
A = 8'h7D; B = 8'hFC; #100;
A = 8'h7D; B = 8'hFD; #100;
A = 8'h7D; B = 8'hFE; #100;
A = 8'h7D; B = 8'hFF; #100;
A = 8'h7E; B = 8'h0; #100;
A = 8'h7E; B = 8'h1; #100;
A = 8'h7E; B = 8'h2; #100;
A = 8'h7E; B = 8'h3; #100;
A = 8'h7E; B = 8'h4; #100;
A = 8'h7E; B = 8'h5; #100;
A = 8'h7E; B = 8'h6; #100;
A = 8'h7E; B = 8'h7; #100;
A = 8'h7E; B = 8'h8; #100;
A = 8'h7E; B = 8'h9; #100;
A = 8'h7E; B = 8'hA; #100;
A = 8'h7E; B = 8'hB; #100;
A = 8'h7E; B = 8'hC; #100;
A = 8'h7E; B = 8'hD; #100;
A = 8'h7E; B = 8'hE; #100;
A = 8'h7E; B = 8'hF; #100;
A = 8'h7E; B = 8'h10; #100;
A = 8'h7E; B = 8'h11; #100;
A = 8'h7E; B = 8'h12; #100;
A = 8'h7E; B = 8'h13; #100;
A = 8'h7E; B = 8'h14; #100;
A = 8'h7E; B = 8'h15; #100;
A = 8'h7E; B = 8'h16; #100;
A = 8'h7E; B = 8'h17; #100;
A = 8'h7E; B = 8'h18; #100;
A = 8'h7E; B = 8'h19; #100;
A = 8'h7E; B = 8'h1A; #100;
A = 8'h7E; B = 8'h1B; #100;
A = 8'h7E; B = 8'h1C; #100;
A = 8'h7E; B = 8'h1D; #100;
A = 8'h7E; B = 8'h1E; #100;
A = 8'h7E; B = 8'h1F; #100;
A = 8'h7E; B = 8'h20; #100;
A = 8'h7E; B = 8'h21; #100;
A = 8'h7E; B = 8'h22; #100;
A = 8'h7E; B = 8'h23; #100;
A = 8'h7E; B = 8'h24; #100;
A = 8'h7E; B = 8'h25; #100;
A = 8'h7E; B = 8'h26; #100;
A = 8'h7E; B = 8'h27; #100;
A = 8'h7E; B = 8'h28; #100;
A = 8'h7E; B = 8'h29; #100;
A = 8'h7E; B = 8'h2A; #100;
A = 8'h7E; B = 8'h2B; #100;
A = 8'h7E; B = 8'h2C; #100;
A = 8'h7E; B = 8'h2D; #100;
A = 8'h7E; B = 8'h2E; #100;
A = 8'h7E; B = 8'h2F; #100;
A = 8'h7E; B = 8'h30; #100;
A = 8'h7E; B = 8'h31; #100;
A = 8'h7E; B = 8'h32; #100;
A = 8'h7E; B = 8'h33; #100;
A = 8'h7E; B = 8'h34; #100;
A = 8'h7E; B = 8'h35; #100;
A = 8'h7E; B = 8'h36; #100;
A = 8'h7E; B = 8'h37; #100;
A = 8'h7E; B = 8'h38; #100;
A = 8'h7E; B = 8'h39; #100;
A = 8'h7E; B = 8'h3A; #100;
A = 8'h7E; B = 8'h3B; #100;
A = 8'h7E; B = 8'h3C; #100;
A = 8'h7E; B = 8'h3D; #100;
A = 8'h7E; B = 8'h3E; #100;
A = 8'h7E; B = 8'h3F; #100;
A = 8'h7E; B = 8'h40; #100;
A = 8'h7E; B = 8'h41; #100;
A = 8'h7E; B = 8'h42; #100;
A = 8'h7E; B = 8'h43; #100;
A = 8'h7E; B = 8'h44; #100;
A = 8'h7E; B = 8'h45; #100;
A = 8'h7E; B = 8'h46; #100;
A = 8'h7E; B = 8'h47; #100;
A = 8'h7E; B = 8'h48; #100;
A = 8'h7E; B = 8'h49; #100;
A = 8'h7E; B = 8'h4A; #100;
A = 8'h7E; B = 8'h4B; #100;
A = 8'h7E; B = 8'h4C; #100;
A = 8'h7E; B = 8'h4D; #100;
A = 8'h7E; B = 8'h4E; #100;
A = 8'h7E; B = 8'h4F; #100;
A = 8'h7E; B = 8'h50; #100;
A = 8'h7E; B = 8'h51; #100;
A = 8'h7E; B = 8'h52; #100;
A = 8'h7E; B = 8'h53; #100;
A = 8'h7E; B = 8'h54; #100;
A = 8'h7E; B = 8'h55; #100;
A = 8'h7E; B = 8'h56; #100;
A = 8'h7E; B = 8'h57; #100;
A = 8'h7E; B = 8'h58; #100;
A = 8'h7E; B = 8'h59; #100;
A = 8'h7E; B = 8'h5A; #100;
A = 8'h7E; B = 8'h5B; #100;
A = 8'h7E; B = 8'h5C; #100;
A = 8'h7E; B = 8'h5D; #100;
A = 8'h7E; B = 8'h5E; #100;
A = 8'h7E; B = 8'h5F; #100;
A = 8'h7E; B = 8'h60; #100;
A = 8'h7E; B = 8'h61; #100;
A = 8'h7E; B = 8'h62; #100;
A = 8'h7E; B = 8'h63; #100;
A = 8'h7E; B = 8'h64; #100;
A = 8'h7E; B = 8'h65; #100;
A = 8'h7E; B = 8'h66; #100;
A = 8'h7E; B = 8'h67; #100;
A = 8'h7E; B = 8'h68; #100;
A = 8'h7E; B = 8'h69; #100;
A = 8'h7E; B = 8'h6A; #100;
A = 8'h7E; B = 8'h6B; #100;
A = 8'h7E; B = 8'h6C; #100;
A = 8'h7E; B = 8'h6D; #100;
A = 8'h7E; B = 8'h6E; #100;
A = 8'h7E; B = 8'h6F; #100;
A = 8'h7E; B = 8'h70; #100;
A = 8'h7E; B = 8'h71; #100;
A = 8'h7E; B = 8'h72; #100;
A = 8'h7E; B = 8'h73; #100;
A = 8'h7E; B = 8'h74; #100;
A = 8'h7E; B = 8'h75; #100;
A = 8'h7E; B = 8'h76; #100;
A = 8'h7E; B = 8'h77; #100;
A = 8'h7E; B = 8'h78; #100;
A = 8'h7E; B = 8'h79; #100;
A = 8'h7E; B = 8'h7A; #100;
A = 8'h7E; B = 8'h7B; #100;
A = 8'h7E; B = 8'h7C; #100;
A = 8'h7E; B = 8'h7D; #100;
A = 8'h7E; B = 8'h7E; #100;
A = 8'h7E; B = 8'h7F; #100;
A = 8'h7E; B = 8'h80; #100;
A = 8'h7E; B = 8'h81; #100;
A = 8'h7E; B = 8'h82; #100;
A = 8'h7E; B = 8'h83; #100;
A = 8'h7E; B = 8'h84; #100;
A = 8'h7E; B = 8'h85; #100;
A = 8'h7E; B = 8'h86; #100;
A = 8'h7E; B = 8'h87; #100;
A = 8'h7E; B = 8'h88; #100;
A = 8'h7E; B = 8'h89; #100;
A = 8'h7E; B = 8'h8A; #100;
A = 8'h7E; B = 8'h8B; #100;
A = 8'h7E; B = 8'h8C; #100;
A = 8'h7E; B = 8'h8D; #100;
A = 8'h7E; B = 8'h8E; #100;
A = 8'h7E; B = 8'h8F; #100;
A = 8'h7E; B = 8'h90; #100;
A = 8'h7E; B = 8'h91; #100;
A = 8'h7E; B = 8'h92; #100;
A = 8'h7E; B = 8'h93; #100;
A = 8'h7E; B = 8'h94; #100;
A = 8'h7E; B = 8'h95; #100;
A = 8'h7E; B = 8'h96; #100;
A = 8'h7E; B = 8'h97; #100;
A = 8'h7E; B = 8'h98; #100;
A = 8'h7E; B = 8'h99; #100;
A = 8'h7E; B = 8'h9A; #100;
A = 8'h7E; B = 8'h9B; #100;
A = 8'h7E; B = 8'h9C; #100;
A = 8'h7E; B = 8'h9D; #100;
A = 8'h7E; B = 8'h9E; #100;
A = 8'h7E; B = 8'h9F; #100;
A = 8'h7E; B = 8'hA0; #100;
A = 8'h7E; B = 8'hA1; #100;
A = 8'h7E; B = 8'hA2; #100;
A = 8'h7E; B = 8'hA3; #100;
A = 8'h7E; B = 8'hA4; #100;
A = 8'h7E; B = 8'hA5; #100;
A = 8'h7E; B = 8'hA6; #100;
A = 8'h7E; B = 8'hA7; #100;
A = 8'h7E; B = 8'hA8; #100;
A = 8'h7E; B = 8'hA9; #100;
A = 8'h7E; B = 8'hAA; #100;
A = 8'h7E; B = 8'hAB; #100;
A = 8'h7E; B = 8'hAC; #100;
A = 8'h7E; B = 8'hAD; #100;
A = 8'h7E; B = 8'hAE; #100;
A = 8'h7E; B = 8'hAF; #100;
A = 8'h7E; B = 8'hB0; #100;
A = 8'h7E; B = 8'hB1; #100;
A = 8'h7E; B = 8'hB2; #100;
A = 8'h7E; B = 8'hB3; #100;
A = 8'h7E; B = 8'hB4; #100;
A = 8'h7E; B = 8'hB5; #100;
A = 8'h7E; B = 8'hB6; #100;
A = 8'h7E; B = 8'hB7; #100;
A = 8'h7E; B = 8'hB8; #100;
A = 8'h7E; B = 8'hB9; #100;
A = 8'h7E; B = 8'hBA; #100;
A = 8'h7E; B = 8'hBB; #100;
A = 8'h7E; B = 8'hBC; #100;
A = 8'h7E; B = 8'hBD; #100;
A = 8'h7E; B = 8'hBE; #100;
A = 8'h7E; B = 8'hBF; #100;
A = 8'h7E; B = 8'hC0; #100;
A = 8'h7E; B = 8'hC1; #100;
A = 8'h7E; B = 8'hC2; #100;
A = 8'h7E; B = 8'hC3; #100;
A = 8'h7E; B = 8'hC4; #100;
A = 8'h7E; B = 8'hC5; #100;
A = 8'h7E; B = 8'hC6; #100;
A = 8'h7E; B = 8'hC7; #100;
A = 8'h7E; B = 8'hC8; #100;
A = 8'h7E; B = 8'hC9; #100;
A = 8'h7E; B = 8'hCA; #100;
A = 8'h7E; B = 8'hCB; #100;
A = 8'h7E; B = 8'hCC; #100;
A = 8'h7E; B = 8'hCD; #100;
A = 8'h7E; B = 8'hCE; #100;
A = 8'h7E; B = 8'hCF; #100;
A = 8'h7E; B = 8'hD0; #100;
A = 8'h7E; B = 8'hD1; #100;
A = 8'h7E; B = 8'hD2; #100;
A = 8'h7E; B = 8'hD3; #100;
A = 8'h7E; B = 8'hD4; #100;
A = 8'h7E; B = 8'hD5; #100;
A = 8'h7E; B = 8'hD6; #100;
A = 8'h7E; B = 8'hD7; #100;
A = 8'h7E; B = 8'hD8; #100;
A = 8'h7E; B = 8'hD9; #100;
A = 8'h7E; B = 8'hDA; #100;
A = 8'h7E; B = 8'hDB; #100;
A = 8'h7E; B = 8'hDC; #100;
A = 8'h7E; B = 8'hDD; #100;
A = 8'h7E; B = 8'hDE; #100;
A = 8'h7E; B = 8'hDF; #100;
A = 8'h7E; B = 8'hE0; #100;
A = 8'h7E; B = 8'hE1; #100;
A = 8'h7E; B = 8'hE2; #100;
A = 8'h7E; B = 8'hE3; #100;
A = 8'h7E; B = 8'hE4; #100;
A = 8'h7E; B = 8'hE5; #100;
A = 8'h7E; B = 8'hE6; #100;
A = 8'h7E; B = 8'hE7; #100;
A = 8'h7E; B = 8'hE8; #100;
A = 8'h7E; B = 8'hE9; #100;
A = 8'h7E; B = 8'hEA; #100;
A = 8'h7E; B = 8'hEB; #100;
A = 8'h7E; B = 8'hEC; #100;
A = 8'h7E; B = 8'hED; #100;
A = 8'h7E; B = 8'hEE; #100;
A = 8'h7E; B = 8'hEF; #100;
A = 8'h7E; B = 8'hF0; #100;
A = 8'h7E; B = 8'hF1; #100;
A = 8'h7E; B = 8'hF2; #100;
A = 8'h7E; B = 8'hF3; #100;
A = 8'h7E; B = 8'hF4; #100;
A = 8'h7E; B = 8'hF5; #100;
A = 8'h7E; B = 8'hF6; #100;
A = 8'h7E; B = 8'hF7; #100;
A = 8'h7E; B = 8'hF8; #100;
A = 8'h7E; B = 8'hF9; #100;
A = 8'h7E; B = 8'hFA; #100;
A = 8'h7E; B = 8'hFB; #100;
A = 8'h7E; B = 8'hFC; #100;
A = 8'h7E; B = 8'hFD; #100;
A = 8'h7E; B = 8'hFE; #100;
A = 8'h7E; B = 8'hFF; #100;
A = 8'h7F; B = 8'h0; #100;
A = 8'h7F; B = 8'h1; #100;
A = 8'h7F; B = 8'h2; #100;
A = 8'h7F; B = 8'h3; #100;
A = 8'h7F; B = 8'h4; #100;
A = 8'h7F; B = 8'h5; #100;
A = 8'h7F; B = 8'h6; #100;
A = 8'h7F; B = 8'h7; #100;
A = 8'h7F; B = 8'h8; #100;
A = 8'h7F; B = 8'h9; #100;
A = 8'h7F; B = 8'hA; #100;
A = 8'h7F; B = 8'hB; #100;
A = 8'h7F; B = 8'hC; #100;
A = 8'h7F; B = 8'hD; #100;
A = 8'h7F; B = 8'hE; #100;
A = 8'h7F; B = 8'hF; #100;
A = 8'h7F; B = 8'h10; #100;
A = 8'h7F; B = 8'h11; #100;
A = 8'h7F; B = 8'h12; #100;
A = 8'h7F; B = 8'h13; #100;
A = 8'h7F; B = 8'h14; #100;
A = 8'h7F; B = 8'h15; #100;
A = 8'h7F; B = 8'h16; #100;
A = 8'h7F; B = 8'h17; #100;
A = 8'h7F; B = 8'h18; #100;
A = 8'h7F; B = 8'h19; #100;
A = 8'h7F; B = 8'h1A; #100;
A = 8'h7F; B = 8'h1B; #100;
A = 8'h7F; B = 8'h1C; #100;
A = 8'h7F; B = 8'h1D; #100;
A = 8'h7F; B = 8'h1E; #100;
A = 8'h7F; B = 8'h1F; #100;
A = 8'h7F; B = 8'h20; #100;
A = 8'h7F; B = 8'h21; #100;
A = 8'h7F; B = 8'h22; #100;
A = 8'h7F; B = 8'h23; #100;
A = 8'h7F; B = 8'h24; #100;
A = 8'h7F; B = 8'h25; #100;
A = 8'h7F; B = 8'h26; #100;
A = 8'h7F; B = 8'h27; #100;
A = 8'h7F; B = 8'h28; #100;
A = 8'h7F; B = 8'h29; #100;
A = 8'h7F; B = 8'h2A; #100;
A = 8'h7F; B = 8'h2B; #100;
A = 8'h7F; B = 8'h2C; #100;
A = 8'h7F; B = 8'h2D; #100;
A = 8'h7F; B = 8'h2E; #100;
A = 8'h7F; B = 8'h2F; #100;
A = 8'h7F; B = 8'h30; #100;
A = 8'h7F; B = 8'h31; #100;
A = 8'h7F; B = 8'h32; #100;
A = 8'h7F; B = 8'h33; #100;
A = 8'h7F; B = 8'h34; #100;
A = 8'h7F; B = 8'h35; #100;
A = 8'h7F; B = 8'h36; #100;
A = 8'h7F; B = 8'h37; #100;
A = 8'h7F; B = 8'h38; #100;
A = 8'h7F; B = 8'h39; #100;
A = 8'h7F; B = 8'h3A; #100;
A = 8'h7F; B = 8'h3B; #100;
A = 8'h7F; B = 8'h3C; #100;
A = 8'h7F; B = 8'h3D; #100;
A = 8'h7F; B = 8'h3E; #100;
A = 8'h7F; B = 8'h3F; #100;
A = 8'h7F; B = 8'h40; #100;
A = 8'h7F; B = 8'h41; #100;
A = 8'h7F; B = 8'h42; #100;
A = 8'h7F; B = 8'h43; #100;
A = 8'h7F; B = 8'h44; #100;
A = 8'h7F; B = 8'h45; #100;
A = 8'h7F; B = 8'h46; #100;
A = 8'h7F; B = 8'h47; #100;
A = 8'h7F; B = 8'h48; #100;
A = 8'h7F; B = 8'h49; #100;
A = 8'h7F; B = 8'h4A; #100;
A = 8'h7F; B = 8'h4B; #100;
A = 8'h7F; B = 8'h4C; #100;
A = 8'h7F; B = 8'h4D; #100;
A = 8'h7F; B = 8'h4E; #100;
A = 8'h7F; B = 8'h4F; #100;
A = 8'h7F; B = 8'h50; #100;
A = 8'h7F; B = 8'h51; #100;
A = 8'h7F; B = 8'h52; #100;
A = 8'h7F; B = 8'h53; #100;
A = 8'h7F; B = 8'h54; #100;
A = 8'h7F; B = 8'h55; #100;
A = 8'h7F; B = 8'h56; #100;
A = 8'h7F; B = 8'h57; #100;
A = 8'h7F; B = 8'h58; #100;
A = 8'h7F; B = 8'h59; #100;
A = 8'h7F; B = 8'h5A; #100;
A = 8'h7F; B = 8'h5B; #100;
A = 8'h7F; B = 8'h5C; #100;
A = 8'h7F; B = 8'h5D; #100;
A = 8'h7F; B = 8'h5E; #100;
A = 8'h7F; B = 8'h5F; #100;
A = 8'h7F; B = 8'h60; #100;
A = 8'h7F; B = 8'h61; #100;
A = 8'h7F; B = 8'h62; #100;
A = 8'h7F; B = 8'h63; #100;
A = 8'h7F; B = 8'h64; #100;
A = 8'h7F; B = 8'h65; #100;
A = 8'h7F; B = 8'h66; #100;
A = 8'h7F; B = 8'h67; #100;
A = 8'h7F; B = 8'h68; #100;
A = 8'h7F; B = 8'h69; #100;
A = 8'h7F; B = 8'h6A; #100;
A = 8'h7F; B = 8'h6B; #100;
A = 8'h7F; B = 8'h6C; #100;
A = 8'h7F; B = 8'h6D; #100;
A = 8'h7F; B = 8'h6E; #100;
A = 8'h7F; B = 8'h6F; #100;
A = 8'h7F; B = 8'h70; #100;
A = 8'h7F; B = 8'h71; #100;
A = 8'h7F; B = 8'h72; #100;
A = 8'h7F; B = 8'h73; #100;
A = 8'h7F; B = 8'h74; #100;
A = 8'h7F; B = 8'h75; #100;
A = 8'h7F; B = 8'h76; #100;
A = 8'h7F; B = 8'h77; #100;
A = 8'h7F; B = 8'h78; #100;
A = 8'h7F; B = 8'h79; #100;
A = 8'h7F; B = 8'h7A; #100;
A = 8'h7F; B = 8'h7B; #100;
A = 8'h7F; B = 8'h7C; #100;
A = 8'h7F; B = 8'h7D; #100;
A = 8'h7F; B = 8'h7E; #100;
A = 8'h7F; B = 8'h7F; #100;
A = 8'h7F; B = 8'h80; #100;
A = 8'h7F; B = 8'h81; #100;
A = 8'h7F; B = 8'h82; #100;
A = 8'h7F; B = 8'h83; #100;
A = 8'h7F; B = 8'h84; #100;
A = 8'h7F; B = 8'h85; #100;
A = 8'h7F; B = 8'h86; #100;
A = 8'h7F; B = 8'h87; #100;
A = 8'h7F; B = 8'h88; #100;
A = 8'h7F; B = 8'h89; #100;
A = 8'h7F; B = 8'h8A; #100;
A = 8'h7F; B = 8'h8B; #100;
A = 8'h7F; B = 8'h8C; #100;
A = 8'h7F; B = 8'h8D; #100;
A = 8'h7F; B = 8'h8E; #100;
A = 8'h7F; B = 8'h8F; #100;
A = 8'h7F; B = 8'h90; #100;
A = 8'h7F; B = 8'h91; #100;
A = 8'h7F; B = 8'h92; #100;
A = 8'h7F; B = 8'h93; #100;
A = 8'h7F; B = 8'h94; #100;
A = 8'h7F; B = 8'h95; #100;
A = 8'h7F; B = 8'h96; #100;
A = 8'h7F; B = 8'h97; #100;
A = 8'h7F; B = 8'h98; #100;
A = 8'h7F; B = 8'h99; #100;
A = 8'h7F; B = 8'h9A; #100;
A = 8'h7F; B = 8'h9B; #100;
A = 8'h7F; B = 8'h9C; #100;
A = 8'h7F; B = 8'h9D; #100;
A = 8'h7F; B = 8'h9E; #100;
A = 8'h7F; B = 8'h9F; #100;
A = 8'h7F; B = 8'hA0; #100;
A = 8'h7F; B = 8'hA1; #100;
A = 8'h7F; B = 8'hA2; #100;
A = 8'h7F; B = 8'hA3; #100;
A = 8'h7F; B = 8'hA4; #100;
A = 8'h7F; B = 8'hA5; #100;
A = 8'h7F; B = 8'hA6; #100;
A = 8'h7F; B = 8'hA7; #100;
A = 8'h7F; B = 8'hA8; #100;
A = 8'h7F; B = 8'hA9; #100;
A = 8'h7F; B = 8'hAA; #100;
A = 8'h7F; B = 8'hAB; #100;
A = 8'h7F; B = 8'hAC; #100;
A = 8'h7F; B = 8'hAD; #100;
A = 8'h7F; B = 8'hAE; #100;
A = 8'h7F; B = 8'hAF; #100;
A = 8'h7F; B = 8'hB0; #100;
A = 8'h7F; B = 8'hB1; #100;
A = 8'h7F; B = 8'hB2; #100;
A = 8'h7F; B = 8'hB3; #100;
A = 8'h7F; B = 8'hB4; #100;
A = 8'h7F; B = 8'hB5; #100;
A = 8'h7F; B = 8'hB6; #100;
A = 8'h7F; B = 8'hB7; #100;
A = 8'h7F; B = 8'hB8; #100;
A = 8'h7F; B = 8'hB9; #100;
A = 8'h7F; B = 8'hBA; #100;
A = 8'h7F; B = 8'hBB; #100;
A = 8'h7F; B = 8'hBC; #100;
A = 8'h7F; B = 8'hBD; #100;
A = 8'h7F; B = 8'hBE; #100;
A = 8'h7F; B = 8'hBF; #100;
A = 8'h7F; B = 8'hC0; #100;
A = 8'h7F; B = 8'hC1; #100;
A = 8'h7F; B = 8'hC2; #100;
A = 8'h7F; B = 8'hC3; #100;
A = 8'h7F; B = 8'hC4; #100;
A = 8'h7F; B = 8'hC5; #100;
A = 8'h7F; B = 8'hC6; #100;
A = 8'h7F; B = 8'hC7; #100;
A = 8'h7F; B = 8'hC8; #100;
A = 8'h7F; B = 8'hC9; #100;
A = 8'h7F; B = 8'hCA; #100;
A = 8'h7F; B = 8'hCB; #100;
A = 8'h7F; B = 8'hCC; #100;
A = 8'h7F; B = 8'hCD; #100;
A = 8'h7F; B = 8'hCE; #100;
A = 8'h7F; B = 8'hCF; #100;
A = 8'h7F; B = 8'hD0; #100;
A = 8'h7F; B = 8'hD1; #100;
A = 8'h7F; B = 8'hD2; #100;
A = 8'h7F; B = 8'hD3; #100;
A = 8'h7F; B = 8'hD4; #100;
A = 8'h7F; B = 8'hD5; #100;
A = 8'h7F; B = 8'hD6; #100;
A = 8'h7F; B = 8'hD7; #100;
A = 8'h7F; B = 8'hD8; #100;
A = 8'h7F; B = 8'hD9; #100;
A = 8'h7F; B = 8'hDA; #100;
A = 8'h7F; B = 8'hDB; #100;
A = 8'h7F; B = 8'hDC; #100;
A = 8'h7F; B = 8'hDD; #100;
A = 8'h7F; B = 8'hDE; #100;
A = 8'h7F; B = 8'hDF; #100;
A = 8'h7F; B = 8'hE0; #100;
A = 8'h7F; B = 8'hE1; #100;
A = 8'h7F; B = 8'hE2; #100;
A = 8'h7F; B = 8'hE3; #100;
A = 8'h7F; B = 8'hE4; #100;
A = 8'h7F; B = 8'hE5; #100;
A = 8'h7F; B = 8'hE6; #100;
A = 8'h7F; B = 8'hE7; #100;
A = 8'h7F; B = 8'hE8; #100;
A = 8'h7F; B = 8'hE9; #100;
A = 8'h7F; B = 8'hEA; #100;
A = 8'h7F; B = 8'hEB; #100;
A = 8'h7F; B = 8'hEC; #100;
A = 8'h7F; B = 8'hED; #100;
A = 8'h7F; B = 8'hEE; #100;
A = 8'h7F; B = 8'hEF; #100;
A = 8'h7F; B = 8'hF0; #100;
A = 8'h7F; B = 8'hF1; #100;
A = 8'h7F; B = 8'hF2; #100;
A = 8'h7F; B = 8'hF3; #100;
A = 8'h7F; B = 8'hF4; #100;
A = 8'h7F; B = 8'hF5; #100;
A = 8'h7F; B = 8'hF6; #100;
A = 8'h7F; B = 8'hF7; #100;
A = 8'h7F; B = 8'hF8; #100;
A = 8'h7F; B = 8'hF9; #100;
A = 8'h7F; B = 8'hFA; #100;
A = 8'h7F; B = 8'hFB; #100;
A = 8'h7F; B = 8'hFC; #100;
A = 8'h7F; B = 8'hFD; #100;
A = 8'h7F; B = 8'hFE; #100;
A = 8'h7F; B = 8'hFF; #100;
A = 8'h80; B = 8'h0; #100;
A = 8'h80; B = 8'h1; #100;
A = 8'h80; B = 8'h2; #100;
A = 8'h80; B = 8'h3; #100;
A = 8'h80; B = 8'h4; #100;
A = 8'h80; B = 8'h5; #100;
A = 8'h80; B = 8'h6; #100;
A = 8'h80; B = 8'h7; #100;
A = 8'h80; B = 8'h8; #100;
A = 8'h80; B = 8'h9; #100;
A = 8'h80; B = 8'hA; #100;
A = 8'h80; B = 8'hB; #100;
A = 8'h80; B = 8'hC; #100;
A = 8'h80; B = 8'hD; #100;
A = 8'h80; B = 8'hE; #100;
A = 8'h80; B = 8'hF; #100;
A = 8'h80; B = 8'h10; #100;
A = 8'h80; B = 8'h11; #100;
A = 8'h80; B = 8'h12; #100;
A = 8'h80; B = 8'h13; #100;
A = 8'h80; B = 8'h14; #100;
A = 8'h80; B = 8'h15; #100;
A = 8'h80; B = 8'h16; #100;
A = 8'h80; B = 8'h17; #100;
A = 8'h80; B = 8'h18; #100;
A = 8'h80; B = 8'h19; #100;
A = 8'h80; B = 8'h1A; #100;
A = 8'h80; B = 8'h1B; #100;
A = 8'h80; B = 8'h1C; #100;
A = 8'h80; B = 8'h1D; #100;
A = 8'h80; B = 8'h1E; #100;
A = 8'h80; B = 8'h1F; #100;
A = 8'h80; B = 8'h20; #100;
A = 8'h80; B = 8'h21; #100;
A = 8'h80; B = 8'h22; #100;
A = 8'h80; B = 8'h23; #100;
A = 8'h80; B = 8'h24; #100;
A = 8'h80; B = 8'h25; #100;
A = 8'h80; B = 8'h26; #100;
A = 8'h80; B = 8'h27; #100;
A = 8'h80; B = 8'h28; #100;
A = 8'h80; B = 8'h29; #100;
A = 8'h80; B = 8'h2A; #100;
A = 8'h80; B = 8'h2B; #100;
A = 8'h80; B = 8'h2C; #100;
A = 8'h80; B = 8'h2D; #100;
A = 8'h80; B = 8'h2E; #100;
A = 8'h80; B = 8'h2F; #100;
A = 8'h80; B = 8'h30; #100;
A = 8'h80; B = 8'h31; #100;
A = 8'h80; B = 8'h32; #100;
A = 8'h80; B = 8'h33; #100;
A = 8'h80; B = 8'h34; #100;
A = 8'h80; B = 8'h35; #100;
A = 8'h80; B = 8'h36; #100;
A = 8'h80; B = 8'h37; #100;
A = 8'h80; B = 8'h38; #100;
A = 8'h80; B = 8'h39; #100;
A = 8'h80; B = 8'h3A; #100;
A = 8'h80; B = 8'h3B; #100;
A = 8'h80; B = 8'h3C; #100;
A = 8'h80; B = 8'h3D; #100;
A = 8'h80; B = 8'h3E; #100;
A = 8'h80; B = 8'h3F; #100;
A = 8'h80; B = 8'h40; #100;
A = 8'h80; B = 8'h41; #100;
A = 8'h80; B = 8'h42; #100;
A = 8'h80; B = 8'h43; #100;
A = 8'h80; B = 8'h44; #100;
A = 8'h80; B = 8'h45; #100;
A = 8'h80; B = 8'h46; #100;
A = 8'h80; B = 8'h47; #100;
A = 8'h80; B = 8'h48; #100;
A = 8'h80; B = 8'h49; #100;
A = 8'h80; B = 8'h4A; #100;
A = 8'h80; B = 8'h4B; #100;
A = 8'h80; B = 8'h4C; #100;
A = 8'h80; B = 8'h4D; #100;
A = 8'h80; B = 8'h4E; #100;
A = 8'h80; B = 8'h4F; #100;
A = 8'h80; B = 8'h50; #100;
A = 8'h80; B = 8'h51; #100;
A = 8'h80; B = 8'h52; #100;
A = 8'h80; B = 8'h53; #100;
A = 8'h80; B = 8'h54; #100;
A = 8'h80; B = 8'h55; #100;
A = 8'h80; B = 8'h56; #100;
A = 8'h80; B = 8'h57; #100;
A = 8'h80; B = 8'h58; #100;
A = 8'h80; B = 8'h59; #100;
A = 8'h80; B = 8'h5A; #100;
A = 8'h80; B = 8'h5B; #100;
A = 8'h80; B = 8'h5C; #100;
A = 8'h80; B = 8'h5D; #100;
A = 8'h80; B = 8'h5E; #100;
A = 8'h80; B = 8'h5F; #100;
A = 8'h80; B = 8'h60; #100;
A = 8'h80; B = 8'h61; #100;
A = 8'h80; B = 8'h62; #100;
A = 8'h80; B = 8'h63; #100;
A = 8'h80; B = 8'h64; #100;
A = 8'h80; B = 8'h65; #100;
A = 8'h80; B = 8'h66; #100;
A = 8'h80; B = 8'h67; #100;
A = 8'h80; B = 8'h68; #100;
A = 8'h80; B = 8'h69; #100;
A = 8'h80; B = 8'h6A; #100;
A = 8'h80; B = 8'h6B; #100;
A = 8'h80; B = 8'h6C; #100;
A = 8'h80; B = 8'h6D; #100;
A = 8'h80; B = 8'h6E; #100;
A = 8'h80; B = 8'h6F; #100;
A = 8'h80; B = 8'h70; #100;
A = 8'h80; B = 8'h71; #100;
A = 8'h80; B = 8'h72; #100;
A = 8'h80; B = 8'h73; #100;
A = 8'h80; B = 8'h74; #100;
A = 8'h80; B = 8'h75; #100;
A = 8'h80; B = 8'h76; #100;
A = 8'h80; B = 8'h77; #100;
A = 8'h80; B = 8'h78; #100;
A = 8'h80; B = 8'h79; #100;
A = 8'h80; B = 8'h7A; #100;
A = 8'h80; B = 8'h7B; #100;
A = 8'h80; B = 8'h7C; #100;
A = 8'h80; B = 8'h7D; #100;
A = 8'h80; B = 8'h7E; #100;
A = 8'h80; B = 8'h7F; #100;
A = 8'h80; B = 8'h80; #100;
A = 8'h80; B = 8'h81; #100;
A = 8'h80; B = 8'h82; #100;
A = 8'h80; B = 8'h83; #100;
A = 8'h80; B = 8'h84; #100;
A = 8'h80; B = 8'h85; #100;
A = 8'h80; B = 8'h86; #100;
A = 8'h80; B = 8'h87; #100;
A = 8'h80; B = 8'h88; #100;
A = 8'h80; B = 8'h89; #100;
A = 8'h80; B = 8'h8A; #100;
A = 8'h80; B = 8'h8B; #100;
A = 8'h80; B = 8'h8C; #100;
A = 8'h80; B = 8'h8D; #100;
A = 8'h80; B = 8'h8E; #100;
A = 8'h80; B = 8'h8F; #100;
A = 8'h80; B = 8'h90; #100;
A = 8'h80; B = 8'h91; #100;
A = 8'h80; B = 8'h92; #100;
A = 8'h80; B = 8'h93; #100;
A = 8'h80; B = 8'h94; #100;
A = 8'h80; B = 8'h95; #100;
A = 8'h80; B = 8'h96; #100;
A = 8'h80; B = 8'h97; #100;
A = 8'h80; B = 8'h98; #100;
A = 8'h80; B = 8'h99; #100;
A = 8'h80; B = 8'h9A; #100;
A = 8'h80; B = 8'h9B; #100;
A = 8'h80; B = 8'h9C; #100;
A = 8'h80; B = 8'h9D; #100;
A = 8'h80; B = 8'h9E; #100;
A = 8'h80; B = 8'h9F; #100;
A = 8'h80; B = 8'hA0; #100;
A = 8'h80; B = 8'hA1; #100;
A = 8'h80; B = 8'hA2; #100;
A = 8'h80; B = 8'hA3; #100;
A = 8'h80; B = 8'hA4; #100;
A = 8'h80; B = 8'hA5; #100;
A = 8'h80; B = 8'hA6; #100;
A = 8'h80; B = 8'hA7; #100;
A = 8'h80; B = 8'hA8; #100;
A = 8'h80; B = 8'hA9; #100;
A = 8'h80; B = 8'hAA; #100;
A = 8'h80; B = 8'hAB; #100;
A = 8'h80; B = 8'hAC; #100;
A = 8'h80; B = 8'hAD; #100;
A = 8'h80; B = 8'hAE; #100;
A = 8'h80; B = 8'hAF; #100;
A = 8'h80; B = 8'hB0; #100;
A = 8'h80; B = 8'hB1; #100;
A = 8'h80; B = 8'hB2; #100;
A = 8'h80; B = 8'hB3; #100;
A = 8'h80; B = 8'hB4; #100;
A = 8'h80; B = 8'hB5; #100;
A = 8'h80; B = 8'hB6; #100;
A = 8'h80; B = 8'hB7; #100;
A = 8'h80; B = 8'hB8; #100;
A = 8'h80; B = 8'hB9; #100;
A = 8'h80; B = 8'hBA; #100;
A = 8'h80; B = 8'hBB; #100;
A = 8'h80; B = 8'hBC; #100;
A = 8'h80; B = 8'hBD; #100;
A = 8'h80; B = 8'hBE; #100;
A = 8'h80; B = 8'hBF; #100;
A = 8'h80; B = 8'hC0; #100;
A = 8'h80; B = 8'hC1; #100;
A = 8'h80; B = 8'hC2; #100;
A = 8'h80; B = 8'hC3; #100;
A = 8'h80; B = 8'hC4; #100;
A = 8'h80; B = 8'hC5; #100;
A = 8'h80; B = 8'hC6; #100;
A = 8'h80; B = 8'hC7; #100;
A = 8'h80; B = 8'hC8; #100;
A = 8'h80; B = 8'hC9; #100;
A = 8'h80; B = 8'hCA; #100;
A = 8'h80; B = 8'hCB; #100;
A = 8'h80; B = 8'hCC; #100;
A = 8'h80; B = 8'hCD; #100;
A = 8'h80; B = 8'hCE; #100;
A = 8'h80; B = 8'hCF; #100;
A = 8'h80; B = 8'hD0; #100;
A = 8'h80; B = 8'hD1; #100;
A = 8'h80; B = 8'hD2; #100;
A = 8'h80; B = 8'hD3; #100;
A = 8'h80; B = 8'hD4; #100;
A = 8'h80; B = 8'hD5; #100;
A = 8'h80; B = 8'hD6; #100;
A = 8'h80; B = 8'hD7; #100;
A = 8'h80; B = 8'hD8; #100;
A = 8'h80; B = 8'hD9; #100;
A = 8'h80; B = 8'hDA; #100;
A = 8'h80; B = 8'hDB; #100;
A = 8'h80; B = 8'hDC; #100;
A = 8'h80; B = 8'hDD; #100;
A = 8'h80; B = 8'hDE; #100;
A = 8'h80; B = 8'hDF; #100;
A = 8'h80; B = 8'hE0; #100;
A = 8'h80; B = 8'hE1; #100;
A = 8'h80; B = 8'hE2; #100;
A = 8'h80; B = 8'hE3; #100;
A = 8'h80; B = 8'hE4; #100;
A = 8'h80; B = 8'hE5; #100;
A = 8'h80; B = 8'hE6; #100;
A = 8'h80; B = 8'hE7; #100;
A = 8'h80; B = 8'hE8; #100;
A = 8'h80; B = 8'hE9; #100;
A = 8'h80; B = 8'hEA; #100;
A = 8'h80; B = 8'hEB; #100;
A = 8'h80; B = 8'hEC; #100;
A = 8'h80; B = 8'hED; #100;
A = 8'h80; B = 8'hEE; #100;
A = 8'h80; B = 8'hEF; #100;
A = 8'h80; B = 8'hF0; #100;
A = 8'h80; B = 8'hF1; #100;
A = 8'h80; B = 8'hF2; #100;
A = 8'h80; B = 8'hF3; #100;
A = 8'h80; B = 8'hF4; #100;
A = 8'h80; B = 8'hF5; #100;
A = 8'h80; B = 8'hF6; #100;
A = 8'h80; B = 8'hF7; #100;
A = 8'h80; B = 8'hF8; #100;
A = 8'h80; B = 8'hF9; #100;
A = 8'h80; B = 8'hFA; #100;
A = 8'h80; B = 8'hFB; #100;
A = 8'h80; B = 8'hFC; #100;
A = 8'h80; B = 8'hFD; #100;
A = 8'h80; B = 8'hFE; #100;
A = 8'h80; B = 8'hFF; #100;
A = 8'h81; B = 8'h0; #100;
A = 8'h81; B = 8'h1; #100;
A = 8'h81; B = 8'h2; #100;
A = 8'h81; B = 8'h3; #100;
A = 8'h81; B = 8'h4; #100;
A = 8'h81; B = 8'h5; #100;
A = 8'h81; B = 8'h6; #100;
A = 8'h81; B = 8'h7; #100;
A = 8'h81; B = 8'h8; #100;
A = 8'h81; B = 8'h9; #100;
A = 8'h81; B = 8'hA; #100;
A = 8'h81; B = 8'hB; #100;
A = 8'h81; B = 8'hC; #100;
A = 8'h81; B = 8'hD; #100;
A = 8'h81; B = 8'hE; #100;
A = 8'h81; B = 8'hF; #100;
A = 8'h81; B = 8'h10; #100;
A = 8'h81; B = 8'h11; #100;
A = 8'h81; B = 8'h12; #100;
A = 8'h81; B = 8'h13; #100;
A = 8'h81; B = 8'h14; #100;
A = 8'h81; B = 8'h15; #100;
A = 8'h81; B = 8'h16; #100;
A = 8'h81; B = 8'h17; #100;
A = 8'h81; B = 8'h18; #100;
A = 8'h81; B = 8'h19; #100;
A = 8'h81; B = 8'h1A; #100;
A = 8'h81; B = 8'h1B; #100;
A = 8'h81; B = 8'h1C; #100;
A = 8'h81; B = 8'h1D; #100;
A = 8'h81; B = 8'h1E; #100;
A = 8'h81; B = 8'h1F; #100;
A = 8'h81; B = 8'h20; #100;
A = 8'h81; B = 8'h21; #100;
A = 8'h81; B = 8'h22; #100;
A = 8'h81; B = 8'h23; #100;
A = 8'h81; B = 8'h24; #100;
A = 8'h81; B = 8'h25; #100;
A = 8'h81; B = 8'h26; #100;
A = 8'h81; B = 8'h27; #100;
A = 8'h81; B = 8'h28; #100;
A = 8'h81; B = 8'h29; #100;
A = 8'h81; B = 8'h2A; #100;
A = 8'h81; B = 8'h2B; #100;
A = 8'h81; B = 8'h2C; #100;
A = 8'h81; B = 8'h2D; #100;
A = 8'h81; B = 8'h2E; #100;
A = 8'h81; B = 8'h2F; #100;
A = 8'h81; B = 8'h30; #100;
A = 8'h81; B = 8'h31; #100;
A = 8'h81; B = 8'h32; #100;
A = 8'h81; B = 8'h33; #100;
A = 8'h81; B = 8'h34; #100;
A = 8'h81; B = 8'h35; #100;
A = 8'h81; B = 8'h36; #100;
A = 8'h81; B = 8'h37; #100;
A = 8'h81; B = 8'h38; #100;
A = 8'h81; B = 8'h39; #100;
A = 8'h81; B = 8'h3A; #100;
A = 8'h81; B = 8'h3B; #100;
A = 8'h81; B = 8'h3C; #100;
A = 8'h81; B = 8'h3D; #100;
A = 8'h81; B = 8'h3E; #100;
A = 8'h81; B = 8'h3F; #100;
A = 8'h81; B = 8'h40; #100;
A = 8'h81; B = 8'h41; #100;
A = 8'h81; B = 8'h42; #100;
A = 8'h81; B = 8'h43; #100;
A = 8'h81; B = 8'h44; #100;
A = 8'h81; B = 8'h45; #100;
A = 8'h81; B = 8'h46; #100;
A = 8'h81; B = 8'h47; #100;
A = 8'h81; B = 8'h48; #100;
A = 8'h81; B = 8'h49; #100;
A = 8'h81; B = 8'h4A; #100;
A = 8'h81; B = 8'h4B; #100;
A = 8'h81; B = 8'h4C; #100;
A = 8'h81; B = 8'h4D; #100;
A = 8'h81; B = 8'h4E; #100;
A = 8'h81; B = 8'h4F; #100;
A = 8'h81; B = 8'h50; #100;
A = 8'h81; B = 8'h51; #100;
A = 8'h81; B = 8'h52; #100;
A = 8'h81; B = 8'h53; #100;
A = 8'h81; B = 8'h54; #100;
A = 8'h81; B = 8'h55; #100;
A = 8'h81; B = 8'h56; #100;
A = 8'h81; B = 8'h57; #100;
A = 8'h81; B = 8'h58; #100;
A = 8'h81; B = 8'h59; #100;
A = 8'h81; B = 8'h5A; #100;
A = 8'h81; B = 8'h5B; #100;
A = 8'h81; B = 8'h5C; #100;
A = 8'h81; B = 8'h5D; #100;
A = 8'h81; B = 8'h5E; #100;
A = 8'h81; B = 8'h5F; #100;
A = 8'h81; B = 8'h60; #100;
A = 8'h81; B = 8'h61; #100;
A = 8'h81; B = 8'h62; #100;
A = 8'h81; B = 8'h63; #100;
A = 8'h81; B = 8'h64; #100;
A = 8'h81; B = 8'h65; #100;
A = 8'h81; B = 8'h66; #100;
A = 8'h81; B = 8'h67; #100;
A = 8'h81; B = 8'h68; #100;
A = 8'h81; B = 8'h69; #100;
A = 8'h81; B = 8'h6A; #100;
A = 8'h81; B = 8'h6B; #100;
A = 8'h81; B = 8'h6C; #100;
A = 8'h81; B = 8'h6D; #100;
A = 8'h81; B = 8'h6E; #100;
A = 8'h81; B = 8'h6F; #100;
A = 8'h81; B = 8'h70; #100;
A = 8'h81; B = 8'h71; #100;
A = 8'h81; B = 8'h72; #100;
A = 8'h81; B = 8'h73; #100;
A = 8'h81; B = 8'h74; #100;
A = 8'h81; B = 8'h75; #100;
A = 8'h81; B = 8'h76; #100;
A = 8'h81; B = 8'h77; #100;
A = 8'h81; B = 8'h78; #100;
A = 8'h81; B = 8'h79; #100;
A = 8'h81; B = 8'h7A; #100;
A = 8'h81; B = 8'h7B; #100;
A = 8'h81; B = 8'h7C; #100;
A = 8'h81; B = 8'h7D; #100;
A = 8'h81; B = 8'h7E; #100;
A = 8'h81; B = 8'h7F; #100;
A = 8'h81; B = 8'h80; #100;
A = 8'h81; B = 8'h81; #100;
A = 8'h81; B = 8'h82; #100;
A = 8'h81; B = 8'h83; #100;
A = 8'h81; B = 8'h84; #100;
A = 8'h81; B = 8'h85; #100;
A = 8'h81; B = 8'h86; #100;
A = 8'h81; B = 8'h87; #100;
A = 8'h81; B = 8'h88; #100;
A = 8'h81; B = 8'h89; #100;
A = 8'h81; B = 8'h8A; #100;
A = 8'h81; B = 8'h8B; #100;
A = 8'h81; B = 8'h8C; #100;
A = 8'h81; B = 8'h8D; #100;
A = 8'h81; B = 8'h8E; #100;
A = 8'h81; B = 8'h8F; #100;
A = 8'h81; B = 8'h90; #100;
A = 8'h81; B = 8'h91; #100;
A = 8'h81; B = 8'h92; #100;
A = 8'h81; B = 8'h93; #100;
A = 8'h81; B = 8'h94; #100;
A = 8'h81; B = 8'h95; #100;
A = 8'h81; B = 8'h96; #100;
A = 8'h81; B = 8'h97; #100;
A = 8'h81; B = 8'h98; #100;
A = 8'h81; B = 8'h99; #100;
A = 8'h81; B = 8'h9A; #100;
A = 8'h81; B = 8'h9B; #100;
A = 8'h81; B = 8'h9C; #100;
A = 8'h81; B = 8'h9D; #100;
A = 8'h81; B = 8'h9E; #100;
A = 8'h81; B = 8'h9F; #100;
A = 8'h81; B = 8'hA0; #100;
A = 8'h81; B = 8'hA1; #100;
A = 8'h81; B = 8'hA2; #100;
A = 8'h81; B = 8'hA3; #100;
A = 8'h81; B = 8'hA4; #100;
A = 8'h81; B = 8'hA5; #100;
A = 8'h81; B = 8'hA6; #100;
A = 8'h81; B = 8'hA7; #100;
A = 8'h81; B = 8'hA8; #100;
A = 8'h81; B = 8'hA9; #100;
A = 8'h81; B = 8'hAA; #100;
A = 8'h81; B = 8'hAB; #100;
A = 8'h81; B = 8'hAC; #100;
A = 8'h81; B = 8'hAD; #100;
A = 8'h81; B = 8'hAE; #100;
A = 8'h81; B = 8'hAF; #100;
A = 8'h81; B = 8'hB0; #100;
A = 8'h81; B = 8'hB1; #100;
A = 8'h81; B = 8'hB2; #100;
A = 8'h81; B = 8'hB3; #100;
A = 8'h81; B = 8'hB4; #100;
A = 8'h81; B = 8'hB5; #100;
A = 8'h81; B = 8'hB6; #100;
A = 8'h81; B = 8'hB7; #100;
A = 8'h81; B = 8'hB8; #100;
A = 8'h81; B = 8'hB9; #100;
A = 8'h81; B = 8'hBA; #100;
A = 8'h81; B = 8'hBB; #100;
A = 8'h81; B = 8'hBC; #100;
A = 8'h81; B = 8'hBD; #100;
A = 8'h81; B = 8'hBE; #100;
A = 8'h81; B = 8'hBF; #100;
A = 8'h81; B = 8'hC0; #100;
A = 8'h81; B = 8'hC1; #100;
A = 8'h81; B = 8'hC2; #100;
A = 8'h81; B = 8'hC3; #100;
A = 8'h81; B = 8'hC4; #100;
A = 8'h81; B = 8'hC5; #100;
A = 8'h81; B = 8'hC6; #100;
A = 8'h81; B = 8'hC7; #100;
A = 8'h81; B = 8'hC8; #100;
A = 8'h81; B = 8'hC9; #100;
A = 8'h81; B = 8'hCA; #100;
A = 8'h81; B = 8'hCB; #100;
A = 8'h81; B = 8'hCC; #100;
A = 8'h81; B = 8'hCD; #100;
A = 8'h81; B = 8'hCE; #100;
A = 8'h81; B = 8'hCF; #100;
A = 8'h81; B = 8'hD0; #100;
A = 8'h81; B = 8'hD1; #100;
A = 8'h81; B = 8'hD2; #100;
A = 8'h81; B = 8'hD3; #100;
A = 8'h81; B = 8'hD4; #100;
A = 8'h81; B = 8'hD5; #100;
A = 8'h81; B = 8'hD6; #100;
A = 8'h81; B = 8'hD7; #100;
A = 8'h81; B = 8'hD8; #100;
A = 8'h81; B = 8'hD9; #100;
A = 8'h81; B = 8'hDA; #100;
A = 8'h81; B = 8'hDB; #100;
A = 8'h81; B = 8'hDC; #100;
A = 8'h81; B = 8'hDD; #100;
A = 8'h81; B = 8'hDE; #100;
A = 8'h81; B = 8'hDF; #100;
A = 8'h81; B = 8'hE0; #100;
A = 8'h81; B = 8'hE1; #100;
A = 8'h81; B = 8'hE2; #100;
A = 8'h81; B = 8'hE3; #100;
A = 8'h81; B = 8'hE4; #100;
A = 8'h81; B = 8'hE5; #100;
A = 8'h81; B = 8'hE6; #100;
A = 8'h81; B = 8'hE7; #100;
A = 8'h81; B = 8'hE8; #100;
A = 8'h81; B = 8'hE9; #100;
A = 8'h81; B = 8'hEA; #100;
A = 8'h81; B = 8'hEB; #100;
A = 8'h81; B = 8'hEC; #100;
A = 8'h81; B = 8'hED; #100;
A = 8'h81; B = 8'hEE; #100;
A = 8'h81; B = 8'hEF; #100;
A = 8'h81; B = 8'hF0; #100;
A = 8'h81; B = 8'hF1; #100;
A = 8'h81; B = 8'hF2; #100;
A = 8'h81; B = 8'hF3; #100;
A = 8'h81; B = 8'hF4; #100;
A = 8'h81; B = 8'hF5; #100;
A = 8'h81; B = 8'hF6; #100;
A = 8'h81; B = 8'hF7; #100;
A = 8'h81; B = 8'hF8; #100;
A = 8'h81; B = 8'hF9; #100;
A = 8'h81; B = 8'hFA; #100;
A = 8'h81; B = 8'hFB; #100;
A = 8'h81; B = 8'hFC; #100;
A = 8'h81; B = 8'hFD; #100;
A = 8'h81; B = 8'hFE; #100;
A = 8'h81; B = 8'hFF; #100;
A = 8'h82; B = 8'h0; #100;
A = 8'h82; B = 8'h1; #100;
A = 8'h82; B = 8'h2; #100;
A = 8'h82; B = 8'h3; #100;
A = 8'h82; B = 8'h4; #100;
A = 8'h82; B = 8'h5; #100;
A = 8'h82; B = 8'h6; #100;
A = 8'h82; B = 8'h7; #100;
A = 8'h82; B = 8'h8; #100;
A = 8'h82; B = 8'h9; #100;
A = 8'h82; B = 8'hA; #100;
A = 8'h82; B = 8'hB; #100;
A = 8'h82; B = 8'hC; #100;
A = 8'h82; B = 8'hD; #100;
A = 8'h82; B = 8'hE; #100;
A = 8'h82; B = 8'hF; #100;
A = 8'h82; B = 8'h10; #100;
A = 8'h82; B = 8'h11; #100;
A = 8'h82; B = 8'h12; #100;
A = 8'h82; B = 8'h13; #100;
A = 8'h82; B = 8'h14; #100;
A = 8'h82; B = 8'h15; #100;
A = 8'h82; B = 8'h16; #100;
A = 8'h82; B = 8'h17; #100;
A = 8'h82; B = 8'h18; #100;
A = 8'h82; B = 8'h19; #100;
A = 8'h82; B = 8'h1A; #100;
A = 8'h82; B = 8'h1B; #100;
A = 8'h82; B = 8'h1C; #100;
A = 8'h82; B = 8'h1D; #100;
A = 8'h82; B = 8'h1E; #100;
A = 8'h82; B = 8'h1F; #100;
A = 8'h82; B = 8'h20; #100;
A = 8'h82; B = 8'h21; #100;
A = 8'h82; B = 8'h22; #100;
A = 8'h82; B = 8'h23; #100;
A = 8'h82; B = 8'h24; #100;
A = 8'h82; B = 8'h25; #100;
A = 8'h82; B = 8'h26; #100;
A = 8'h82; B = 8'h27; #100;
A = 8'h82; B = 8'h28; #100;
A = 8'h82; B = 8'h29; #100;
A = 8'h82; B = 8'h2A; #100;
A = 8'h82; B = 8'h2B; #100;
A = 8'h82; B = 8'h2C; #100;
A = 8'h82; B = 8'h2D; #100;
A = 8'h82; B = 8'h2E; #100;
A = 8'h82; B = 8'h2F; #100;
A = 8'h82; B = 8'h30; #100;
A = 8'h82; B = 8'h31; #100;
A = 8'h82; B = 8'h32; #100;
A = 8'h82; B = 8'h33; #100;
A = 8'h82; B = 8'h34; #100;
A = 8'h82; B = 8'h35; #100;
A = 8'h82; B = 8'h36; #100;
A = 8'h82; B = 8'h37; #100;
A = 8'h82; B = 8'h38; #100;
A = 8'h82; B = 8'h39; #100;
A = 8'h82; B = 8'h3A; #100;
A = 8'h82; B = 8'h3B; #100;
A = 8'h82; B = 8'h3C; #100;
A = 8'h82; B = 8'h3D; #100;
A = 8'h82; B = 8'h3E; #100;
A = 8'h82; B = 8'h3F; #100;
A = 8'h82; B = 8'h40; #100;
A = 8'h82; B = 8'h41; #100;
A = 8'h82; B = 8'h42; #100;
A = 8'h82; B = 8'h43; #100;
A = 8'h82; B = 8'h44; #100;
A = 8'h82; B = 8'h45; #100;
A = 8'h82; B = 8'h46; #100;
A = 8'h82; B = 8'h47; #100;
A = 8'h82; B = 8'h48; #100;
A = 8'h82; B = 8'h49; #100;
A = 8'h82; B = 8'h4A; #100;
A = 8'h82; B = 8'h4B; #100;
A = 8'h82; B = 8'h4C; #100;
A = 8'h82; B = 8'h4D; #100;
A = 8'h82; B = 8'h4E; #100;
A = 8'h82; B = 8'h4F; #100;
A = 8'h82; B = 8'h50; #100;
A = 8'h82; B = 8'h51; #100;
A = 8'h82; B = 8'h52; #100;
A = 8'h82; B = 8'h53; #100;
A = 8'h82; B = 8'h54; #100;
A = 8'h82; B = 8'h55; #100;
A = 8'h82; B = 8'h56; #100;
A = 8'h82; B = 8'h57; #100;
A = 8'h82; B = 8'h58; #100;
A = 8'h82; B = 8'h59; #100;
A = 8'h82; B = 8'h5A; #100;
A = 8'h82; B = 8'h5B; #100;
A = 8'h82; B = 8'h5C; #100;
A = 8'h82; B = 8'h5D; #100;
A = 8'h82; B = 8'h5E; #100;
A = 8'h82; B = 8'h5F; #100;
A = 8'h82; B = 8'h60; #100;
A = 8'h82; B = 8'h61; #100;
A = 8'h82; B = 8'h62; #100;
A = 8'h82; B = 8'h63; #100;
A = 8'h82; B = 8'h64; #100;
A = 8'h82; B = 8'h65; #100;
A = 8'h82; B = 8'h66; #100;
A = 8'h82; B = 8'h67; #100;
A = 8'h82; B = 8'h68; #100;
A = 8'h82; B = 8'h69; #100;
A = 8'h82; B = 8'h6A; #100;
A = 8'h82; B = 8'h6B; #100;
A = 8'h82; B = 8'h6C; #100;
A = 8'h82; B = 8'h6D; #100;
A = 8'h82; B = 8'h6E; #100;
A = 8'h82; B = 8'h6F; #100;
A = 8'h82; B = 8'h70; #100;
A = 8'h82; B = 8'h71; #100;
A = 8'h82; B = 8'h72; #100;
A = 8'h82; B = 8'h73; #100;
A = 8'h82; B = 8'h74; #100;
A = 8'h82; B = 8'h75; #100;
A = 8'h82; B = 8'h76; #100;
A = 8'h82; B = 8'h77; #100;
A = 8'h82; B = 8'h78; #100;
A = 8'h82; B = 8'h79; #100;
A = 8'h82; B = 8'h7A; #100;
A = 8'h82; B = 8'h7B; #100;
A = 8'h82; B = 8'h7C; #100;
A = 8'h82; B = 8'h7D; #100;
A = 8'h82; B = 8'h7E; #100;
A = 8'h82; B = 8'h7F; #100;
A = 8'h82; B = 8'h80; #100;
A = 8'h82; B = 8'h81; #100;
A = 8'h82; B = 8'h82; #100;
A = 8'h82; B = 8'h83; #100;
A = 8'h82; B = 8'h84; #100;
A = 8'h82; B = 8'h85; #100;
A = 8'h82; B = 8'h86; #100;
A = 8'h82; B = 8'h87; #100;
A = 8'h82; B = 8'h88; #100;
A = 8'h82; B = 8'h89; #100;
A = 8'h82; B = 8'h8A; #100;
A = 8'h82; B = 8'h8B; #100;
A = 8'h82; B = 8'h8C; #100;
A = 8'h82; B = 8'h8D; #100;
A = 8'h82; B = 8'h8E; #100;
A = 8'h82; B = 8'h8F; #100;
A = 8'h82; B = 8'h90; #100;
A = 8'h82; B = 8'h91; #100;
A = 8'h82; B = 8'h92; #100;
A = 8'h82; B = 8'h93; #100;
A = 8'h82; B = 8'h94; #100;
A = 8'h82; B = 8'h95; #100;
A = 8'h82; B = 8'h96; #100;
A = 8'h82; B = 8'h97; #100;
A = 8'h82; B = 8'h98; #100;
A = 8'h82; B = 8'h99; #100;
A = 8'h82; B = 8'h9A; #100;
A = 8'h82; B = 8'h9B; #100;
A = 8'h82; B = 8'h9C; #100;
A = 8'h82; B = 8'h9D; #100;
A = 8'h82; B = 8'h9E; #100;
A = 8'h82; B = 8'h9F; #100;
A = 8'h82; B = 8'hA0; #100;
A = 8'h82; B = 8'hA1; #100;
A = 8'h82; B = 8'hA2; #100;
A = 8'h82; B = 8'hA3; #100;
A = 8'h82; B = 8'hA4; #100;
A = 8'h82; B = 8'hA5; #100;
A = 8'h82; B = 8'hA6; #100;
A = 8'h82; B = 8'hA7; #100;
A = 8'h82; B = 8'hA8; #100;
A = 8'h82; B = 8'hA9; #100;
A = 8'h82; B = 8'hAA; #100;
A = 8'h82; B = 8'hAB; #100;
A = 8'h82; B = 8'hAC; #100;
A = 8'h82; B = 8'hAD; #100;
A = 8'h82; B = 8'hAE; #100;
A = 8'h82; B = 8'hAF; #100;
A = 8'h82; B = 8'hB0; #100;
A = 8'h82; B = 8'hB1; #100;
A = 8'h82; B = 8'hB2; #100;
A = 8'h82; B = 8'hB3; #100;
A = 8'h82; B = 8'hB4; #100;
A = 8'h82; B = 8'hB5; #100;
A = 8'h82; B = 8'hB6; #100;
A = 8'h82; B = 8'hB7; #100;
A = 8'h82; B = 8'hB8; #100;
A = 8'h82; B = 8'hB9; #100;
A = 8'h82; B = 8'hBA; #100;
A = 8'h82; B = 8'hBB; #100;
A = 8'h82; B = 8'hBC; #100;
A = 8'h82; B = 8'hBD; #100;
A = 8'h82; B = 8'hBE; #100;
A = 8'h82; B = 8'hBF; #100;
A = 8'h82; B = 8'hC0; #100;
A = 8'h82; B = 8'hC1; #100;
A = 8'h82; B = 8'hC2; #100;
A = 8'h82; B = 8'hC3; #100;
A = 8'h82; B = 8'hC4; #100;
A = 8'h82; B = 8'hC5; #100;
A = 8'h82; B = 8'hC6; #100;
A = 8'h82; B = 8'hC7; #100;
A = 8'h82; B = 8'hC8; #100;
A = 8'h82; B = 8'hC9; #100;
A = 8'h82; B = 8'hCA; #100;
A = 8'h82; B = 8'hCB; #100;
A = 8'h82; B = 8'hCC; #100;
A = 8'h82; B = 8'hCD; #100;
A = 8'h82; B = 8'hCE; #100;
A = 8'h82; B = 8'hCF; #100;
A = 8'h82; B = 8'hD0; #100;
A = 8'h82; B = 8'hD1; #100;
A = 8'h82; B = 8'hD2; #100;
A = 8'h82; B = 8'hD3; #100;
A = 8'h82; B = 8'hD4; #100;
A = 8'h82; B = 8'hD5; #100;
A = 8'h82; B = 8'hD6; #100;
A = 8'h82; B = 8'hD7; #100;
A = 8'h82; B = 8'hD8; #100;
A = 8'h82; B = 8'hD9; #100;
A = 8'h82; B = 8'hDA; #100;
A = 8'h82; B = 8'hDB; #100;
A = 8'h82; B = 8'hDC; #100;
A = 8'h82; B = 8'hDD; #100;
A = 8'h82; B = 8'hDE; #100;
A = 8'h82; B = 8'hDF; #100;
A = 8'h82; B = 8'hE0; #100;
A = 8'h82; B = 8'hE1; #100;
A = 8'h82; B = 8'hE2; #100;
A = 8'h82; B = 8'hE3; #100;
A = 8'h82; B = 8'hE4; #100;
A = 8'h82; B = 8'hE5; #100;
A = 8'h82; B = 8'hE6; #100;
A = 8'h82; B = 8'hE7; #100;
A = 8'h82; B = 8'hE8; #100;
A = 8'h82; B = 8'hE9; #100;
A = 8'h82; B = 8'hEA; #100;
A = 8'h82; B = 8'hEB; #100;
A = 8'h82; B = 8'hEC; #100;
A = 8'h82; B = 8'hED; #100;
A = 8'h82; B = 8'hEE; #100;
A = 8'h82; B = 8'hEF; #100;
A = 8'h82; B = 8'hF0; #100;
A = 8'h82; B = 8'hF1; #100;
A = 8'h82; B = 8'hF2; #100;
A = 8'h82; B = 8'hF3; #100;
A = 8'h82; B = 8'hF4; #100;
A = 8'h82; B = 8'hF5; #100;
A = 8'h82; B = 8'hF6; #100;
A = 8'h82; B = 8'hF7; #100;
A = 8'h82; B = 8'hF8; #100;
A = 8'h82; B = 8'hF9; #100;
A = 8'h82; B = 8'hFA; #100;
A = 8'h82; B = 8'hFB; #100;
A = 8'h82; B = 8'hFC; #100;
A = 8'h82; B = 8'hFD; #100;
A = 8'h82; B = 8'hFE; #100;
A = 8'h82; B = 8'hFF; #100;
A = 8'h83; B = 8'h0; #100;
A = 8'h83; B = 8'h1; #100;
A = 8'h83; B = 8'h2; #100;
A = 8'h83; B = 8'h3; #100;
A = 8'h83; B = 8'h4; #100;
A = 8'h83; B = 8'h5; #100;
A = 8'h83; B = 8'h6; #100;
A = 8'h83; B = 8'h7; #100;
A = 8'h83; B = 8'h8; #100;
A = 8'h83; B = 8'h9; #100;
A = 8'h83; B = 8'hA; #100;
A = 8'h83; B = 8'hB; #100;
A = 8'h83; B = 8'hC; #100;
A = 8'h83; B = 8'hD; #100;
A = 8'h83; B = 8'hE; #100;
A = 8'h83; B = 8'hF; #100;
A = 8'h83; B = 8'h10; #100;
A = 8'h83; B = 8'h11; #100;
A = 8'h83; B = 8'h12; #100;
A = 8'h83; B = 8'h13; #100;
A = 8'h83; B = 8'h14; #100;
A = 8'h83; B = 8'h15; #100;
A = 8'h83; B = 8'h16; #100;
A = 8'h83; B = 8'h17; #100;
A = 8'h83; B = 8'h18; #100;
A = 8'h83; B = 8'h19; #100;
A = 8'h83; B = 8'h1A; #100;
A = 8'h83; B = 8'h1B; #100;
A = 8'h83; B = 8'h1C; #100;
A = 8'h83; B = 8'h1D; #100;
A = 8'h83; B = 8'h1E; #100;
A = 8'h83; B = 8'h1F; #100;
A = 8'h83; B = 8'h20; #100;
A = 8'h83; B = 8'h21; #100;
A = 8'h83; B = 8'h22; #100;
A = 8'h83; B = 8'h23; #100;
A = 8'h83; B = 8'h24; #100;
A = 8'h83; B = 8'h25; #100;
A = 8'h83; B = 8'h26; #100;
A = 8'h83; B = 8'h27; #100;
A = 8'h83; B = 8'h28; #100;
A = 8'h83; B = 8'h29; #100;
A = 8'h83; B = 8'h2A; #100;
A = 8'h83; B = 8'h2B; #100;
A = 8'h83; B = 8'h2C; #100;
A = 8'h83; B = 8'h2D; #100;
A = 8'h83; B = 8'h2E; #100;
A = 8'h83; B = 8'h2F; #100;
A = 8'h83; B = 8'h30; #100;
A = 8'h83; B = 8'h31; #100;
A = 8'h83; B = 8'h32; #100;
A = 8'h83; B = 8'h33; #100;
A = 8'h83; B = 8'h34; #100;
A = 8'h83; B = 8'h35; #100;
A = 8'h83; B = 8'h36; #100;
A = 8'h83; B = 8'h37; #100;
A = 8'h83; B = 8'h38; #100;
A = 8'h83; B = 8'h39; #100;
A = 8'h83; B = 8'h3A; #100;
A = 8'h83; B = 8'h3B; #100;
A = 8'h83; B = 8'h3C; #100;
A = 8'h83; B = 8'h3D; #100;
A = 8'h83; B = 8'h3E; #100;
A = 8'h83; B = 8'h3F; #100;
A = 8'h83; B = 8'h40; #100;
A = 8'h83; B = 8'h41; #100;
A = 8'h83; B = 8'h42; #100;
A = 8'h83; B = 8'h43; #100;
A = 8'h83; B = 8'h44; #100;
A = 8'h83; B = 8'h45; #100;
A = 8'h83; B = 8'h46; #100;
A = 8'h83; B = 8'h47; #100;
A = 8'h83; B = 8'h48; #100;
A = 8'h83; B = 8'h49; #100;
A = 8'h83; B = 8'h4A; #100;
A = 8'h83; B = 8'h4B; #100;
A = 8'h83; B = 8'h4C; #100;
A = 8'h83; B = 8'h4D; #100;
A = 8'h83; B = 8'h4E; #100;
A = 8'h83; B = 8'h4F; #100;
A = 8'h83; B = 8'h50; #100;
A = 8'h83; B = 8'h51; #100;
A = 8'h83; B = 8'h52; #100;
A = 8'h83; B = 8'h53; #100;
A = 8'h83; B = 8'h54; #100;
A = 8'h83; B = 8'h55; #100;
A = 8'h83; B = 8'h56; #100;
A = 8'h83; B = 8'h57; #100;
A = 8'h83; B = 8'h58; #100;
A = 8'h83; B = 8'h59; #100;
A = 8'h83; B = 8'h5A; #100;
A = 8'h83; B = 8'h5B; #100;
A = 8'h83; B = 8'h5C; #100;
A = 8'h83; B = 8'h5D; #100;
A = 8'h83; B = 8'h5E; #100;
A = 8'h83; B = 8'h5F; #100;
A = 8'h83; B = 8'h60; #100;
A = 8'h83; B = 8'h61; #100;
A = 8'h83; B = 8'h62; #100;
A = 8'h83; B = 8'h63; #100;
A = 8'h83; B = 8'h64; #100;
A = 8'h83; B = 8'h65; #100;
A = 8'h83; B = 8'h66; #100;
A = 8'h83; B = 8'h67; #100;
A = 8'h83; B = 8'h68; #100;
A = 8'h83; B = 8'h69; #100;
A = 8'h83; B = 8'h6A; #100;
A = 8'h83; B = 8'h6B; #100;
A = 8'h83; B = 8'h6C; #100;
A = 8'h83; B = 8'h6D; #100;
A = 8'h83; B = 8'h6E; #100;
A = 8'h83; B = 8'h6F; #100;
A = 8'h83; B = 8'h70; #100;
A = 8'h83; B = 8'h71; #100;
A = 8'h83; B = 8'h72; #100;
A = 8'h83; B = 8'h73; #100;
A = 8'h83; B = 8'h74; #100;
A = 8'h83; B = 8'h75; #100;
A = 8'h83; B = 8'h76; #100;
A = 8'h83; B = 8'h77; #100;
A = 8'h83; B = 8'h78; #100;
A = 8'h83; B = 8'h79; #100;
A = 8'h83; B = 8'h7A; #100;
A = 8'h83; B = 8'h7B; #100;
A = 8'h83; B = 8'h7C; #100;
A = 8'h83; B = 8'h7D; #100;
A = 8'h83; B = 8'h7E; #100;
A = 8'h83; B = 8'h7F; #100;
A = 8'h83; B = 8'h80; #100;
A = 8'h83; B = 8'h81; #100;
A = 8'h83; B = 8'h82; #100;
A = 8'h83; B = 8'h83; #100;
A = 8'h83; B = 8'h84; #100;
A = 8'h83; B = 8'h85; #100;
A = 8'h83; B = 8'h86; #100;
A = 8'h83; B = 8'h87; #100;
A = 8'h83; B = 8'h88; #100;
A = 8'h83; B = 8'h89; #100;
A = 8'h83; B = 8'h8A; #100;
A = 8'h83; B = 8'h8B; #100;
A = 8'h83; B = 8'h8C; #100;
A = 8'h83; B = 8'h8D; #100;
A = 8'h83; B = 8'h8E; #100;
A = 8'h83; B = 8'h8F; #100;
A = 8'h83; B = 8'h90; #100;
A = 8'h83; B = 8'h91; #100;
A = 8'h83; B = 8'h92; #100;
A = 8'h83; B = 8'h93; #100;
A = 8'h83; B = 8'h94; #100;
A = 8'h83; B = 8'h95; #100;
A = 8'h83; B = 8'h96; #100;
A = 8'h83; B = 8'h97; #100;
A = 8'h83; B = 8'h98; #100;
A = 8'h83; B = 8'h99; #100;
A = 8'h83; B = 8'h9A; #100;
A = 8'h83; B = 8'h9B; #100;
A = 8'h83; B = 8'h9C; #100;
A = 8'h83; B = 8'h9D; #100;
A = 8'h83; B = 8'h9E; #100;
A = 8'h83; B = 8'h9F; #100;
A = 8'h83; B = 8'hA0; #100;
A = 8'h83; B = 8'hA1; #100;
A = 8'h83; B = 8'hA2; #100;
A = 8'h83; B = 8'hA3; #100;
A = 8'h83; B = 8'hA4; #100;
A = 8'h83; B = 8'hA5; #100;
A = 8'h83; B = 8'hA6; #100;
A = 8'h83; B = 8'hA7; #100;
A = 8'h83; B = 8'hA8; #100;
A = 8'h83; B = 8'hA9; #100;
A = 8'h83; B = 8'hAA; #100;
A = 8'h83; B = 8'hAB; #100;
A = 8'h83; B = 8'hAC; #100;
A = 8'h83; B = 8'hAD; #100;
A = 8'h83; B = 8'hAE; #100;
A = 8'h83; B = 8'hAF; #100;
A = 8'h83; B = 8'hB0; #100;
A = 8'h83; B = 8'hB1; #100;
A = 8'h83; B = 8'hB2; #100;
A = 8'h83; B = 8'hB3; #100;
A = 8'h83; B = 8'hB4; #100;
A = 8'h83; B = 8'hB5; #100;
A = 8'h83; B = 8'hB6; #100;
A = 8'h83; B = 8'hB7; #100;
A = 8'h83; B = 8'hB8; #100;
A = 8'h83; B = 8'hB9; #100;
A = 8'h83; B = 8'hBA; #100;
A = 8'h83; B = 8'hBB; #100;
A = 8'h83; B = 8'hBC; #100;
A = 8'h83; B = 8'hBD; #100;
A = 8'h83; B = 8'hBE; #100;
A = 8'h83; B = 8'hBF; #100;
A = 8'h83; B = 8'hC0; #100;
A = 8'h83; B = 8'hC1; #100;
A = 8'h83; B = 8'hC2; #100;
A = 8'h83; B = 8'hC3; #100;
A = 8'h83; B = 8'hC4; #100;
A = 8'h83; B = 8'hC5; #100;
A = 8'h83; B = 8'hC6; #100;
A = 8'h83; B = 8'hC7; #100;
A = 8'h83; B = 8'hC8; #100;
A = 8'h83; B = 8'hC9; #100;
A = 8'h83; B = 8'hCA; #100;
A = 8'h83; B = 8'hCB; #100;
A = 8'h83; B = 8'hCC; #100;
A = 8'h83; B = 8'hCD; #100;
A = 8'h83; B = 8'hCE; #100;
A = 8'h83; B = 8'hCF; #100;
A = 8'h83; B = 8'hD0; #100;
A = 8'h83; B = 8'hD1; #100;
A = 8'h83; B = 8'hD2; #100;
A = 8'h83; B = 8'hD3; #100;
A = 8'h83; B = 8'hD4; #100;
A = 8'h83; B = 8'hD5; #100;
A = 8'h83; B = 8'hD6; #100;
A = 8'h83; B = 8'hD7; #100;
A = 8'h83; B = 8'hD8; #100;
A = 8'h83; B = 8'hD9; #100;
A = 8'h83; B = 8'hDA; #100;
A = 8'h83; B = 8'hDB; #100;
A = 8'h83; B = 8'hDC; #100;
A = 8'h83; B = 8'hDD; #100;
A = 8'h83; B = 8'hDE; #100;
A = 8'h83; B = 8'hDF; #100;
A = 8'h83; B = 8'hE0; #100;
A = 8'h83; B = 8'hE1; #100;
A = 8'h83; B = 8'hE2; #100;
A = 8'h83; B = 8'hE3; #100;
A = 8'h83; B = 8'hE4; #100;
A = 8'h83; B = 8'hE5; #100;
A = 8'h83; B = 8'hE6; #100;
A = 8'h83; B = 8'hE7; #100;
A = 8'h83; B = 8'hE8; #100;
A = 8'h83; B = 8'hE9; #100;
A = 8'h83; B = 8'hEA; #100;
A = 8'h83; B = 8'hEB; #100;
A = 8'h83; B = 8'hEC; #100;
A = 8'h83; B = 8'hED; #100;
A = 8'h83; B = 8'hEE; #100;
A = 8'h83; B = 8'hEF; #100;
A = 8'h83; B = 8'hF0; #100;
A = 8'h83; B = 8'hF1; #100;
A = 8'h83; B = 8'hF2; #100;
A = 8'h83; B = 8'hF3; #100;
A = 8'h83; B = 8'hF4; #100;
A = 8'h83; B = 8'hF5; #100;
A = 8'h83; B = 8'hF6; #100;
A = 8'h83; B = 8'hF7; #100;
A = 8'h83; B = 8'hF8; #100;
A = 8'h83; B = 8'hF9; #100;
A = 8'h83; B = 8'hFA; #100;
A = 8'h83; B = 8'hFB; #100;
A = 8'h83; B = 8'hFC; #100;
A = 8'h83; B = 8'hFD; #100;
A = 8'h83; B = 8'hFE; #100;
A = 8'h83; B = 8'hFF; #100;
A = 8'h84; B = 8'h0; #100;
A = 8'h84; B = 8'h1; #100;
A = 8'h84; B = 8'h2; #100;
A = 8'h84; B = 8'h3; #100;
A = 8'h84; B = 8'h4; #100;
A = 8'h84; B = 8'h5; #100;
A = 8'h84; B = 8'h6; #100;
A = 8'h84; B = 8'h7; #100;
A = 8'h84; B = 8'h8; #100;
A = 8'h84; B = 8'h9; #100;
A = 8'h84; B = 8'hA; #100;
A = 8'h84; B = 8'hB; #100;
A = 8'h84; B = 8'hC; #100;
A = 8'h84; B = 8'hD; #100;
A = 8'h84; B = 8'hE; #100;
A = 8'h84; B = 8'hF; #100;
A = 8'h84; B = 8'h10; #100;
A = 8'h84; B = 8'h11; #100;
A = 8'h84; B = 8'h12; #100;
A = 8'h84; B = 8'h13; #100;
A = 8'h84; B = 8'h14; #100;
A = 8'h84; B = 8'h15; #100;
A = 8'h84; B = 8'h16; #100;
A = 8'h84; B = 8'h17; #100;
A = 8'h84; B = 8'h18; #100;
A = 8'h84; B = 8'h19; #100;
A = 8'h84; B = 8'h1A; #100;
A = 8'h84; B = 8'h1B; #100;
A = 8'h84; B = 8'h1C; #100;
A = 8'h84; B = 8'h1D; #100;
A = 8'h84; B = 8'h1E; #100;
A = 8'h84; B = 8'h1F; #100;
A = 8'h84; B = 8'h20; #100;
A = 8'h84; B = 8'h21; #100;
A = 8'h84; B = 8'h22; #100;
A = 8'h84; B = 8'h23; #100;
A = 8'h84; B = 8'h24; #100;
A = 8'h84; B = 8'h25; #100;
A = 8'h84; B = 8'h26; #100;
A = 8'h84; B = 8'h27; #100;
A = 8'h84; B = 8'h28; #100;
A = 8'h84; B = 8'h29; #100;
A = 8'h84; B = 8'h2A; #100;
A = 8'h84; B = 8'h2B; #100;
A = 8'h84; B = 8'h2C; #100;
A = 8'h84; B = 8'h2D; #100;
A = 8'h84; B = 8'h2E; #100;
A = 8'h84; B = 8'h2F; #100;
A = 8'h84; B = 8'h30; #100;
A = 8'h84; B = 8'h31; #100;
A = 8'h84; B = 8'h32; #100;
A = 8'h84; B = 8'h33; #100;
A = 8'h84; B = 8'h34; #100;
A = 8'h84; B = 8'h35; #100;
A = 8'h84; B = 8'h36; #100;
A = 8'h84; B = 8'h37; #100;
A = 8'h84; B = 8'h38; #100;
A = 8'h84; B = 8'h39; #100;
A = 8'h84; B = 8'h3A; #100;
A = 8'h84; B = 8'h3B; #100;
A = 8'h84; B = 8'h3C; #100;
A = 8'h84; B = 8'h3D; #100;
A = 8'h84; B = 8'h3E; #100;
A = 8'h84; B = 8'h3F; #100;
A = 8'h84; B = 8'h40; #100;
A = 8'h84; B = 8'h41; #100;
A = 8'h84; B = 8'h42; #100;
A = 8'h84; B = 8'h43; #100;
A = 8'h84; B = 8'h44; #100;
A = 8'h84; B = 8'h45; #100;
A = 8'h84; B = 8'h46; #100;
A = 8'h84; B = 8'h47; #100;
A = 8'h84; B = 8'h48; #100;
A = 8'h84; B = 8'h49; #100;
A = 8'h84; B = 8'h4A; #100;
A = 8'h84; B = 8'h4B; #100;
A = 8'h84; B = 8'h4C; #100;
A = 8'h84; B = 8'h4D; #100;
A = 8'h84; B = 8'h4E; #100;
A = 8'h84; B = 8'h4F; #100;
A = 8'h84; B = 8'h50; #100;
A = 8'h84; B = 8'h51; #100;
A = 8'h84; B = 8'h52; #100;
A = 8'h84; B = 8'h53; #100;
A = 8'h84; B = 8'h54; #100;
A = 8'h84; B = 8'h55; #100;
A = 8'h84; B = 8'h56; #100;
A = 8'h84; B = 8'h57; #100;
A = 8'h84; B = 8'h58; #100;
A = 8'h84; B = 8'h59; #100;
A = 8'h84; B = 8'h5A; #100;
A = 8'h84; B = 8'h5B; #100;
A = 8'h84; B = 8'h5C; #100;
A = 8'h84; B = 8'h5D; #100;
A = 8'h84; B = 8'h5E; #100;
A = 8'h84; B = 8'h5F; #100;
A = 8'h84; B = 8'h60; #100;
A = 8'h84; B = 8'h61; #100;
A = 8'h84; B = 8'h62; #100;
A = 8'h84; B = 8'h63; #100;
A = 8'h84; B = 8'h64; #100;
A = 8'h84; B = 8'h65; #100;
A = 8'h84; B = 8'h66; #100;
A = 8'h84; B = 8'h67; #100;
A = 8'h84; B = 8'h68; #100;
A = 8'h84; B = 8'h69; #100;
A = 8'h84; B = 8'h6A; #100;
A = 8'h84; B = 8'h6B; #100;
A = 8'h84; B = 8'h6C; #100;
A = 8'h84; B = 8'h6D; #100;
A = 8'h84; B = 8'h6E; #100;
A = 8'h84; B = 8'h6F; #100;
A = 8'h84; B = 8'h70; #100;
A = 8'h84; B = 8'h71; #100;
A = 8'h84; B = 8'h72; #100;
A = 8'h84; B = 8'h73; #100;
A = 8'h84; B = 8'h74; #100;
A = 8'h84; B = 8'h75; #100;
A = 8'h84; B = 8'h76; #100;
A = 8'h84; B = 8'h77; #100;
A = 8'h84; B = 8'h78; #100;
A = 8'h84; B = 8'h79; #100;
A = 8'h84; B = 8'h7A; #100;
A = 8'h84; B = 8'h7B; #100;
A = 8'h84; B = 8'h7C; #100;
A = 8'h84; B = 8'h7D; #100;
A = 8'h84; B = 8'h7E; #100;
A = 8'h84; B = 8'h7F; #100;
A = 8'h84; B = 8'h80; #100;
A = 8'h84; B = 8'h81; #100;
A = 8'h84; B = 8'h82; #100;
A = 8'h84; B = 8'h83; #100;
A = 8'h84; B = 8'h84; #100;
A = 8'h84; B = 8'h85; #100;
A = 8'h84; B = 8'h86; #100;
A = 8'h84; B = 8'h87; #100;
A = 8'h84; B = 8'h88; #100;
A = 8'h84; B = 8'h89; #100;
A = 8'h84; B = 8'h8A; #100;
A = 8'h84; B = 8'h8B; #100;
A = 8'h84; B = 8'h8C; #100;
A = 8'h84; B = 8'h8D; #100;
A = 8'h84; B = 8'h8E; #100;
A = 8'h84; B = 8'h8F; #100;
A = 8'h84; B = 8'h90; #100;
A = 8'h84; B = 8'h91; #100;
A = 8'h84; B = 8'h92; #100;
A = 8'h84; B = 8'h93; #100;
A = 8'h84; B = 8'h94; #100;
A = 8'h84; B = 8'h95; #100;
A = 8'h84; B = 8'h96; #100;
A = 8'h84; B = 8'h97; #100;
A = 8'h84; B = 8'h98; #100;
A = 8'h84; B = 8'h99; #100;
A = 8'h84; B = 8'h9A; #100;
A = 8'h84; B = 8'h9B; #100;
A = 8'h84; B = 8'h9C; #100;
A = 8'h84; B = 8'h9D; #100;
A = 8'h84; B = 8'h9E; #100;
A = 8'h84; B = 8'h9F; #100;
A = 8'h84; B = 8'hA0; #100;
A = 8'h84; B = 8'hA1; #100;
A = 8'h84; B = 8'hA2; #100;
A = 8'h84; B = 8'hA3; #100;
A = 8'h84; B = 8'hA4; #100;
A = 8'h84; B = 8'hA5; #100;
A = 8'h84; B = 8'hA6; #100;
A = 8'h84; B = 8'hA7; #100;
A = 8'h84; B = 8'hA8; #100;
A = 8'h84; B = 8'hA9; #100;
A = 8'h84; B = 8'hAA; #100;
A = 8'h84; B = 8'hAB; #100;
A = 8'h84; B = 8'hAC; #100;
A = 8'h84; B = 8'hAD; #100;
A = 8'h84; B = 8'hAE; #100;
A = 8'h84; B = 8'hAF; #100;
A = 8'h84; B = 8'hB0; #100;
A = 8'h84; B = 8'hB1; #100;
A = 8'h84; B = 8'hB2; #100;
A = 8'h84; B = 8'hB3; #100;
A = 8'h84; B = 8'hB4; #100;
A = 8'h84; B = 8'hB5; #100;
A = 8'h84; B = 8'hB6; #100;
A = 8'h84; B = 8'hB7; #100;
A = 8'h84; B = 8'hB8; #100;
A = 8'h84; B = 8'hB9; #100;
A = 8'h84; B = 8'hBA; #100;
A = 8'h84; B = 8'hBB; #100;
A = 8'h84; B = 8'hBC; #100;
A = 8'h84; B = 8'hBD; #100;
A = 8'h84; B = 8'hBE; #100;
A = 8'h84; B = 8'hBF; #100;
A = 8'h84; B = 8'hC0; #100;
A = 8'h84; B = 8'hC1; #100;
A = 8'h84; B = 8'hC2; #100;
A = 8'h84; B = 8'hC3; #100;
A = 8'h84; B = 8'hC4; #100;
A = 8'h84; B = 8'hC5; #100;
A = 8'h84; B = 8'hC6; #100;
A = 8'h84; B = 8'hC7; #100;
A = 8'h84; B = 8'hC8; #100;
A = 8'h84; B = 8'hC9; #100;
A = 8'h84; B = 8'hCA; #100;
A = 8'h84; B = 8'hCB; #100;
A = 8'h84; B = 8'hCC; #100;
A = 8'h84; B = 8'hCD; #100;
A = 8'h84; B = 8'hCE; #100;
A = 8'h84; B = 8'hCF; #100;
A = 8'h84; B = 8'hD0; #100;
A = 8'h84; B = 8'hD1; #100;
A = 8'h84; B = 8'hD2; #100;
A = 8'h84; B = 8'hD3; #100;
A = 8'h84; B = 8'hD4; #100;
A = 8'h84; B = 8'hD5; #100;
A = 8'h84; B = 8'hD6; #100;
A = 8'h84; B = 8'hD7; #100;
A = 8'h84; B = 8'hD8; #100;
A = 8'h84; B = 8'hD9; #100;
A = 8'h84; B = 8'hDA; #100;
A = 8'h84; B = 8'hDB; #100;
A = 8'h84; B = 8'hDC; #100;
A = 8'h84; B = 8'hDD; #100;
A = 8'h84; B = 8'hDE; #100;
A = 8'h84; B = 8'hDF; #100;
A = 8'h84; B = 8'hE0; #100;
A = 8'h84; B = 8'hE1; #100;
A = 8'h84; B = 8'hE2; #100;
A = 8'h84; B = 8'hE3; #100;
A = 8'h84; B = 8'hE4; #100;
A = 8'h84; B = 8'hE5; #100;
A = 8'h84; B = 8'hE6; #100;
A = 8'h84; B = 8'hE7; #100;
A = 8'h84; B = 8'hE8; #100;
A = 8'h84; B = 8'hE9; #100;
A = 8'h84; B = 8'hEA; #100;
A = 8'h84; B = 8'hEB; #100;
A = 8'h84; B = 8'hEC; #100;
A = 8'h84; B = 8'hED; #100;
A = 8'h84; B = 8'hEE; #100;
A = 8'h84; B = 8'hEF; #100;
A = 8'h84; B = 8'hF0; #100;
A = 8'h84; B = 8'hF1; #100;
A = 8'h84; B = 8'hF2; #100;
A = 8'h84; B = 8'hF3; #100;
A = 8'h84; B = 8'hF4; #100;
A = 8'h84; B = 8'hF5; #100;
A = 8'h84; B = 8'hF6; #100;
A = 8'h84; B = 8'hF7; #100;
A = 8'h84; B = 8'hF8; #100;
A = 8'h84; B = 8'hF9; #100;
A = 8'h84; B = 8'hFA; #100;
A = 8'h84; B = 8'hFB; #100;
A = 8'h84; B = 8'hFC; #100;
A = 8'h84; B = 8'hFD; #100;
A = 8'h84; B = 8'hFE; #100;
A = 8'h84; B = 8'hFF; #100;
A = 8'h85; B = 8'h0; #100;
A = 8'h85; B = 8'h1; #100;
A = 8'h85; B = 8'h2; #100;
A = 8'h85; B = 8'h3; #100;
A = 8'h85; B = 8'h4; #100;
A = 8'h85; B = 8'h5; #100;
A = 8'h85; B = 8'h6; #100;
A = 8'h85; B = 8'h7; #100;
A = 8'h85; B = 8'h8; #100;
A = 8'h85; B = 8'h9; #100;
A = 8'h85; B = 8'hA; #100;
A = 8'h85; B = 8'hB; #100;
A = 8'h85; B = 8'hC; #100;
A = 8'h85; B = 8'hD; #100;
A = 8'h85; B = 8'hE; #100;
A = 8'h85; B = 8'hF; #100;
A = 8'h85; B = 8'h10; #100;
A = 8'h85; B = 8'h11; #100;
A = 8'h85; B = 8'h12; #100;
A = 8'h85; B = 8'h13; #100;
A = 8'h85; B = 8'h14; #100;
A = 8'h85; B = 8'h15; #100;
A = 8'h85; B = 8'h16; #100;
A = 8'h85; B = 8'h17; #100;
A = 8'h85; B = 8'h18; #100;
A = 8'h85; B = 8'h19; #100;
A = 8'h85; B = 8'h1A; #100;
A = 8'h85; B = 8'h1B; #100;
A = 8'h85; B = 8'h1C; #100;
A = 8'h85; B = 8'h1D; #100;
A = 8'h85; B = 8'h1E; #100;
A = 8'h85; B = 8'h1F; #100;
A = 8'h85; B = 8'h20; #100;
A = 8'h85; B = 8'h21; #100;
A = 8'h85; B = 8'h22; #100;
A = 8'h85; B = 8'h23; #100;
A = 8'h85; B = 8'h24; #100;
A = 8'h85; B = 8'h25; #100;
A = 8'h85; B = 8'h26; #100;
A = 8'h85; B = 8'h27; #100;
A = 8'h85; B = 8'h28; #100;
A = 8'h85; B = 8'h29; #100;
A = 8'h85; B = 8'h2A; #100;
A = 8'h85; B = 8'h2B; #100;
A = 8'h85; B = 8'h2C; #100;
A = 8'h85; B = 8'h2D; #100;
A = 8'h85; B = 8'h2E; #100;
A = 8'h85; B = 8'h2F; #100;
A = 8'h85; B = 8'h30; #100;
A = 8'h85; B = 8'h31; #100;
A = 8'h85; B = 8'h32; #100;
A = 8'h85; B = 8'h33; #100;
A = 8'h85; B = 8'h34; #100;
A = 8'h85; B = 8'h35; #100;
A = 8'h85; B = 8'h36; #100;
A = 8'h85; B = 8'h37; #100;
A = 8'h85; B = 8'h38; #100;
A = 8'h85; B = 8'h39; #100;
A = 8'h85; B = 8'h3A; #100;
A = 8'h85; B = 8'h3B; #100;
A = 8'h85; B = 8'h3C; #100;
A = 8'h85; B = 8'h3D; #100;
A = 8'h85; B = 8'h3E; #100;
A = 8'h85; B = 8'h3F; #100;
A = 8'h85; B = 8'h40; #100;
A = 8'h85; B = 8'h41; #100;
A = 8'h85; B = 8'h42; #100;
A = 8'h85; B = 8'h43; #100;
A = 8'h85; B = 8'h44; #100;
A = 8'h85; B = 8'h45; #100;
A = 8'h85; B = 8'h46; #100;
A = 8'h85; B = 8'h47; #100;
A = 8'h85; B = 8'h48; #100;
A = 8'h85; B = 8'h49; #100;
A = 8'h85; B = 8'h4A; #100;
A = 8'h85; B = 8'h4B; #100;
A = 8'h85; B = 8'h4C; #100;
A = 8'h85; B = 8'h4D; #100;
A = 8'h85; B = 8'h4E; #100;
A = 8'h85; B = 8'h4F; #100;
A = 8'h85; B = 8'h50; #100;
A = 8'h85; B = 8'h51; #100;
A = 8'h85; B = 8'h52; #100;
A = 8'h85; B = 8'h53; #100;
A = 8'h85; B = 8'h54; #100;
A = 8'h85; B = 8'h55; #100;
A = 8'h85; B = 8'h56; #100;
A = 8'h85; B = 8'h57; #100;
A = 8'h85; B = 8'h58; #100;
A = 8'h85; B = 8'h59; #100;
A = 8'h85; B = 8'h5A; #100;
A = 8'h85; B = 8'h5B; #100;
A = 8'h85; B = 8'h5C; #100;
A = 8'h85; B = 8'h5D; #100;
A = 8'h85; B = 8'h5E; #100;
A = 8'h85; B = 8'h5F; #100;
A = 8'h85; B = 8'h60; #100;
A = 8'h85; B = 8'h61; #100;
A = 8'h85; B = 8'h62; #100;
A = 8'h85; B = 8'h63; #100;
A = 8'h85; B = 8'h64; #100;
A = 8'h85; B = 8'h65; #100;
A = 8'h85; B = 8'h66; #100;
A = 8'h85; B = 8'h67; #100;
A = 8'h85; B = 8'h68; #100;
A = 8'h85; B = 8'h69; #100;
A = 8'h85; B = 8'h6A; #100;
A = 8'h85; B = 8'h6B; #100;
A = 8'h85; B = 8'h6C; #100;
A = 8'h85; B = 8'h6D; #100;
A = 8'h85; B = 8'h6E; #100;
A = 8'h85; B = 8'h6F; #100;
A = 8'h85; B = 8'h70; #100;
A = 8'h85; B = 8'h71; #100;
A = 8'h85; B = 8'h72; #100;
A = 8'h85; B = 8'h73; #100;
A = 8'h85; B = 8'h74; #100;
A = 8'h85; B = 8'h75; #100;
A = 8'h85; B = 8'h76; #100;
A = 8'h85; B = 8'h77; #100;
A = 8'h85; B = 8'h78; #100;
A = 8'h85; B = 8'h79; #100;
A = 8'h85; B = 8'h7A; #100;
A = 8'h85; B = 8'h7B; #100;
A = 8'h85; B = 8'h7C; #100;
A = 8'h85; B = 8'h7D; #100;
A = 8'h85; B = 8'h7E; #100;
A = 8'h85; B = 8'h7F; #100;
A = 8'h85; B = 8'h80; #100;
A = 8'h85; B = 8'h81; #100;
A = 8'h85; B = 8'h82; #100;
A = 8'h85; B = 8'h83; #100;
A = 8'h85; B = 8'h84; #100;
A = 8'h85; B = 8'h85; #100;
A = 8'h85; B = 8'h86; #100;
A = 8'h85; B = 8'h87; #100;
A = 8'h85; B = 8'h88; #100;
A = 8'h85; B = 8'h89; #100;
A = 8'h85; B = 8'h8A; #100;
A = 8'h85; B = 8'h8B; #100;
A = 8'h85; B = 8'h8C; #100;
A = 8'h85; B = 8'h8D; #100;
A = 8'h85; B = 8'h8E; #100;
A = 8'h85; B = 8'h8F; #100;
A = 8'h85; B = 8'h90; #100;
A = 8'h85; B = 8'h91; #100;
A = 8'h85; B = 8'h92; #100;
A = 8'h85; B = 8'h93; #100;
A = 8'h85; B = 8'h94; #100;
A = 8'h85; B = 8'h95; #100;
A = 8'h85; B = 8'h96; #100;
A = 8'h85; B = 8'h97; #100;
A = 8'h85; B = 8'h98; #100;
A = 8'h85; B = 8'h99; #100;
A = 8'h85; B = 8'h9A; #100;
A = 8'h85; B = 8'h9B; #100;
A = 8'h85; B = 8'h9C; #100;
A = 8'h85; B = 8'h9D; #100;
A = 8'h85; B = 8'h9E; #100;
A = 8'h85; B = 8'h9F; #100;
A = 8'h85; B = 8'hA0; #100;
A = 8'h85; B = 8'hA1; #100;
A = 8'h85; B = 8'hA2; #100;
A = 8'h85; B = 8'hA3; #100;
A = 8'h85; B = 8'hA4; #100;
A = 8'h85; B = 8'hA5; #100;
A = 8'h85; B = 8'hA6; #100;
A = 8'h85; B = 8'hA7; #100;
A = 8'h85; B = 8'hA8; #100;
A = 8'h85; B = 8'hA9; #100;
A = 8'h85; B = 8'hAA; #100;
A = 8'h85; B = 8'hAB; #100;
A = 8'h85; B = 8'hAC; #100;
A = 8'h85; B = 8'hAD; #100;
A = 8'h85; B = 8'hAE; #100;
A = 8'h85; B = 8'hAF; #100;
A = 8'h85; B = 8'hB0; #100;
A = 8'h85; B = 8'hB1; #100;
A = 8'h85; B = 8'hB2; #100;
A = 8'h85; B = 8'hB3; #100;
A = 8'h85; B = 8'hB4; #100;
A = 8'h85; B = 8'hB5; #100;
A = 8'h85; B = 8'hB6; #100;
A = 8'h85; B = 8'hB7; #100;
A = 8'h85; B = 8'hB8; #100;
A = 8'h85; B = 8'hB9; #100;
A = 8'h85; B = 8'hBA; #100;
A = 8'h85; B = 8'hBB; #100;
A = 8'h85; B = 8'hBC; #100;
A = 8'h85; B = 8'hBD; #100;
A = 8'h85; B = 8'hBE; #100;
A = 8'h85; B = 8'hBF; #100;
A = 8'h85; B = 8'hC0; #100;
A = 8'h85; B = 8'hC1; #100;
A = 8'h85; B = 8'hC2; #100;
A = 8'h85; B = 8'hC3; #100;
A = 8'h85; B = 8'hC4; #100;
A = 8'h85; B = 8'hC5; #100;
A = 8'h85; B = 8'hC6; #100;
A = 8'h85; B = 8'hC7; #100;
A = 8'h85; B = 8'hC8; #100;
A = 8'h85; B = 8'hC9; #100;
A = 8'h85; B = 8'hCA; #100;
A = 8'h85; B = 8'hCB; #100;
A = 8'h85; B = 8'hCC; #100;
A = 8'h85; B = 8'hCD; #100;
A = 8'h85; B = 8'hCE; #100;
A = 8'h85; B = 8'hCF; #100;
A = 8'h85; B = 8'hD0; #100;
A = 8'h85; B = 8'hD1; #100;
A = 8'h85; B = 8'hD2; #100;
A = 8'h85; B = 8'hD3; #100;
A = 8'h85; B = 8'hD4; #100;
A = 8'h85; B = 8'hD5; #100;
A = 8'h85; B = 8'hD6; #100;
A = 8'h85; B = 8'hD7; #100;
A = 8'h85; B = 8'hD8; #100;
A = 8'h85; B = 8'hD9; #100;
A = 8'h85; B = 8'hDA; #100;
A = 8'h85; B = 8'hDB; #100;
A = 8'h85; B = 8'hDC; #100;
A = 8'h85; B = 8'hDD; #100;
A = 8'h85; B = 8'hDE; #100;
A = 8'h85; B = 8'hDF; #100;
A = 8'h85; B = 8'hE0; #100;
A = 8'h85; B = 8'hE1; #100;
A = 8'h85; B = 8'hE2; #100;
A = 8'h85; B = 8'hE3; #100;
A = 8'h85; B = 8'hE4; #100;
A = 8'h85; B = 8'hE5; #100;
A = 8'h85; B = 8'hE6; #100;
A = 8'h85; B = 8'hE7; #100;
A = 8'h85; B = 8'hE8; #100;
A = 8'h85; B = 8'hE9; #100;
A = 8'h85; B = 8'hEA; #100;
A = 8'h85; B = 8'hEB; #100;
A = 8'h85; B = 8'hEC; #100;
A = 8'h85; B = 8'hED; #100;
A = 8'h85; B = 8'hEE; #100;
A = 8'h85; B = 8'hEF; #100;
A = 8'h85; B = 8'hF0; #100;
A = 8'h85; B = 8'hF1; #100;
A = 8'h85; B = 8'hF2; #100;
A = 8'h85; B = 8'hF3; #100;
A = 8'h85; B = 8'hF4; #100;
A = 8'h85; B = 8'hF5; #100;
A = 8'h85; B = 8'hF6; #100;
A = 8'h85; B = 8'hF7; #100;
A = 8'h85; B = 8'hF8; #100;
A = 8'h85; B = 8'hF9; #100;
A = 8'h85; B = 8'hFA; #100;
A = 8'h85; B = 8'hFB; #100;
A = 8'h85; B = 8'hFC; #100;
A = 8'h85; B = 8'hFD; #100;
A = 8'h85; B = 8'hFE; #100;
A = 8'h85; B = 8'hFF; #100;
A = 8'h86; B = 8'h0; #100;
A = 8'h86; B = 8'h1; #100;
A = 8'h86; B = 8'h2; #100;
A = 8'h86; B = 8'h3; #100;
A = 8'h86; B = 8'h4; #100;
A = 8'h86; B = 8'h5; #100;
A = 8'h86; B = 8'h6; #100;
A = 8'h86; B = 8'h7; #100;
A = 8'h86; B = 8'h8; #100;
A = 8'h86; B = 8'h9; #100;
A = 8'h86; B = 8'hA; #100;
A = 8'h86; B = 8'hB; #100;
A = 8'h86; B = 8'hC; #100;
A = 8'h86; B = 8'hD; #100;
A = 8'h86; B = 8'hE; #100;
A = 8'h86; B = 8'hF; #100;
A = 8'h86; B = 8'h10; #100;
A = 8'h86; B = 8'h11; #100;
A = 8'h86; B = 8'h12; #100;
A = 8'h86; B = 8'h13; #100;
A = 8'h86; B = 8'h14; #100;
A = 8'h86; B = 8'h15; #100;
A = 8'h86; B = 8'h16; #100;
A = 8'h86; B = 8'h17; #100;
A = 8'h86; B = 8'h18; #100;
A = 8'h86; B = 8'h19; #100;
A = 8'h86; B = 8'h1A; #100;
A = 8'h86; B = 8'h1B; #100;
A = 8'h86; B = 8'h1C; #100;
A = 8'h86; B = 8'h1D; #100;
A = 8'h86; B = 8'h1E; #100;
A = 8'h86; B = 8'h1F; #100;
A = 8'h86; B = 8'h20; #100;
A = 8'h86; B = 8'h21; #100;
A = 8'h86; B = 8'h22; #100;
A = 8'h86; B = 8'h23; #100;
A = 8'h86; B = 8'h24; #100;
A = 8'h86; B = 8'h25; #100;
A = 8'h86; B = 8'h26; #100;
A = 8'h86; B = 8'h27; #100;
A = 8'h86; B = 8'h28; #100;
A = 8'h86; B = 8'h29; #100;
A = 8'h86; B = 8'h2A; #100;
A = 8'h86; B = 8'h2B; #100;
A = 8'h86; B = 8'h2C; #100;
A = 8'h86; B = 8'h2D; #100;
A = 8'h86; B = 8'h2E; #100;
A = 8'h86; B = 8'h2F; #100;
A = 8'h86; B = 8'h30; #100;
A = 8'h86; B = 8'h31; #100;
A = 8'h86; B = 8'h32; #100;
A = 8'h86; B = 8'h33; #100;
A = 8'h86; B = 8'h34; #100;
A = 8'h86; B = 8'h35; #100;
A = 8'h86; B = 8'h36; #100;
A = 8'h86; B = 8'h37; #100;
A = 8'h86; B = 8'h38; #100;
A = 8'h86; B = 8'h39; #100;
A = 8'h86; B = 8'h3A; #100;
A = 8'h86; B = 8'h3B; #100;
A = 8'h86; B = 8'h3C; #100;
A = 8'h86; B = 8'h3D; #100;
A = 8'h86; B = 8'h3E; #100;
A = 8'h86; B = 8'h3F; #100;
A = 8'h86; B = 8'h40; #100;
A = 8'h86; B = 8'h41; #100;
A = 8'h86; B = 8'h42; #100;
A = 8'h86; B = 8'h43; #100;
A = 8'h86; B = 8'h44; #100;
A = 8'h86; B = 8'h45; #100;
A = 8'h86; B = 8'h46; #100;
A = 8'h86; B = 8'h47; #100;
A = 8'h86; B = 8'h48; #100;
A = 8'h86; B = 8'h49; #100;
A = 8'h86; B = 8'h4A; #100;
A = 8'h86; B = 8'h4B; #100;
A = 8'h86; B = 8'h4C; #100;
A = 8'h86; B = 8'h4D; #100;
A = 8'h86; B = 8'h4E; #100;
A = 8'h86; B = 8'h4F; #100;
A = 8'h86; B = 8'h50; #100;
A = 8'h86; B = 8'h51; #100;
A = 8'h86; B = 8'h52; #100;
A = 8'h86; B = 8'h53; #100;
A = 8'h86; B = 8'h54; #100;
A = 8'h86; B = 8'h55; #100;
A = 8'h86; B = 8'h56; #100;
A = 8'h86; B = 8'h57; #100;
A = 8'h86; B = 8'h58; #100;
A = 8'h86; B = 8'h59; #100;
A = 8'h86; B = 8'h5A; #100;
A = 8'h86; B = 8'h5B; #100;
A = 8'h86; B = 8'h5C; #100;
A = 8'h86; B = 8'h5D; #100;
A = 8'h86; B = 8'h5E; #100;
A = 8'h86; B = 8'h5F; #100;
A = 8'h86; B = 8'h60; #100;
A = 8'h86; B = 8'h61; #100;
A = 8'h86; B = 8'h62; #100;
A = 8'h86; B = 8'h63; #100;
A = 8'h86; B = 8'h64; #100;
A = 8'h86; B = 8'h65; #100;
A = 8'h86; B = 8'h66; #100;
A = 8'h86; B = 8'h67; #100;
A = 8'h86; B = 8'h68; #100;
A = 8'h86; B = 8'h69; #100;
A = 8'h86; B = 8'h6A; #100;
A = 8'h86; B = 8'h6B; #100;
A = 8'h86; B = 8'h6C; #100;
A = 8'h86; B = 8'h6D; #100;
A = 8'h86; B = 8'h6E; #100;
A = 8'h86; B = 8'h6F; #100;
A = 8'h86; B = 8'h70; #100;
A = 8'h86; B = 8'h71; #100;
A = 8'h86; B = 8'h72; #100;
A = 8'h86; B = 8'h73; #100;
A = 8'h86; B = 8'h74; #100;
A = 8'h86; B = 8'h75; #100;
A = 8'h86; B = 8'h76; #100;
A = 8'h86; B = 8'h77; #100;
A = 8'h86; B = 8'h78; #100;
A = 8'h86; B = 8'h79; #100;
A = 8'h86; B = 8'h7A; #100;
A = 8'h86; B = 8'h7B; #100;
A = 8'h86; B = 8'h7C; #100;
A = 8'h86; B = 8'h7D; #100;
A = 8'h86; B = 8'h7E; #100;
A = 8'h86; B = 8'h7F; #100;
A = 8'h86; B = 8'h80; #100;
A = 8'h86; B = 8'h81; #100;
A = 8'h86; B = 8'h82; #100;
A = 8'h86; B = 8'h83; #100;
A = 8'h86; B = 8'h84; #100;
A = 8'h86; B = 8'h85; #100;
A = 8'h86; B = 8'h86; #100;
A = 8'h86; B = 8'h87; #100;
A = 8'h86; B = 8'h88; #100;
A = 8'h86; B = 8'h89; #100;
A = 8'h86; B = 8'h8A; #100;
A = 8'h86; B = 8'h8B; #100;
A = 8'h86; B = 8'h8C; #100;
A = 8'h86; B = 8'h8D; #100;
A = 8'h86; B = 8'h8E; #100;
A = 8'h86; B = 8'h8F; #100;
A = 8'h86; B = 8'h90; #100;
A = 8'h86; B = 8'h91; #100;
A = 8'h86; B = 8'h92; #100;
A = 8'h86; B = 8'h93; #100;
A = 8'h86; B = 8'h94; #100;
A = 8'h86; B = 8'h95; #100;
A = 8'h86; B = 8'h96; #100;
A = 8'h86; B = 8'h97; #100;
A = 8'h86; B = 8'h98; #100;
A = 8'h86; B = 8'h99; #100;
A = 8'h86; B = 8'h9A; #100;
A = 8'h86; B = 8'h9B; #100;
A = 8'h86; B = 8'h9C; #100;
A = 8'h86; B = 8'h9D; #100;
A = 8'h86; B = 8'h9E; #100;
A = 8'h86; B = 8'h9F; #100;
A = 8'h86; B = 8'hA0; #100;
A = 8'h86; B = 8'hA1; #100;
A = 8'h86; B = 8'hA2; #100;
A = 8'h86; B = 8'hA3; #100;
A = 8'h86; B = 8'hA4; #100;
A = 8'h86; B = 8'hA5; #100;
A = 8'h86; B = 8'hA6; #100;
A = 8'h86; B = 8'hA7; #100;
A = 8'h86; B = 8'hA8; #100;
A = 8'h86; B = 8'hA9; #100;
A = 8'h86; B = 8'hAA; #100;
A = 8'h86; B = 8'hAB; #100;
A = 8'h86; B = 8'hAC; #100;
A = 8'h86; B = 8'hAD; #100;
A = 8'h86; B = 8'hAE; #100;
A = 8'h86; B = 8'hAF; #100;
A = 8'h86; B = 8'hB0; #100;
A = 8'h86; B = 8'hB1; #100;
A = 8'h86; B = 8'hB2; #100;
A = 8'h86; B = 8'hB3; #100;
A = 8'h86; B = 8'hB4; #100;
A = 8'h86; B = 8'hB5; #100;
A = 8'h86; B = 8'hB6; #100;
A = 8'h86; B = 8'hB7; #100;
A = 8'h86; B = 8'hB8; #100;
A = 8'h86; B = 8'hB9; #100;
A = 8'h86; B = 8'hBA; #100;
A = 8'h86; B = 8'hBB; #100;
A = 8'h86; B = 8'hBC; #100;
A = 8'h86; B = 8'hBD; #100;
A = 8'h86; B = 8'hBE; #100;
A = 8'h86; B = 8'hBF; #100;
A = 8'h86; B = 8'hC0; #100;
A = 8'h86; B = 8'hC1; #100;
A = 8'h86; B = 8'hC2; #100;
A = 8'h86; B = 8'hC3; #100;
A = 8'h86; B = 8'hC4; #100;
A = 8'h86; B = 8'hC5; #100;
A = 8'h86; B = 8'hC6; #100;
A = 8'h86; B = 8'hC7; #100;
A = 8'h86; B = 8'hC8; #100;
A = 8'h86; B = 8'hC9; #100;
A = 8'h86; B = 8'hCA; #100;
A = 8'h86; B = 8'hCB; #100;
A = 8'h86; B = 8'hCC; #100;
A = 8'h86; B = 8'hCD; #100;
A = 8'h86; B = 8'hCE; #100;
A = 8'h86; B = 8'hCF; #100;
A = 8'h86; B = 8'hD0; #100;
A = 8'h86; B = 8'hD1; #100;
A = 8'h86; B = 8'hD2; #100;
A = 8'h86; B = 8'hD3; #100;
A = 8'h86; B = 8'hD4; #100;
A = 8'h86; B = 8'hD5; #100;
A = 8'h86; B = 8'hD6; #100;
A = 8'h86; B = 8'hD7; #100;
A = 8'h86; B = 8'hD8; #100;
A = 8'h86; B = 8'hD9; #100;
A = 8'h86; B = 8'hDA; #100;
A = 8'h86; B = 8'hDB; #100;
A = 8'h86; B = 8'hDC; #100;
A = 8'h86; B = 8'hDD; #100;
A = 8'h86; B = 8'hDE; #100;
A = 8'h86; B = 8'hDF; #100;
A = 8'h86; B = 8'hE0; #100;
A = 8'h86; B = 8'hE1; #100;
A = 8'h86; B = 8'hE2; #100;
A = 8'h86; B = 8'hE3; #100;
A = 8'h86; B = 8'hE4; #100;
A = 8'h86; B = 8'hE5; #100;
A = 8'h86; B = 8'hE6; #100;
A = 8'h86; B = 8'hE7; #100;
A = 8'h86; B = 8'hE8; #100;
A = 8'h86; B = 8'hE9; #100;
A = 8'h86; B = 8'hEA; #100;
A = 8'h86; B = 8'hEB; #100;
A = 8'h86; B = 8'hEC; #100;
A = 8'h86; B = 8'hED; #100;
A = 8'h86; B = 8'hEE; #100;
A = 8'h86; B = 8'hEF; #100;
A = 8'h86; B = 8'hF0; #100;
A = 8'h86; B = 8'hF1; #100;
A = 8'h86; B = 8'hF2; #100;
A = 8'h86; B = 8'hF3; #100;
A = 8'h86; B = 8'hF4; #100;
A = 8'h86; B = 8'hF5; #100;
A = 8'h86; B = 8'hF6; #100;
A = 8'h86; B = 8'hF7; #100;
A = 8'h86; B = 8'hF8; #100;
A = 8'h86; B = 8'hF9; #100;
A = 8'h86; B = 8'hFA; #100;
A = 8'h86; B = 8'hFB; #100;
A = 8'h86; B = 8'hFC; #100;
A = 8'h86; B = 8'hFD; #100;
A = 8'h86; B = 8'hFE; #100;
A = 8'h86; B = 8'hFF; #100;
A = 8'h87; B = 8'h0; #100;
A = 8'h87; B = 8'h1; #100;
A = 8'h87; B = 8'h2; #100;
A = 8'h87; B = 8'h3; #100;
A = 8'h87; B = 8'h4; #100;
A = 8'h87; B = 8'h5; #100;
A = 8'h87; B = 8'h6; #100;
A = 8'h87; B = 8'h7; #100;
A = 8'h87; B = 8'h8; #100;
A = 8'h87; B = 8'h9; #100;
A = 8'h87; B = 8'hA; #100;
A = 8'h87; B = 8'hB; #100;
A = 8'h87; B = 8'hC; #100;
A = 8'h87; B = 8'hD; #100;
A = 8'h87; B = 8'hE; #100;
A = 8'h87; B = 8'hF; #100;
A = 8'h87; B = 8'h10; #100;
A = 8'h87; B = 8'h11; #100;
A = 8'h87; B = 8'h12; #100;
A = 8'h87; B = 8'h13; #100;
A = 8'h87; B = 8'h14; #100;
A = 8'h87; B = 8'h15; #100;
A = 8'h87; B = 8'h16; #100;
A = 8'h87; B = 8'h17; #100;
A = 8'h87; B = 8'h18; #100;
A = 8'h87; B = 8'h19; #100;
A = 8'h87; B = 8'h1A; #100;
A = 8'h87; B = 8'h1B; #100;
A = 8'h87; B = 8'h1C; #100;
A = 8'h87; B = 8'h1D; #100;
A = 8'h87; B = 8'h1E; #100;
A = 8'h87; B = 8'h1F; #100;
A = 8'h87; B = 8'h20; #100;
A = 8'h87; B = 8'h21; #100;
A = 8'h87; B = 8'h22; #100;
A = 8'h87; B = 8'h23; #100;
A = 8'h87; B = 8'h24; #100;
A = 8'h87; B = 8'h25; #100;
A = 8'h87; B = 8'h26; #100;
A = 8'h87; B = 8'h27; #100;
A = 8'h87; B = 8'h28; #100;
A = 8'h87; B = 8'h29; #100;
A = 8'h87; B = 8'h2A; #100;
A = 8'h87; B = 8'h2B; #100;
A = 8'h87; B = 8'h2C; #100;
A = 8'h87; B = 8'h2D; #100;
A = 8'h87; B = 8'h2E; #100;
A = 8'h87; B = 8'h2F; #100;
A = 8'h87; B = 8'h30; #100;
A = 8'h87; B = 8'h31; #100;
A = 8'h87; B = 8'h32; #100;
A = 8'h87; B = 8'h33; #100;
A = 8'h87; B = 8'h34; #100;
A = 8'h87; B = 8'h35; #100;
A = 8'h87; B = 8'h36; #100;
A = 8'h87; B = 8'h37; #100;
A = 8'h87; B = 8'h38; #100;
A = 8'h87; B = 8'h39; #100;
A = 8'h87; B = 8'h3A; #100;
A = 8'h87; B = 8'h3B; #100;
A = 8'h87; B = 8'h3C; #100;
A = 8'h87; B = 8'h3D; #100;
A = 8'h87; B = 8'h3E; #100;
A = 8'h87; B = 8'h3F; #100;
A = 8'h87; B = 8'h40; #100;
A = 8'h87; B = 8'h41; #100;
A = 8'h87; B = 8'h42; #100;
A = 8'h87; B = 8'h43; #100;
A = 8'h87; B = 8'h44; #100;
A = 8'h87; B = 8'h45; #100;
A = 8'h87; B = 8'h46; #100;
A = 8'h87; B = 8'h47; #100;
A = 8'h87; B = 8'h48; #100;
A = 8'h87; B = 8'h49; #100;
A = 8'h87; B = 8'h4A; #100;
A = 8'h87; B = 8'h4B; #100;
A = 8'h87; B = 8'h4C; #100;
A = 8'h87; B = 8'h4D; #100;
A = 8'h87; B = 8'h4E; #100;
A = 8'h87; B = 8'h4F; #100;
A = 8'h87; B = 8'h50; #100;
A = 8'h87; B = 8'h51; #100;
A = 8'h87; B = 8'h52; #100;
A = 8'h87; B = 8'h53; #100;
A = 8'h87; B = 8'h54; #100;
A = 8'h87; B = 8'h55; #100;
A = 8'h87; B = 8'h56; #100;
A = 8'h87; B = 8'h57; #100;
A = 8'h87; B = 8'h58; #100;
A = 8'h87; B = 8'h59; #100;
A = 8'h87; B = 8'h5A; #100;
A = 8'h87; B = 8'h5B; #100;
A = 8'h87; B = 8'h5C; #100;
A = 8'h87; B = 8'h5D; #100;
A = 8'h87; B = 8'h5E; #100;
A = 8'h87; B = 8'h5F; #100;
A = 8'h87; B = 8'h60; #100;
A = 8'h87; B = 8'h61; #100;
A = 8'h87; B = 8'h62; #100;
A = 8'h87; B = 8'h63; #100;
A = 8'h87; B = 8'h64; #100;
A = 8'h87; B = 8'h65; #100;
A = 8'h87; B = 8'h66; #100;
A = 8'h87; B = 8'h67; #100;
A = 8'h87; B = 8'h68; #100;
A = 8'h87; B = 8'h69; #100;
A = 8'h87; B = 8'h6A; #100;
A = 8'h87; B = 8'h6B; #100;
A = 8'h87; B = 8'h6C; #100;
A = 8'h87; B = 8'h6D; #100;
A = 8'h87; B = 8'h6E; #100;
A = 8'h87; B = 8'h6F; #100;
A = 8'h87; B = 8'h70; #100;
A = 8'h87; B = 8'h71; #100;
A = 8'h87; B = 8'h72; #100;
A = 8'h87; B = 8'h73; #100;
A = 8'h87; B = 8'h74; #100;
A = 8'h87; B = 8'h75; #100;
A = 8'h87; B = 8'h76; #100;
A = 8'h87; B = 8'h77; #100;
A = 8'h87; B = 8'h78; #100;
A = 8'h87; B = 8'h79; #100;
A = 8'h87; B = 8'h7A; #100;
A = 8'h87; B = 8'h7B; #100;
A = 8'h87; B = 8'h7C; #100;
A = 8'h87; B = 8'h7D; #100;
A = 8'h87; B = 8'h7E; #100;
A = 8'h87; B = 8'h7F; #100;
A = 8'h87; B = 8'h80; #100;
A = 8'h87; B = 8'h81; #100;
A = 8'h87; B = 8'h82; #100;
A = 8'h87; B = 8'h83; #100;
A = 8'h87; B = 8'h84; #100;
A = 8'h87; B = 8'h85; #100;
A = 8'h87; B = 8'h86; #100;
A = 8'h87; B = 8'h87; #100;
A = 8'h87; B = 8'h88; #100;
A = 8'h87; B = 8'h89; #100;
A = 8'h87; B = 8'h8A; #100;
A = 8'h87; B = 8'h8B; #100;
A = 8'h87; B = 8'h8C; #100;
A = 8'h87; B = 8'h8D; #100;
A = 8'h87; B = 8'h8E; #100;
A = 8'h87; B = 8'h8F; #100;
A = 8'h87; B = 8'h90; #100;
A = 8'h87; B = 8'h91; #100;
A = 8'h87; B = 8'h92; #100;
A = 8'h87; B = 8'h93; #100;
A = 8'h87; B = 8'h94; #100;
A = 8'h87; B = 8'h95; #100;
A = 8'h87; B = 8'h96; #100;
A = 8'h87; B = 8'h97; #100;
A = 8'h87; B = 8'h98; #100;
A = 8'h87; B = 8'h99; #100;
A = 8'h87; B = 8'h9A; #100;
A = 8'h87; B = 8'h9B; #100;
A = 8'h87; B = 8'h9C; #100;
A = 8'h87; B = 8'h9D; #100;
A = 8'h87; B = 8'h9E; #100;
A = 8'h87; B = 8'h9F; #100;
A = 8'h87; B = 8'hA0; #100;
A = 8'h87; B = 8'hA1; #100;
A = 8'h87; B = 8'hA2; #100;
A = 8'h87; B = 8'hA3; #100;
A = 8'h87; B = 8'hA4; #100;
A = 8'h87; B = 8'hA5; #100;
A = 8'h87; B = 8'hA6; #100;
A = 8'h87; B = 8'hA7; #100;
A = 8'h87; B = 8'hA8; #100;
A = 8'h87; B = 8'hA9; #100;
A = 8'h87; B = 8'hAA; #100;
A = 8'h87; B = 8'hAB; #100;
A = 8'h87; B = 8'hAC; #100;
A = 8'h87; B = 8'hAD; #100;
A = 8'h87; B = 8'hAE; #100;
A = 8'h87; B = 8'hAF; #100;
A = 8'h87; B = 8'hB0; #100;
A = 8'h87; B = 8'hB1; #100;
A = 8'h87; B = 8'hB2; #100;
A = 8'h87; B = 8'hB3; #100;
A = 8'h87; B = 8'hB4; #100;
A = 8'h87; B = 8'hB5; #100;
A = 8'h87; B = 8'hB6; #100;
A = 8'h87; B = 8'hB7; #100;
A = 8'h87; B = 8'hB8; #100;
A = 8'h87; B = 8'hB9; #100;
A = 8'h87; B = 8'hBA; #100;
A = 8'h87; B = 8'hBB; #100;
A = 8'h87; B = 8'hBC; #100;
A = 8'h87; B = 8'hBD; #100;
A = 8'h87; B = 8'hBE; #100;
A = 8'h87; B = 8'hBF; #100;
A = 8'h87; B = 8'hC0; #100;
A = 8'h87; B = 8'hC1; #100;
A = 8'h87; B = 8'hC2; #100;
A = 8'h87; B = 8'hC3; #100;
A = 8'h87; B = 8'hC4; #100;
A = 8'h87; B = 8'hC5; #100;
A = 8'h87; B = 8'hC6; #100;
A = 8'h87; B = 8'hC7; #100;
A = 8'h87; B = 8'hC8; #100;
A = 8'h87; B = 8'hC9; #100;
A = 8'h87; B = 8'hCA; #100;
A = 8'h87; B = 8'hCB; #100;
A = 8'h87; B = 8'hCC; #100;
A = 8'h87; B = 8'hCD; #100;
A = 8'h87; B = 8'hCE; #100;
A = 8'h87; B = 8'hCF; #100;
A = 8'h87; B = 8'hD0; #100;
A = 8'h87; B = 8'hD1; #100;
A = 8'h87; B = 8'hD2; #100;
A = 8'h87; B = 8'hD3; #100;
A = 8'h87; B = 8'hD4; #100;
A = 8'h87; B = 8'hD5; #100;
A = 8'h87; B = 8'hD6; #100;
A = 8'h87; B = 8'hD7; #100;
A = 8'h87; B = 8'hD8; #100;
A = 8'h87; B = 8'hD9; #100;
A = 8'h87; B = 8'hDA; #100;
A = 8'h87; B = 8'hDB; #100;
A = 8'h87; B = 8'hDC; #100;
A = 8'h87; B = 8'hDD; #100;
A = 8'h87; B = 8'hDE; #100;
A = 8'h87; B = 8'hDF; #100;
A = 8'h87; B = 8'hE0; #100;
A = 8'h87; B = 8'hE1; #100;
A = 8'h87; B = 8'hE2; #100;
A = 8'h87; B = 8'hE3; #100;
A = 8'h87; B = 8'hE4; #100;
A = 8'h87; B = 8'hE5; #100;
A = 8'h87; B = 8'hE6; #100;
A = 8'h87; B = 8'hE7; #100;
A = 8'h87; B = 8'hE8; #100;
A = 8'h87; B = 8'hE9; #100;
A = 8'h87; B = 8'hEA; #100;
A = 8'h87; B = 8'hEB; #100;
A = 8'h87; B = 8'hEC; #100;
A = 8'h87; B = 8'hED; #100;
A = 8'h87; B = 8'hEE; #100;
A = 8'h87; B = 8'hEF; #100;
A = 8'h87; B = 8'hF0; #100;
A = 8'h87; B = 8'hF1; #100;
A = 8'h87; B = 8'hF2; #100;
A = 8'h87; B = 8'hF3; #100;
A = 8'h87; B = 8'hF4; #100;
A = 8'h87; B = 8'hF5; #100;
A = 8'h87; B = 8'hF6; #100;
A = 8'h87; B = 8'hF7; #100;
A = 8'h87; B = 8'hF8; #100;
A = 8'h87; B = 8'hF9; #100;
A = 8'h87; B = 8'hFA; #100;
A = 8'h87; B = 8'hFB; #100;
A = 8'h87; B = 8'hFC; #100;
A = 8'h87; B = 8'hFD; #100;
A = 8'h87; B = 8'hFE; #100;
A = 8'h87; B = 8'hFF; #100;
A = 8'h88; B = 8'h0; #100;
A = 8'h88; B = 8'h1; #100;
A = 8'h88; B = 8'h2; #100;
A = 8'h88; B = 8'h3; #100;
A = 8'h88; B = 8'h4; #100;
A = 8'h88; B = 8'h5; #100;
A = 8'h88; B = 8'h6; #100;
A = 8'h88; B = 8'h7; #100;
A = 8'h88; B = 8'h8; #100;
A = 8'h88; B = 8'h9; #100;
A = 8'h88; B = 8'hA; #100;
A = 8'h88; B = 8'hB; #100;
A = 8'h88; B = 8'hC; #100;
A = 8'h88; B = 8'hD; #100;
A = 8'h88; B = 8'hE; #100;
A = 8'h88; B = 8'hF; #100;
A = 8'h88; B = 8'h10; #100;
A = 8'h88; B = 8'h11; #100;
A = 8'h88; B = 8'h12; #100;
A = 8'h88; B = 8'h13; #100;
A = 8'h88; B = 8'h14; #100;
A = 8'h88; B = 8'h15; #100;
A = 8'h88; B = 8'h16; #100;
A = 8'h88; B = 8'h17; #100;
A = 8'h88; B = 8'h18; #100;
A = 8'h88; B = 8'h19; #100;
A = 8'h88; B = 8'h1A; #100;
A = 8'h88; B = 8'h1B; #100;
A = 8'h88; B = 8'h1C; #100;
A = 8'h88; B = 8'h1D; #100;
A = 8'h88; B = 8'h1E; #100;
A = 8'h88; B = 8'h1F; #100;
A = 8'h88; B = 8'h20; #100;
A = 8'h88; B = 8'h21; #100;
A = 8'h88; B = 8'h22; #100;
A = 8'h88; B = 8'h23; #100;
A = 8'h88; B = 8'h24; #100;
A = 8'h88; B = 8'h25; #100;
A = 8'h88; B = 8'h26; #100;
A = 8'h88; B = 8'h27; #100;
A = 8'h88; B = 8'h28; #100;
A = 8'h88; B = 8'h29; #100;
A = 8'h88; B = 8'h2A; #100;
A = 8'h88; B = 8'h2B; #100;
A = 8'h88; B = 8'h2C; #100;
A = 8'h88; B = 8'h2D; #100;
A = 8'h88; B = 8'h2E; #100;
A = 8'h88; B = 8'h2F; #100;
A = 8'h88; B = 8'h30; #100;
A = 8'h88; B = 8'h31; #100;
A = 8'h88; B = 8'h32; #100;
A = 8'h88; B = 8'h33; #100;
A = 8'h88; B = 8'h34; #100;
A = 8'h88; B = 8'h35; #100;
A = 8'h88; B = 8'h36; #100;
A = 8'h88; B = 8'h37; #100;
A = 8'h88; B = 8'h38; #100;
A = 8'h88; B = 8'h39; #100;
A = 8'h88; B = 8'h3A; #100;
A = 8'h88; B = 8'h3B; #100;
A = 8'h88; B = 8'h3C; #100;
A = 8'h88; B = 8'h3D; #100;
A = 8'h88; B = 8'h3E; #100;
A = 8'h88; B = 8'h3F; #100;
A = 8'h88; B = 8'h40; #100;
A = 8'h88; B = 8'h41; #100;
A = 8'h88; B = 8'h42; #100;
A = 8'h88; B = 8'h43; #100;
A = 8'h88; B = 8'h44; #100;
A = 8'h88; B = 8'h45; #100;
A = 8'h88; B = 8'h46; #100;
A = 8'h88; B = 8'h47; #100;
A = 8'h88; B = 8'h48; #100;
A = 8'h88; B = 8'h49; #100;
A = 8'h88; B = 8'h4A; #100;
A = 8'h88; B = 8'h4B; #100;
A = 8'h88; B = 8'h4C; #100;
A = 8'h88; B = 8'h4D; #100;
A = 8'h88; B = 8'h4E; #100;
A = 8'h88; B = 8'h4F; #100;
A = 8'h88; B = 8'h50; #100;
A = 8'h88; B = 8'h51; #100;
A = 8'h88; B = 8'h52; #100;
A = 8'h88; B = 8'h53; #100;
A = 8'h88; B = 8'h54; #100;
A = 8'h88; B = 8'h55; #100;
A = 8'h88; B = 8'h56; #100;
A = 8'h88; B = 8'h57; #100;
A = 8'h88; B = 8'h58; #100;
A = 8'h88; B = 8'h59; #100;
A = 8'h88; B = 8'h5A; #100;
A = 8'h88; B = 8'h5B; #100;
A = 8'h88; B = 8'h5C; #100;
A = 8'h88; B = 8'h5D; #100;
A = 8'h88; B = 8'h5E; #100;
A = 8'h88; B = 8'h5F; #100;
A = 8'h88; B = 8'h60; #100;
A = 8'h88; B = 8'h61; #100;
A = 8'h88; B = 8'h62; #100;
A = 8'h88; B = 8'h63; #100;
A = 8'h88; B = 8'h64; #100;
A = 8'h88; B = 8'h65; #100;
A = 8'h88; B = 8'h66; #100;
A = 8'h88; B = 8'h67; #100;
A = 8'h88; B = 8'h68; #100;
A = 8'h88; B = 8'h69; #100;
A = 8'h88; B = 8'h6A; #100;
A = 8'h88; B = 8'h6B; #100;
A = 8'h88; B = 8'h6C; #100;
A = 8'h88; B = 8'h6D; #100;
A = 8'h88; B = 8'h6E; #100;
A = 8'h88; B = 8'h6F; #100;
A = 8'h88; B = 8'h70; #100;
A = 8'h88; B = 8'h71; #100;
A = 8'h88; B = 8'h72; #100;
A = 8'h88; B = 8'h73; #100;
A = 8'h88; B = 8'h74; #100;
A = 8'h88; B = 8'h75; #100;
A = 8'h88; B = 8'h76; #100;
A = 8'h88; B = 8'h77; #100;
A = 8'h88; B = 8'h78; #100;
A = 8'h88; B = 8'h79; #100;
A = 8'h88; B = 8'h7A; #100;
A = 8'h88; B = 8'h7B; #100;
A = 8'h88; B = 8'h7C; #100;
A = 8'h88; B = 8'h7D; #100;
A = 8'h88; B = 8'h7E; #100;
A = 8'h88; B = 8'h7F; #100;
A = 8'h88; B = 8'h80; #100;
A = 8'h88; B = 8'h81; #100;
A = 8'h88; B = 8'h82; #100;
A = 8'h88; B = 8'h83; #100;
A = 8'h88; B = 8'h84; #100;
A = 8'h88; B = 8'h85; #100;
A = 8'h88; B = 8'h86; #100;
A = 8'h88; B = 8'h87; #100;
A = 8'h88; B = 8'h88; #100;
A = 8'h88; B = 8'h89; #100;
A = 8'h88; B = 8'h8A; #100;
A = 8'h88; B = 8'h8B; #100;
A = 8'h88; B = 8'h8C; #100;
A = 8'h88; B = 8'h8D; #100;
A = 8'h88; B = 8'h8E; #100;
A = 8'h88; B = 8'h8F; #100;
A = 8'h88; B = 8'h90; #100;
A = 8'h88; B = 8'h91; #100;
A = 8'h88; B = 8'h92; #100;
A = 8'h88; B = 8'h93; #100;
A = 8'h88; B = 8'h94; #100;
A = 8'h88; B = 8'h95; #100;
A = 8'h88; B = 8'h96; #100;
A = 8'h88; B = 8'h97; #100;
A = 8'h88; B = 8'h98; #100;
A = 8'h88; B = 8'h99; #100;
A = 8'h88; B = 8'h9A; #100;
A = 8'h88; B = 8'h9B; #100;
A = 8'h88; B = 8'h9C; #100;
A = 8'h88; B = 8'h9D; #100;
A = 8'h88; B = 8'h9E; #100;
A = 8'h88; B = 8'h9F; #100;
A = 8'h88; B = 8'hA0; #100;
A = 8'h88; B = 8'hA1; #100;
A = 8'h88; B = 8'hA2; #100;
A = 8'h88; B = 8'hA3; #100;
A = 8'h88; B = 8'hA4; #100;
A = 8'h88; B = 8'hA5; #100;
A = 8'h88; B = 8'hA6; #100;
A = 8'h88; B = 8'hA7; #100;
A = 8'h88; B = 8'hA8; #100;
A = 8'h88; B = 8'hA9; #100;
A = 8'h88; B = 8'hAA; #100;
A = 8'h88; B = 8'hAB; #100;
A = 8'h88; B = 8'hAC; #100;
A = 8'h88; B = 8'hAD; #100;
A = 8'h88; B = 8'hAE; #100;
A = 8'h88; B = 8'hAF; #100;
A = 8'h88; B = 8'hB0; #100;
A = 8'h88; B = 8'hB1; #100;
A = 8'h88; B = 8'hB2; #100;
A = 8'h88; B = 8'hB3; #100;
A = 8'h88; B = 8'hB4; #100;
A = 8'h88; B = 8'hB5; #100;
A = 8'h88; B = 8'hB6; #100;
A = 8'h88; B = 8'hB7; #100;
A = 8'h88; B = 8'hB8; #100;
A = 8'h88; B = 8'hB9; #100;
A = 8'h88; B = 8'hBA; #100;
A = 8'h88; B = 8'hBB; #100;
A = 8'h88; B = 8'hBC; #100;
A = 8'h88; B = 8'hBD; #100;
A = 8'h88; B = 8'hBE; #100;
A = 8'h88; B = 8'hBF; #100;
A = 8'h88; B = 8'hC0; #100;
A = 8'h88; B = 8'hC1; #100;
A = 8'h88; B = 8'hC2; #100;
A = 8'h88; B = 8'hC3; #100;
A = 8'h88; B = 8'hC4; #100;
A = 8'h88; B = 8'hC5; #100;
A = 8'h88; B = 8'hC6; #100;
A = 8'h88; B = 8'hC7; #100;
A = 8'h88; B = 8'hC8; #100;
A = 8'h88; B = 8'hC9; #100;
A = 8'h88; B = 8'hCA; #100;
A = 8'h88; B = 8'hCB; #100;
A = 8'h88; B = 8'hCC; #100;
A = 8'h88; B = 8'hCD; #100;
A = 8'h88; B = 8'hCE; #100;
A = 8'h88; B = 8'hCF; #100;
A = 8'h88; B = 8'hD0; #100;
A = 8'h88; B = 8'hD1; #100;
A = 8'h88; B = 8'hD2; #100;
A = 8'h88; B = 8'hD3; #100;
A = 8'h88; B = 8'hD4; #100;
A = 8'h88; B = 8'hD5; #100;
A = 8'h88; B = 8'hD6; #100;
A = 8'h88; B = 8'hD7; #100;
A = 8'h88; B = 8'hD8; #100;
A = 8'h88; B = 8'hD9; #100;
A = 8'h88; B = 8'hDA; #100;
A = 8'h88; B = 8'hDB; #100;
A = 8'h88; B = 8'hDC; #100;
A = 8'h88; B = 8'hDD; #100;
A = 8'h88; B = 8'hDE; #100;
A = 8'h88; B = 8'hDF; #100;
A = 8'h88; B = 8'hE0; #100;
A = 8'h88; B = 8'hE1; #100;
A = 8'h88; B = 8'hE2; #100;
A = 8'h88; B = 8'hE3; #100;
A = 8'h88; B = 8'hE4; #100;
A = 8'h88; B = 8'hE5; #100;
A = 8'h88; B = 8'hE6; #100;
A = 8'h88; B = 8'hE7; #100;
A = 8'h88; B = 8'hE8; #100;
A = 8'h88; B = 8'hE9; #100;
A = 8'h88; B = 8'hEA; #100;
A = 8'h88; B = 8'hEB; #100;
A = 8'h88; B = 8'hEC; #100;
A = 8'h88; B = 8'hED; #100;
A = 8'h88; B = 8'hEE; #100;
A = 8'h88; B = 8'hEF; #100;
A = 8'h88; B = 8'hF0; #100;
A = 8'h88; B = 8'hF1; #100;
A = 8'h88; B = 8'hF2; #100;
A = 8'h88; B = 8'hF3; #100;
A = 8'h88; B = 8'hF4; #100;
A = 8'h88; B = 8'hF5; #100;
A = 8'h88; B = 8'hF6; #100;
A = 8'h88; B = 8'hF7; #100;
A = 8'h88; B = 8'hF8; #100;
A = 8'h88; B = 8'hF9; #100;
A = 8'h88; B = 8'hFA; #100;
A = 8'h88; B = 8'hFB; #100;
A = 8'h88; B = 8'hFC; #100;
A = 8'h88; B = 8'hFD; #100;
A = 8'h88; B = 8'hFE; #100;
A = 8'h88; B = 8'hFF; #100;
A = 8'h89; B = 8'h0; #100;
A = 8'h89; B = 8'h1; #100;
A = 8'h89; B = 8'h2; #100;
A = 8'h89; B = 8'h3; #100;
A = 8'h89; B = 8'h4; #100;
A = 8'h89; B = 8'h5; #100;
A = 8'h89; B = 8'h6; #100;
A = 8'h89; B = 8'h7; #100;
A = 8'h89; B = 8'h8; #100;
A = 8'h89; B = 8'h9; #100;
A = 8'h89; B = 8'hA; #100;
A = 8'h89; B = 8'hB; #100;
A = 8'h89; B = 8'hC; #100;
A = 8'h89; B = 8'hD; #100;
A = 8'h89; B = 8'hE; #100;
A = 8'h89; B = 8'hF; #100;
A = 8'h89; B = 8'h10; #100;
A = 8'h89; B = 8'h11; #100;
A = 8'h89; B = 8'h12; #100;
A = 8'h89; B = 8'h13; #100;
A = 8'h89; B = 8'h14; #100;
A = 8'h89; B = 8'h15; #100;
A = 8'h89; B = 8'h16; #100;
A = 8'h89; B = 8'h17; #100;
A = 8'h89; B = 8'h18; #100;
A = 8'h89; B = 8'h19; #100;
A = 8'h89; B = 8'h1A; #100;
A = 8'h89; B = 8'h1B; #100;
A = 8'h89; B = 8'h1C; #100;
A = 8'h89; B = 8'h1D; #100;
A = 8'h89; B = 8'h1E; #100;
A = 8'h89; B = 8'h1F; #100;
A = 8'h89; B = 8'h20; #100;
A = 8'h89; B = 8'h21; #100;
A = 8'h89; B = 8'h22; #100;
A = 8'h89; B = 8'h23; #100;
A = 8'h89; B = 8'h24; #100;
A = 8'h89; B = 8'h25; #100;
A = 8'h89; B = 8'h26; #100;
A = 8'h89; B = 8'h27; #100;
A = 8'h89; B = 8'h28; #100;
A = 8'h89; B = 8'h29; #100;
A = 8'h89; B = 8'h2A; #100;
A = 8'h89; B = 8'h2B; #100;
A = 8'h89; B = 8'h2C; #100;
A = 8'h89; B = 8'h2D; #100;
A = 8'h89; B = 8'h2E; #100;
A = 8'h89; B = 8'h2F; #100;
A = 8'h89; B = 8'h30; #100;
A = 8'h89; B = 8'h31; #100;
A = 8'h89; B = 8'h32; #100;
A = 8'h89; B = 8'h33; #100;
A = 8'h89; B = 8'h34; #100;
A = 8'h89; B = 8'h35; #100;
A = 8'h89; B = 8'h36; #100;
A = 8'h89; B = 8'h37; #100;
A = 8'h89; B = 8'h38; #100;
A = 8'h89; B = 8'h39; #100;
A = 8'h89; B = 8'h3A; #100;
A = 8'h89; B = 8'h3B; #100;
A = 8'h89; B = 8'h3C; #100;
A = 8'h89; B = 8'h3D; #100;
A = 8'h89; B = 8'h3E; #100;
A = 8'h89; B = 8'h3F; #100;
A = 8'h89; B = 8'h40; #100;
A = 8'h89; B = 8'h41; #100;
A = 8'h89; B = 8'h42; #100;
A = 8'h89; B = 8'h43; #100;
A = 8'h89; B = 8'h44; #100;
A = 8'h89; B = 8'h45; #100;
A = 8'h89; B = 8'h46; #100;
A = 8'h89; B = 8'h47; #100;
A = 8'h89; B = 8'h48; #100;
A = 8'h89; B = 8'h49; #100;
A = 8'h89; B = 8'h4A; #100;
A = 8'h89; B = 8'h4B; #100;
A = 8'h89; B = 8'h4C; #100;
A = 8'h89; B = 8'h4D; #100;
A = 8'h89; B = 8'h4E; #100;
A = 8'h89; B = 8'h4F; #100;
A = 8'h89; B = 8'h50; #100;
A = 8'h89; B = 8'h51; #100;
A = 8'h89; B = 8'h52; #100;
A = 8'h89; B = 8'h53; #100;
A = 8'h89; B = 8'h54; #100;
A = 8'h89; B = 8'h55; #100;
A = 8'h89; B = 8'h56; #100;
A = 8'h89; B = 8'h57; #100;
A = 8'h89; B = 8'h58; #100;
A = 8'h89; B = 8'h59; #100;
A = 8'h89; B = 8'h5A; #100;
A = 8'h89; B = 8'h5B; #100;
A = 8'h89; B = 8'h5C; #100;
A = 8'h89; B = 8'h5D; #100;
A = 8'h89; B = 8'h5E; #100;
A = 8'h89; B = 8'h5F; #100;
A = 8'h89; B = 8'h60; #100;
A = 8'h89; B = 8'h61; #100;
A = 8'h89; B = 8'h62; #100;
A = 8'h89; B = 8'h63; #100;
A = 8'h89; B = 8'h64; #100;
A = 8'h89; B = 8'h65; #100;
A = 8'h89; B = 8'h66; #100;
A = 8'h89; B = 8'h67; #100;
A = 8'h89; B = 8'h68; #100;
A = 8'h89; B = 8'h69; #100;
A = 8'h89; B = 8'h6A; #100;
A = 8'h89; B = 8'h6B; #100;
A = 8'h89; B = 8'h6C; #100;
A = 8'h89; B = 8'h6D; #100;
A = 8'h89; B = 8'h6E; #100;
A = 8'h89; B = 8'h6F; #100;
A = 8'h89; B = 8'h70; #100;
A = 8'h89; B = 8'h71; #100;
A = 8'h89; B = 8'h72; #100;
A = 8'h89; B = 8'h73; #100;
A = 8'h89; B = 8'h74; #100;
A = 8'h89; B = 8'h75; #100;
A = 8'h89; B = 8'h76; #100;
A = 8'h89; B = 8'h77; #100;
A = 8'h89; B = 8'h78; #100;
A = 8'h89; B = 8'h79; #100;
A = 8'h89; B = 8'h7A; #100;
A = 8'h89; B = 8'h7B; #100;
A = 8'h89; B = 8'h7C; #100;
A = 8'h89; B = 8'h7D; #100;
A = 8'h89; B = 8'h7E; #100;
A = 8'h89; B = 8'h7F; #100;
A = 8'h89; B = 8'h80; #100;
A = 8'h89; B = 8'h81; #100;
A = 8'h89; B = 8'h82; #100;
A = 8'h89; B = 8'h83; #100;
A = 8'h89; B = 8'h84; #100;
A = 8'h89; B = 8'h85; #100;
A = 8'h89; B = 8'h86; #100;
A = 8'h89; B = 8'h87; #100;
A = 8'h89; B = 8'h88; #100;
A = 8'h89; B = 8'h89; #100;
A = 8'h89; B = 8'h8A; #100;
A = 8'h89; B = 8'h8B; #100;
A = 8'h89; B = 8'h8C; #100;
A = 8'h89; B = 8'h8D; #100;
A = 8'h89; B = 8'h8E; #100;
A = 8'h89; B = 8'h8F; #100;
A = 8'h89; B = 8'h90; #100;
A = 8'h89; B = 8'h91; #100;
A = 8'h89; B = 8'h92; #100;
A = 8'h89; B = 8'h93; #100;
A = 8'h89; B = 8'h94; #100;
A = 8'h89; B = 8'h95; #100;
A = 8'h89; B = 8'h96; #100;
A = 8'h89; B = 8'h97; #100;
A = 8'h89; B = 8'h98; #100;
A = 8'h89; B = 8'h99; #100;
A = 8'h89; B = 8'h9A; #100;
A = 8'h89; B = 8'h9B; #100;
A = 8'h89; B = 8'h9C; #100;
A = 8'h89; B = 8'h9D; #100;
A = 8'h89; B = 8'h9E; #100;
A = 8'h89; B = 8'h9F; #100;
A = 8'h89; B = 8'hA0; #100;
A = 8'h89; B = 8'hA1; #100;
A = 8'h89; B = 8'hA2; #100;
A = 8'h89; B = 8'hA3; #100;
A = 8'h89; B = 8'hA4; #100;
A = 8'h89; B = 8'hA5; #100;
A = 8'h89; B = 8'hA6; #100;
A = 8'h89; B = 8'hA7; #100;
A = 8'h89; B = 8'hA8; #100;
A = 8'h89; B = 8'hA9; #100;
A = 8'h89; B = 8'hAA; #100;
A = 8'h89; B = 8'hAB; #100;
A = 8'h89; B = 8'hAC; #100;
A = 8'h89; B = 8'hAD; #100;
A = 8'h89; B = 8'hAE; #100;
A = 8'h89; B = 8'hAF; #100;
A = 8'h89; B = 8'hB0; #100;
A = 8'h89; B = 8'hB1; #100;
A = 8'h89; B = 8'hB2; #100;
A = 8'h89; B = 8'hB3; #100;
A = 8'h89; B = 8'hB4; #100;
A = 8'h89; B = 8'hB5; #100;
A = 8'h89; B = 8'hB6; #100;
A = 8'h89; B = 8'hB7; #100;
A = 8'h89; B = 8'hB8; #100;
A = 8'h89; B = 8'hB9; #100;
A = 8'h89; B = 8'hBA; #100;
A = 8'h89; B = 8'hBB; #100;
A = 8'h89; B = 8'hBC; #100;
A = 8'h89; B = 8'hBD; #100;
A = 8'h89; B = 8'hBE; #100;
A = 8'h89; B = 8'hBF; #100;
A = 8'h89; B = 8'hC0; #100;
A = 8'h89; B = 8'hC1; #100;
A = 8'h89; B = 8'hC2; #100;
A = 8'h89; B = 8'hC3; #100;
A = 8'h89; B = 8'hC4; #100;
A = 8'h89; B = 8'hC5; #100;
A = 8'h89; B = 8'hC6; #100;
A = 8'h89; B = 8'hC7; #100;
A = 8'h89; B = 8'hC8; #100;
A = 8'h89; B = 8'hC9; #100;
A = 8'h89; B = 8'hCA; #100;
A = 8'h89; B = 8'hCB; #100;
A = 8'h89; B = 8'hCC; #100;
A = 8'h89; B = 8'hCD; #100;
A = 8'h89; B = 8'hCE; #100;
A = 8'h89; B = 8'hCF; #100;
A = 8'h89; B = 8'hD0; #100;
A = 8'h89; B = 8'hD1; #100;
A = 8'h89; B = 8'hD2; #100;
A = 8'h89; B = 8'hD3; #100;
A = 8'h89; B = 8'hD4; #100;
A = 8'h89; B = 8'hD5; #100;
A = 8'h89; B = 8'hD6; #100;
A = 8'h89; B = 8'hD7; #100;
A = 8'h89; B = 8'hD8; #100;
A = 8'h89; B = 8'hD9; #100;
A = 8'h89; B = 8'hDA; #100;
A = 8'h89; B = 8'hDB; #100;
A = 8'h89; B = 8'hDC; #100;
A = 8'h89; B = 8'hDD; #100;
A = 8'h89; B = 8'hDE; #100;
A = 8'h89; B = 8'hDF; #100;
A = 8'h89; B = 8'hE0; #100;
A = 8'h89; B = 8'hE1; #100;
A = 8'h89; B = 8'hE2; #100;
A = 8'h89; B = 8'hE3; #100;
A = 8'h89; B = 8'hE4; #100;
A = 8'h89; B = 8'hE5; #100;
A = 8'h89; B = 8'hE6; #100;
A = 8'h89; B = 8'hE7; #100;
A = 8'h89; B = 8'hE8; #100;
A = 8'h89; B = 8'hE9; #100;
A = 8'h89; B = 8'hEA; #100;
A = 8'h89; B = 8'hEB; #100;
A = 8'h89; B = 8'hEC; #100;
A = 8'h89; B = 8'hED; #100;
A = 8'h89; B = 8'hEE; #100;
A = 8'h89; B = 8'hEF; #100;
A = 8'h89; B = 8'hF0; #100;
A = 8'h89; B = 8'hF1; #100;
A = 8'h89; B = 8'hF2; #100;
A = 8'h89; B = 8'hF3; #100;
A = 8'h89; B = 8'hF4; #100;
A = 8'h89; B = 8'hF5; #100;
A = 8'h89; B = 8'hF6; #100;
A = 8'h89; B = 8'hF7; #100;
A = 8'h89; B = 8'hF8; #100;
A = 8'h89; B = 8'hF9; #100;
A = 8'h89; B = 8'hFA; #100;
A = 8'h89; B = 8'hFB; #100;
A = 8'h89; B = 8'hFC; #100;
A = 8'h89; B = 8'hFD; #100;
A = 8'h89; B = 8'hFE; #100;
A = 8'h89; B = 8'hFF; #100;
A = 8'h8A; B = 8'h0; #100;
A = 8'h8A; B = 8'h1; #100;
A = 8'h8A; B = 8'h2; #100;
A = 8'h8A; B = 8'h3; #100;
A = 8'h8A; B = 8'h4; #100;
A = 8'h8A; B = 8'h5; #100;
A = 8'h8A; B = 8'h6; #100;
A = 8'h8A; B = 8'h7; #100;
A = 8'h8A; B = 8'h8; #100;
A = 8'h8A; B = 8'h9; #100;
A = 8'h8A; B = 8'hA; #100;
A = 8'h8A; B = 8'hB; #100;
A = 8'h8A; B = 8'hC; #100;
A = 8'h8A; B = 8'hD; #100;
A = 8'h8A; B = 8'hE; #100;
A = 8'h8A; B = 8'hF; #100;
A = 8'h8A; B = 8'h10; #100;
A = 8'h8A; B = 8'h11; #100;
A = 8'h8A; B = 8'h12; #100;
A = 8'h8A; B = 8'h13; #100;
A = 8'h8A; B = 8'h14; #100;
A = 8'h8A; B = 8'h15; #100;
A = 8'h8A; B = 8'h16; #100;
A = 8'h8A; B = 8'h17; #100;
A = 8'h8A; B = 8'h18; #100;
A = 8'h8A; B = 8'h19; #100;
A = 8'h8A; B = 8'h1A; #100;
A = 8'h8A; B = 8'h1B; #100;
A = 8'h8A; B = 8'h1C; #100;
A = 8'h8A; B = 8'h1D; #100;
A = 8'h8A; B = 8'h1E; #100;
A = 8'h8A; B = 8'h1F; #100;
A = 8'h8A; B = 8'h20; #100;
A = 8'h8A; B = 8'h21; #100;
A = 8'h8A; B = 8'h22; #100;
A = 8'h8A; B = 8'h23; #100;
A = 8'h8A; B = 8'h24; #100;
A = 8'h8A; B = 8'h25; #100;
A = 8'h8A; B = 8'h26; #100;
A = 8'h8A; B = 8'h27; #100;
A = 8'h8A; B = 8'h28; #100;
A = 8'h8A; B = 8'h29; #100;
A = 8'h8A; B = 8'h2A; #100;
A = 8'h8A; B = 8'h2B; #100;
A = 8'h8A; B = 8'h2C; #100;
A = 8'h8A; B = 8'h2D; #100;
A = 8'h8A; B = 8'h2E; #100;
A = 8'h8A; B = 8'h2F; #100;
A = 8'h8A; B = 8'h30; #100;
A = 8'h8A; B = 8'h31; #100;
A = 8'h8A; B = 8'h32; #100;
A = 8'h8A; B = 8'h33; #100;
A = 8'h8A; B = 8'h34; #100;
A = 8'h8A; B = 8'h35; #100;
A = 8'h8A; B = 8'h36; #100;
A = 8'h8A; B = 8'h37; #100;
A = 8'h8A; B = 8'h38; #100;
A = 8'h8A; B = 8'h39; #100;
A = 8'h8A; B = 8'h3A; #100;
A = 8'h8A; B = 8'h3B; #100;
A = 8'h8A; B = 8'h3C; #100;
A = 8'h8A; B = 8'h3D; #100;
A = 8'h8A; B = 8'h3E; #100;
A = 8'h8A; B = 8'h3F; #100;
A = 8'h8A; B = 8'h40; #100;
A = 8'h8A; B = 8'h41; #100;
A = 8'h8A; B = 8'h42; #100;
A = 8'h8A; B = 8'h43; #100;
A = 8'h8A; B = 8'h44; #100;
A = 8'h8A; B = 8'h45; #100;
A = 8'h8A; B = 8'h46; #100;
A = 8'h8A; B = 8'h47; #100;
A = 8'h8A; B = 8'h48; #100;
A = 8'h8A; B = 8'h49; #100;
A = 8'h8A; B = 8'h4A; #100;
A = 8'h8A; B = 8'h4B; #100;
A = 8'h8A; B = 8'h4C; #100;
A = 8'h8A; B = 8'h4D; #100;
A = 8'h8A; B = 8'h4E; #100;
A = 8'h8A; B = 8'h4F; #100;
A = 8'h8A; B = 8'h50; #100;
A = 8'h8A; B = 8'h51; #100;
A = 8'h8A; B = 8'h52; #100;
A = 8'h8A; B = 8'h53; #100;
A = 8'h8A; B = 8'h54; #100;
A = 8'h8A; B = 8'h55; #100;
A = 8'h8A; B = 8'h56; #100;
A = 8'h8A; B = 8'h57; #100;
A = 8'h8A; B = 8'h58; #100;
A = 8'h8A; B = 8'h59; #100;
A = 8'h8A; B = 8'h5A; #100;
A = 8'h8A; B = 8'h5B; #100;
A = 8'h8A; B = 8'h5C; #100;
A = 8'h8A; B = 8'h5D; #100;
A = 8'h8A; B = 8'h5E; #100;
A = 8'h8A; B = 8'h5F; #100;
A = 8'h8A; B = 8'h60; #100;
A = 8'h8A; B = 8'h61; #100;
A = 8'h8A; B = 8'h62; #100;
A = 8'h8A; B = 8'h63; #100;
A = 8'h8A; B = 8'h64; #100;
A = 8'h8A; B = 8'h65; #100;
A = 8'h8A; B = 8'h66; #100;
A = 8'h8A; B = 8'h67; #100;
A = 8'h8A; B = 8'h68; #100;
A = 8'h8A; B = 8'h69; #100;
A = 8'h8A; B = 8'h6A; #100;
A = 8'h8A; B = 8'h6B; #100;
A = 8'h8A; B = 8'h6C; #100;
A = 8'h8A; B = 8'h6D; #100;
A = 8'h8A; B = 8'h6E; #100;
A = 8'h8A; B = 8'h6F; #100;
A = 8'h8A; B = 8'h70; #100;
A = 8'h8A; B = 8'h71; #100;
A = 8'h8A; B = 8'h72; #100;
A = 8'h8A; B = 8'h73; #100;
A = 8'h8A; B = 8'h74; #100;
A = 8'h8A; B = 8'h75; #100;
A = 8'h8A; B = 8'h76; #100;
A = 8'h8A; B = 8'h77; #100;
A = 8'h8A; B = 8'h78; #100;
A = 8'h8A; B = 8'h79; #100;
A = 8'h8A; B = 8'h7A; #100;
A = 8'h8A; B = 8'h7B; #100;
A = 8'h8A; B = 8'h7C; #100;
A = 8'h8A; B = 8'h7D; #100;
A = 8'h8A; B = 8'h7E; #100;
A = 8'h8A; B = 8'h7F; #100;
A = 8'h8A; B = 8'h80; #100;
A = 8'h8A; B = 8'h81; #100;
A = 8'h8A; B = 8'h82; #100;
A = 8'h8A; B = 8'h83; #100;
A = 8'h8A; B = 8'h84; #100;
A = 8'h8A; B = 8'h85; #100;
A = 8'h8A; B = 8'h86; #100;
A = 8'h8A; B = 8'h87; #100;
A = 8'h8A; B = 8'h88; #100;
A = 8'h8A; B = 8'h89; #100;
A = 8'h8A; B = 8'h8A; #100;
A = 8'h8A; B = 8'h8B; #100;
A = 8'h8A; B = 8'h8C; #100;
A = 8'h8A; B = 8'h8D; #100;
A = 8'h8A; B = 8'h8E; #100;
A = 8'h8A; B = 8'h8F; #100;
A = 8'h8A; B = 8'h90; #100;
A = 8'h8A; B = 8'h91; #100;
A = 8'h8A; B = 8'h92; #100;
A = 8'h8A; B = 8'h93; #100;
A = 8'h8A; B = 8'h94; #100;
A = 8'h8A; B = 8'h95; #100;
A = 8'h8A; B = 8'h96; #100;
A = 8'h8A; B = 8'h97; #100;
A = 8'h8A; B = 8'h98; #100;
A = 8'h8A; B = 8'h99; #100;
A = 8'h8A; B = 8'h9A; #100;
A = 8'h8A; B = 8'h9B; #100;
A = 8'h8A; B = 8'h9C; #100;
A = 8'h8A; B = 8'h9D; #100;
A = 8'h8A; B = 8'h9E; #100;
A = 8'h8A; B = 8'h9F; #100;
A = 8'h8A; B = 8'hA0; #100;
A = 8'h8A; B = 8'hA1; #100;
A = 8'h8A; B = 8'hA2; #100;
A = 8'h8A; B = 8'hA3; #100;
A = 8'h8A; B = 8'hA4; #100;
A = 8'h8A; B = 8'hA5; #100;
A = 8'h8A; B = 8'hA6; #100;
A = 8'h8A; B = 8'hA7; #100;
A = 8'h8A; B = 8'hA8; #100;
A = 8'h8A; B = 8'hA9; #100;
A = 8'h8A; B = 8'hAA; #100;
A = 8'h8A; B = 8'hAB; #100;
A = 8'h8A; B = 8'hAC; #100;
A = 8'h8A; B = 8'hAD; #100;
A = 8'h8A; B = 8'hAE; #100;
A = 8'h8A; B = 8'hAF; #100;
A = 8'h8A; B = 8'hB0; #100;
A = 8'h8A; B = 8'hB1; #100;
A = 8'h8A; B = 8'hB2; #100;
A = 8'h8A; B = 8'hB3; #100;
A = 8'h8A; B = 8'hB4; #100;
A = 8'h8A; B = 8'hB5; #100;
A = 8'h8A; B = 8'hB6; #100;
A = 8'h8A; B = 8'hB7; #100;
A = 8'h8A; B = 8'hB8; #100;
A = 8'h8A; B = 8'hB9; #100;
A = 8'h8A; B = 8'hBA; #100;
A = 8'h8A; B = 8'hBB; #100;
A = 8'h8A; B = 8'hBC; #100;
A = 8'h8A; B = 8'hBD; #100;
A = 8'h8A; B = 8'hBE; #100;
A = 8'h8A; B = 8'hBF; #100;
A = 8'h8A; B = 8'hC0; #100;
A = 8'h8A; B = 8'hC1; #100;
A = 8'h8A; B = 8'hC2; #100;
A = 8'h8A; B = 8'hC3; #100;
A = 8'h8A; B = 8'hC4; #100;
A = 8'h8A; B = 8'hC5; #100;
A = 8'h8A; B = 8'hC6; #100;
A = 8'h8A; B = 8'hC7; #100;
A = 8'h8A; B = 8'hC8; #100;
A = 8'h8A; B = 8'hC9; #100;
A = 8'h8A; B = 8'hCA; #100;
A = 8'h8A; B = 8'hCB; #100;
A = 8'h8A; B = 8'hCC; #100;
A = 8'h8A; B = 8'hCD; #100;
A = 8'h8A; B = 8'hCE; #100;
A = 8'h8A; B = 8'hCF; #100;
A = 8'h8A; B = 8'hD0; #100;
A = 8'h8A; B = 8'hD1; #100;
A = 8'h8A; B = 8'hD2; #100;
A = 8'h8A; B = 8'hD3; #100;
A = 8'h8A; B = 8'hD4; #100;
A = 8'h8A; B = 8'hD5; #100;
A = 8'h8A; B = 8'hD6; #100;
A = 8'h8A; B = 8'hD7; #100;
A = 8'h8A; B = 8'hD8; #100;
A = 8'h8A; B = 8'hD9; #100;
A = 8'h8A; B = 8'hDA; #100;
A = 8'h8A; B = 8'hDB; #100;
A = 8'h8A; B = 8'hDC; #100;
A = 8'h8A; B = 8'hDD; #100;
A = 8'h8A; B = 8'hDE; #100;
A = 8'h8A; B = 8'hDF; #100;
A = 8'h8A; B = 8'hE0; #100;
A = 8'h8A; B = 8'hE1; #100;
A = 8'h8A; B = 8'hE2; #100;
A = 8'h8A; B = 8'hE3; #100;
A = 8'h8A; B = 8'hE4; #100;
A = 8'h8A; B = 8'hE5; #100;
A = 8'h8A; B = 8'hE6; #100;
A = 8'h8A; B = 8'hE7; #100;
A = 8'h8A; B = 8'hE8; #100;
A = 8'h8A; B = 8'hE9; #100;
A = 8'h8A; B = 8'hEA; #100;
A = 8'h8A; B = 8'hEB; #100;
A = 8'h8A; B = 8'hEC; #100;
A = 8'h8A; B = 8'hED; #100;
A = 8'h8A; B = 8'hEE; #100;
A = 8'h8A; B = 8'hEF; #100;
A = 8'h8A; B = 8'hF0; #100;
A = 8'h8A; B = 8'hF1; #100;
A = 8'h8A; B = 8'hF2; #100;
A = 8'h8A; B = 8'hF3; #100;
A = 8'h8A; B = 8'hF4; #100;
A = 8'h8A; B = 8'hF5; #100;
A = 8'h8A; B = 8'hF6; #100;
A = 8'h8A; B = 8'hF7; #100;
A = 8'h8A; B = 8'hF8; #100;
A = 8'h8A; B = 8'hF9; #100;
A = 8'h8A; B = 8'hFA; #100;
A = 8'h8A; B = 8'hFB; #100;
A = 8'h8A; B = 8'hFC; #100;
A = 8'h8A; B = 8'hFD; #100;
A = 8'h8A; B = 8'hFE; #100;
A = 8'h8A; B = 8'hFF; #100;
A = 8'h8B; B = 8'h0; #100;
A = 8'h8B; B = 8'h1; #100;
A = 8'h8B; B = 8'h2; #100;
A = 8'h8B; B = 8'h3; #100;
A = 8'h8B; B = 8'h4; #100;
A = 8'h8B; B = 8'h5; #100;
A = 8'h8B; B = 8'h6; #100;
A = 8'h8B; B = 8'h7; #100;
A = 8'h8B; B = 8'h8; #100;
A = 8'h8B; B = 8'h9; #100;
A = 8'h8B; B = 8'hA; #100;
A = 8'h8B; B = 8'hB; #100;
A = 8'h8B; B = 8'hC; #100;
A = 8'h8B; B = 8'hD; #100;
A = 8'h8B; B = 8'hE; #100;
A = 8'h8B; B = 8'hF; #100;
A = 8'h8B; B = 8'h10; #100;
A = 8'h8B; B = 8'h11; #100;
A = 8'h8B; B = 8'h12; #100;
A = 8'h8B; B = 8'h13; #100;
A = 8'h8B; B = 8'h14; #100;
A = 8'h8B; B = 8'h15; #100;
A = 8'h8B; B = 8'h16; #100;
A = 8'h8B; B = 8'h17; #100;
A = 8'h8B; B = 8'h18; #100;
A = 8'h8B; B = 8'h19; #100;
A = 8'h8B; B = 8'h1A; #100;
A = 8'h8B; B = 8'h1B; #100;
A = 8'h8B; B = 8'h1C; #100;
A = 8'h8B; B = 8'h1D; #100;
A = 8'h8B; B = 8'h1E; #100;
A = 8'h8B; B = 8'h1F; #100;
A = 8'h8B; B = 8'h20; #100;
A = 8'h8B; B = 8'h21; #100;
A = 8'h8B; B = 8'h22; #100;
A = 8'h8B; B = 8'h23; #100;
A = 8'h8B; B = 8'h24; #100;
A = 8'h8B; B = 8'h25; #100;
A = 8'h8B; B = 8'h26; #100;
A = 8'h8B; B = 8'h27; #100;
A = 8'h8B; B = 8'h28; #100;
A = 8'h8B; B = 8'h29; #100;
A = 8'h8B; B = 8'h2A; #100;
A = 8'h8B; B = 8'h2B; #100;
A = 8'h8B; B = 8'h2C; #100;
A = 8'h8B; B = 8'h2D; #100;
A = 8'h8B; B = 8'h2E; #100;
A = 8'h8B; B = 8'h2F; #100;
A = 8'h8B; B = 8'h30; #100;
A = 8'h8B; B = 8'h31; #100;
A = 8'h8B; B = 8'h32; #100;
A = 8'h8B; B = 8'h33; #100;
A = 8'h8B; B = 8'h34; #100;
A = 8'h8B; B = 8'h35; #100;
A = 8'h8B; B = 8'h36; #100;
A = 8'h8B; B = 8'h37; #100;
A = 8'h8B; B = 8'h38; #100;
A = 8'h8B; B = 8'h39; #100;
A = 8'h8B; B = 8'h3A; #100;
A = 8'h8B; B = 8'h3B; #100;
A = 8'h8B; B = 8'h3C; #100;
A = 8'h8B; B = 8'h3D; #100;
A = 8'h8B; B = 8'h3E; #100;
A = 8'h8B; B = 8'h3F; #100;
A = 8'h8B; B = 8'h40; #100;
A = 8'h8B; B = 8'h41; #100;
A = 8'h8B; B = 8'h42; #100;
A = 8'h8B; B = 8'h43; #100;
A = 8'h8B; B = 8'h44; #100;
A = 8'h8B; B = 8'h45; #100;
A = 8'h8B; B = 8'h46; #100;
A = 8'h8B; B = 8'h47; #100;
A = 8'h8B; B = 8'h48; #100;
A = 8'h8B; B = 8'h49; #100;
A = 8'h8B; B = 8'h4A; #100;
A = 8'h8B; B = 8'h4B; #100;
A = 8'h8B; B = 8'h4C; #100;
A = 8'h8B; B = 8'h4D; #100;
A = 8'h8B; B = 8'h4E; #100;
A = 8'h8B; B = 8'h4F; #100;
A = 8'h8B; B = 8'h50; #100;
A = 8'h8B; B = 8'h51; #100;
A = 8'h8B; B = 8'h52; #100;
A = 8'h8B; B = 8'h53; #100;
A = 8'h8B; B = 8'h54; #100;
A = 8'h8B; B = 8'h55; #100;
A = 8'h8B; B = 8'h56; #100;
A = 8'h8B; B = 8'h57; #100;
A = 8'h8B; B = 8'h58; #100;
A = 8'h8B; B = 8'h59; #100;
A = 8'h8B; B = 8'h5A; #100;
A = 8'h8B; B = 8'h5B; #100;
A = 8'h8B; B = 8'h5C; #100;
A = 8'h8B; B = 8'h5D; #100;
A = 8'h8B; B = 8'h5E; #100;
A = 8'h8B; B = 8'h5F; #100;
A = 8'h8B; B = 8'h60; #100;
A = 8'h8B; B = 8'h61; #100;
A = 8'h8B; B = 8'h62; #100;
A = 8'h8B; B = 8'h63; #100;
A = 8'h8B; B = 8'h64; #100;
A = 8'h8B; B = 8'h65; #100;
A = 8'h8B; B = 8'h66; #100;
A = 8'h8B; B = 8'h67; #100;
A = 8'h8B; B = 8'h68; #100;
A = 8'h8B; B = 8'h69; #100;
A = 8'h8B; B = 8'h6A; #100;
A = 8'h8B; B = 8'h6B; #100;
A = 8'h8B; B = 8'h6C; #100;
A = 8'h8B; B = 8'h6D; #100;
A = 8'h8B; B = 8'h6E; #100;
A = 8'h8B; B = 8'h6F; #100;
A = 8'h8B; B = 8'h70; #100;
A = 8'h8B; B = 8'h71; #100;
A = 8'h8B; B = 8'h72; #100;
A = 8'h8B; B = 8'h73; #100;
A = 8'h8B; B = 8'h74; #100;
A = 8'h8B; B = 8'h75; #100;
A = 8'h8B; B = 8'h76; #100;
A = 8'h8B; B = 8'h77; #100;
A = 8'h8B; B = 8'h78; #100;
A = 8'h8B; B = 8'h79; #100;
A = 8'h8B; B = 8'h7A; #100;
A = 8'h8B; B = 8'h7B; #100;
A = 8'h8B; B = 8'h7C; #100;
A = 8'h8B; B = 8'h7D; #100;
A = 8'h8B; B = 8'h7E; #100;
A = 8'h8B; B = 8'h7F; #100;
A = 8'h8B; B = 8'h80; #100;
A = 8'h8B; B = 8'h81; #100;
A = 8'h8B; B = 8'h82; #100;
A = 8'h8B; B = 8'h83; #100;
A = 8'h8B; B = 8'h84; #100;
A = 8'h8B; B = 8'h85; #100;
A = 8'h8B; B = 8'h86; #100;
A = 8'h8B; B = 8'h87; #100;
A = 8'h8B; B = 8'h88; #100;
A = 8'h8B; B = 8'h89; #100;
A = 8'h8B; B = 8'h8A; #100;
A = 8'h8B; B = 8'h8B; #100;
A = 8'h8B; B = 8'h8C; #100;
A = 8'h8B; B = 8'h8D; #100;
A = 8'h8B; B = 8'h8E; #100;
A = 8'h8B; B = 8'h8F; #100;
A = 8'h8B; B = 8'h90; #100;
A = 8'h8B; B = 8'h91; #100;
A = 8'h8B; B = 8'h92; #100;
A = 8'h8B; B = 8'h93; #100;
A = 8'h8B; B = 8'h94; #100;
A = 8'h8B; B = 8'h95; #100;
A = 8'h8B; B = 8'h96; #100;
A = 8'h8B; B = 8'h97; #100;
A = 8'h8B; B = 8'h98; #100;
A = 8'h8B; B = 8'h99; #100;
A = 8'h8B; B = 8'h9A; #100;
A = 8'h8B; B = 8'h9B; #100;
A = 8'h8B; B = 8'h9C; #100;
A = 8'h8B; B = 8'h9D; #100;
A = 8'h8B; B = 8'h9E; #100;
A = 8'h8B; B = 8'h9F; #100;
A = 8'h8B; B = 8'hA0; #100;
A = 8'h8B; B = 8'hA1; #100;
A = 8'h8B; B = 8'hA2; #100;
A = 8'h8B; B = 8'hA3; #100;
A = 8'h8B; B = 8'hA4; #100;
A = 8'h8B; B = 8'hA5; #100;
A = 8'h8B; B = 8'hA6; #100;
A = 8'h8B; B = 8'hA7; #100;
A = 8'h8B; B = 8'hA8; #100;
A = 8'h8B; B = 8'hA9; #100;
A = 8'h8B; B = 8'hAA; #100;
A = 8'h8B; B = 8'hAB; #100;
A = 8'h8B; B = 8'hAC; #100;
A = 8'h8B; B = 8'hAD; #100;
A = 8'h8B; B = 8'hAE; #100;
A = 8'h8B; B = 8'hAF; #100;
A = 8'h8B; B = 8'hB0; #100;
A = 8'h8B; B = 8'hB1; #100;
A = 8'h8B; B = 8'hB2; #100;
A = 8'h8B; B = 8'hB3; #100;
A = 8'h8B; B = 8'hB4; #100;
A = 8'h8B; B = 8'hB5; #100;
A = 8'h8B; B = 8'hB6; #100;
A = 8'h8B; B = 8'hB7; #100;
A = 8'h8B; B = 8'hB8; #100;
A = 8'h8B; B = 8'hB9; #100;
A = 8'h8B; B = 8'hBA; #100;
A = 8'h8B; B = 8'hBB; #100;
A = 8'h8B; B = 8'hBC; #100;
A = 8'h8B; B = 8'hBD; #100;
A = 8'h8B; B = 8'hBE; #100;
A = 8'h8B; B = 8'hBF; #100;
A = 8'h8B; B = 8'hC0; #100;
A = 8'h8B; B = 8'hC1; #100;
A = 8'h8B; B = 8'hC2; #100;
A = 8'h8B; B = 8'hC3; #100;
A = 8'h8B; B = 8'hC4; #100;
A = 8'h8B; B = 8'hC5; #100;
A = 8'h8B; B = 8'hC6; #100;
A = 8'h8B; B = 8'hC7; #100;
A = 8'h8B; B = 8'hC8; #100;
A = 8'h8B; B = 8'hC9; #100;
A = 8'h8B; B = 8'hCA; #100;
A = 8'h8B; B = 8'hCB; #100;
A = 8'h8B; B = 8'hCC; #100;
A = 8'h8B; B = 8'hCD; #100;
A = 8'h8B; B = 8'hCE; #100;
A = 8'h8B; B = 8'hCF; #100;
A = 8'h8B; B = 8'hD0; #100;
A = 8'h8B; B = 8'hD1; #100;
A = 8'h8B; B = 8'hD2; #100;
A = 8'h8B; B = 8'hD3; #100;
A = 8'h8B; B = 8'hD4; #100;
A = 8'h8B; B = 8'hD5; #100;
A = 8'h8B; B = 8'hD6; #100;
A = 8'h8B; B = 8'hD7; #100;
A = 8'h8B; B = 8'hD8; #100;
A = 8'h8B; B = 8'hD9; #100;
A = 8'h8B; B = 8'hDA; #100;
A = 8'h8B; B = 8'hDB; #100;
A = 8'h8B; B = 8'hDC; #100;
A = 8'h8B; B = 8'hDD; #100;
A = 8'h8B; B = 8'hDE; #100;
A = 8'h8B; B = 8'hDF; #100;
A = 8'h8B; B = 8'hE0; #100;
A = 8'h8B; B = 8'hE1; #100;
A = 8'h8B; B = 8'hE2; #100;
A = 8'h8B; B = 8'hE3; #100;
A = 8'h8B; B = 8'hE4; #100;
A = 8'h8B; B = 8'hE5; #100;
A = 8'h8B; B = 8'hE6; #100;
A = 8'h8B; B = 8'hE7; #100;
A = 8'h8B; B = 8'hE8; #100;
A = 8'h8B; B = 8'hE9; #100;
A = 8'h8B; B = 8'hEA; #100;
A = 8'h8B; B = 8'hEB; #100;
A = 8'h8B; B = 8'hEC; #100;
A = 8'h8B; B = 8'hED; #100;
A = 8'h8B; B = 8'hEE; #100;
A = 8'h8B; B = 8'hEF; #100;
A = 8'h8B; B = 8'hF0; #100;
A = 8'h8B; B = 8'hF1; #100;
A = 8'h8B; B = 8'hF2; #100;
A = 8'h8B; B = 8'hF3; #100;
A = 8'h8B; B = 8'hF4; #100;
A = 8'h8B; B = 8'hF5; #100;
A = 8'h8B; B = 8'hF6; #100;
A = 8'h8B; B = 8'hF7; #100;
A = 8'h8B; B = 8'hF8; #100;
A = 8'h8B; B = 8'hF9; #100;
A = 8'h8B; B = 8'hFA; #100;
A = 8'h8B; B = 8'hFB; #100;
A = 8'h8B; B = 8'hFC; #100;
A = 8'h8B; B = 8'hFD; #100;
A = 8'h8B; B = 8'hFE; #100;
A = 8'h8B; B = 8'hFF; #100;
A = 8'h8C; B = 8'h0; #100;
A = 8'h8C; B = 8'h1; #100;
A = 8'h8C; B = 8'h2; #100;
A = 8'h8C; B = 8'h3; #100;
A = 8'h8C; B = 8'h4; #100;
A = 8'h8C; B = 8'h5; #100;
A = 8'h8C; B = 8'h6; #100;
A = 8'h8C; B = 8'h7; #100;
A = 8'h8C; B = 8'h8; #100;
A = 8'h8C; B = 8'h9; #100;
A = 8'h8C; B = 8'hA; #100;
A = 8'h8C; B = 8'hB; #100;
A = 8'h8C; B = 8'hC; #100;
A = 8'h8C; B = 8'hD; #100;
A = 8'h8C; B = 8'hE; #100;
A = 8'h8C; B = 8'hF; #100;
A = 8'h8C; B = 8'h10; #100;
A = 8'h8C; B = 8'h11; #100;
A = 8'h8C; B = 8'h12; #100;
A = 8'h8C; B = 8'h13; #100;
A = 8'h8C; B = 8'h14; #100;
A = 8'h8C; B = 8'h15; #100;
A = 8'h8C; B = 8'h16; #100;
A = 8'h8C; B = 8'h17; #100;
A = 8'h8C; B = 8'h18; #100;
A = 8'h8C; B = 8'h19; #100;
A = 8'h8C; B = 8'h1A; #100;
A = 8'h8C; B = 8'h1B; #100;
A = 8'h8C; B = 8'h1C; #100;
A = 8'h8C; B = 8'h1D; #100;
A = 8'h8C; B = 8'h1E; #100;
A = 8'h8C; B = 8'h1F; #100;
A = 8'h8C; B = 8'h20; #100;
A = 8'h8C; B = 8'h21; #100;
A = 8'h8C; B = 8'h22; #100;
A = 8'h8C; B = 8'h23; #100;
A = 8'h8C; B = 8'h24; #100;
A = 8'h8C; B = 8'h25; #100;
A = 8'h8C; B = 8'h26; #100;
A = 8'h8C; B = 8'h27; #100;
A = 8'h8C; B = 8'h28; #100;
A = 8'h8C; B = 8'h29; #100;
A = 8'h8C; B = 8'h2A; #100;
A = 8'h8C; B = 8'h2B; #100;
A = 8'h8C; B = 8'h2C; #100;
A = 8'h8C; B = 8'h2D; #100;
A = 8'h8C; B = 8'h2E; #100;
A = 8'h8C; B = 8'h2F; #100;
A = 8'h8C; B = 8'h30; #100;
A = 8'h8C; B = 8'h31; #100;
A = 8'h8C; B = 8'h32; #100;
A = 8'h8C; B = 8'h33; #100;
A = 8'h8C; B = 8'h34; #100;
A = 8'h8C; B = 8'h35; #100;
A = 8'h8C; B = 8'h36; #100;
A = 8'h8C; B = 8'h37; #100;
A = 8'h8C; B = 8'h38; #100;
A = 8'h8C; B = 8'h39; #100;
A = 8'h8C; B = 8'h3A; #100;
A = 8'h8C; B = 8'h3B; #100;
A = 8'h8C; B = 8'h3C; #100;
A = 8'h8C; B = 8'h3D; #100;
A = 8'h8C; B = 8'h3E; #100;
A = 8'h8C; B = 8'h3F; #100;
A = 8'h8C; B = 8'h40; #100;
A = 8'h8C; B = 8'h41; #100;
A = 8'h8C; B = 8'h42; #100;
A = 8'h8C; B = 8'h43; #100;
A = 8'h8C; B = 8'h44; #100;
A = 8'h8C; B = 8'h45; #100;
A = 8'h8C; B = 8'h46; #100;
A = 8'h8C; B = 8'h47; #100;
A = 8'h8C; B = 8'h48; #100;
A = 8'h8C; B = 8'h49; #100;
A = 8'h8C; B = 8'h4A; #100;
A = 8'h8C; B = 8'h4B; #100;
A = 8'h8C; B = 8'h4C; #100;
A = 8'h8C; B = 8'h4D; #100;
A = 8'h8C; B = 8'h4E; #100;
A = 8'h8C; B = 8'h4F; #100;
A = 8'h8C; B = 8'h50; #100;
A = 8'h8C; B = 8'h51; #100;
A = 8'h8C; B = 8'h52; #100;
A = 8'h8C; B = 8'h53; #100;
A = 8'h8C; B = 8'h54; #100;
A = 8'h8C; B = 8'h55; #100;
A = 8'h8C; B = 8'h56; #100;
A = 8'h8C; B = 8'h57; #100;
A = 8'h8C; B = 8'h58; #100;
A = 8'h8C; B = 8'h59; #100;
A = 8'h8C; B = 8'h5A; #100;
A = 8'h8C; B = 8'h5B; #100;
A = 8'h8C; B = 8'h5C; #100;
A = 8'h8C; B = 8'h5D; #100;
A = 8'h8C; B = 8'h5E; #100;
A = 8'h8C; B = 8'h5F; #100;
A = 8'h8C; B = 8'h60; #100;
A = 8'h8C; B = 8'h61; #100;
A = 8'h8C; B = 8'h62; #100;
A = 8'h8C; B = 8'h63; #100;
A = 8'h8C; B = 8'h64; #100;
A = 8'h8C; B = 8'h65; #100;
A = 8'h8C; B = 8'h66; #100;
A = 8'h8C; B = 8'h67; #100;
A = 8'h8C; B = 8'h68; #100;
A = 8'h8C; B = 8'h69; #100;
A = 8'h8C; B = 8'h6A; #100;
A = 8'h8C; B = 8'h6B; #100;
A = 8'h8C; B = 8'h6C; #100;
A = 8'h8C; B = 8'h6D; #100;
A = 8'h8C; B = 8'h6E; #100;
A = 8'h8C; B = 8'h6F; #100;
A = 8'h8C; B = 8'h70; #100;
A = 8'h8C; B = 8'h71; #100;
A = 8'h8C; B = 8'h72; #100;
A = 8'h8C; B = 8'h73; #100;
A = 8'h8C; B = 8'h74; #100;
A = 8'h8C; B = 8'h75; #100;
A = 8'h8C; B = 8'h76; #100;
A = 8'h8C; B = 8'h77; #100;
A = 8'h8C; B = 8'h78; #100;
A = 8'h8C; B = 8'h79; #100;
A = 8'h8C; B = 8'h7A; #100;
A = 8'h8C; B = 8'h7B; #100;
A = 8'h8C; B = 8'h7C; #100;
A = 8'h8C; B = 8'h7D; #100;
A = 8'h8C; B = 8'h7E; #100;
A = 8'h8C; B = 8'h7F; #100;
A = 8'h8C; B = 8'h80; #100;
A = 8'h8C; B = 8'h81; #100;
A = 8'h8C; B = 8'h82; #100;
A = 8'h8C; B = 8'h83; #100;
A = 8'h8C; B = 8'h84; #100;
A = 8'h8C; B = 8'h85; #100;
A = 8'h8C; B = 8'h86; #100;
A = 8'h8C; B = 8'h87; #100;
A = 8'h8C; B = 8'h88; #100;
A = 8'h8C; B = 8'h89; #100;
A = 8'h8C; B = 8'h8A; #100;
A = 8'h8C; B = 8'h8B; #100;
A = 8'h8C; B = 8'h8C; #100;
A = 8'h8C; B = 8'h8D; #100;
A = 8'h8C; B = 8'h8E; #100;
A = 8'h8C; B = 8'h8F; #100;
A = 8'h8C; B = 8'h90; #100;
A = 8'h8C; B = 8'h91; #100;
A = 8'h8C; B = 8'h92; #100;
A = 8'h8C; B = 8'h93; #100;
A = 8'h8C; B = 8'h94; #100;
A = 8'h8C; B = 8'h95; #100;
A = 8'h8C; B = 8'h96; #100;
A = 8'h8C; B = 8'h97; #100;
A = 8'h8C; B = 8'h98; #100;
A = 8'h8C; B = 8'h99; #100;
A = 8'h8C; B = 8'h9A; #100;
A = 8'h8C; B = 8'h9B; #100;
A = 8'h8C; B = 8'h9C; #100;
A = 8'h8C; B = 8'h9D; #100;
A = 8'h8C; B = 8'h9E; #100;
A = 8'h8C; B = 8'h9F; #100;
A = 8'h8C; B = 8'hA0; #100;
A = 8'h8C; B = 8'hA1; #100;
A = 8'h8C; B = 8'hA2; #100;
A = 8'h8C; B = 8'hA3; #100;
A = 8'h8C; B = 8'hA4; #100;
A = 8'h8C; B = 8'hA5; #100;
A = 8'h8C; B = 8'hA6; #100;
A = 8'h8C; B = 8'hA7; #100;
A = 8'h8C; B = 8'hA8; #100;
A = 8'h8C; B = 8'hA9; #100;
A = 8'h8C; B = 8'hAA; #100;
A = 8'h8C; B = 8'hAB; #100;
A = 8'h8C; B = 8'hAC; #100;
A = 8'h8C; B = 8'hAD; #100;
A = 8'h8C; B = 8'hAE; #100;
A = 8'h8C; B = 8'hAF; #100;
A = 8'h8C; B = 8'hB0; #100;
A = 8'h8C; B = 8'hB1; #100;
A = 8'h8C; B = 8'hB2; #100;
A = 8'h8C; B = 8'hB3; #100;
A = 8'h8C; B = 8'hB4; #100;
A = 8'h8C; B = 8'hB5; #100;
A = 8'h8C; B = 8'hB6; #100;
A = 8'h8C; B = 8'hB7; #100;
A = 8'h8C; B = 8'hB8; #100;
A = 8'h8C; B = 8'hB9; #100;
A = 8'h8C; B = 8'hBA; #100;
A = 8'h8C; B = 8'hBB; #100;
A = 8'h8C; B = 8'hBC; #100;
A = 8'h8C; B = 8'hBD; #100;
A = 8'h8C; B = 8'hBE; #100;
A = 8'h8C; B = 8'hBF; #100;
A = 8'h8C; B = 8'hC0; #100;
A = 8'h8C; B = 8'hC1; #100;
A = 8'h8C; B = 8'hC2; #100;
A = 8'h8C; B = 8'hC3; #100;
A = 8'h8C; B = 8'hC4; #100;
A = 8'h8C; B = 8'hC5; #100;
A = 8'h8C; B = 8'hC6; #100;
A = 8'h8C; B = 8'hC7; #100;
A = 8'h8C; B = 8'hC8; #100;
A = 8'h8C; B = 8'hC9; #100;
A = 8'h8C; B = 8'hCA; #100;
A = 8'h8C; B = 8'hCB; #100;
A = 8'h8C; B = 8'hCC; #100;
A = 8'h8C; B = 8'hCD; #100;
A = 8'h8C; B = 8'hCE; #100;
A = 8'h8C; B = 8'hCF; #100;
A = 8'h8C; B = 8'hD0; #100;
A = 8'h8C; B = 8'hD1; #100;
A = 8'h8C; B = 8'hD2; #100;
A = 8'h8C; B = 8'hD3; #100;
A = 8'h8C; B = 8'hD4; #100;
A = 8'h8C; B = 8'hD5; #100;
A = 8'h8C; B = 8'hD6; #100;
A = 8'h8C; B = 8'hD7; #100;
A = 8'h8C; B = 8'hD8; #100;
A = 8'h8C; B = 8'hD9; #100;
A = 8'h8C; B = 8'hDA; #100;
A = 8'h8C; B = 8'hDB; #100;
A = 8'h8C; B = 8'hDC; #100;
A = 8'h8C; B = 8'hDD; #100;
A = 8'h8C; B = 8'hDE; #100;
A = 8'h8C; B = 8'hDF; #100;
A = 8'h8C; B = 8'hE0; #100;
A = 8'h8C; B = 8'hE1; #100;
A = 8'h8C; B = 8'hE2; #100;
A = 8'h8C; B = 8'hE3; #100;
A = 8'h8C; B = 8'hE4; #100;
A = 8'h8C; B = 8'hE5; #100;
A = 8'h8C; B = 8'hE6; #100;
A = 8'h8C; B = 8'hE7; #100;
A = 8'h8C; B = 8'hE8; #100;
A = 8'h8C; B = 8'hE9; #100;
A = 8'h8C; B = 8'hEA; #100;
A = 8'h8C; B = 8'hEB; #100;
A = 8'h8C; B = 8'hEC; #100;
A = 8'h8C; B = 8'hED; #100;
A = 8'h8C; B = 8'hEE; #100;
A = 8'h8C; B = 8'hEF; #100;
A = 8'h8C; B = 8'hF0; #100;
A = 8'h8C; B = 8'hF1; #100;
A = 8'h8C; B = 8'hF2; #100;
A = 8'h8C; B = 8'hF3; #100;
A = 8'h8C; B = 8'hF4; #100;
A = 8'h8C; B = 8'hF5; #100;
A = 8'h8C; B = 8'hF6; #100;
A = 8'h8C; B = 8'hF7; #100;
A = 8'h8C; B = 8'hF8; #100;
A = 8'h8C; B = 8'hF9; #100;
A = 8'h8C; B = 8'hFA; #100;
A = 8'h8C; B = 8'hFB; #100;
A = 8'h8C; B = 8'hFC; #100;
A = 8'h8C; B = 8'hFD; #100;
A = 8'h8C; B = 8'hFE; #100;
A = 8'h8C; B = 8'hFF; #100;
A = 8'h8D; B = 8'h0; #100;
A = 8'h8D; B = 8'h1; #100;
A = 8'h8D; B = 8'h2; #100;
A = 8'h8D; B = 8'h3; #100;
A = 8'h8D; B = 8'h4; #100;
A = 8'h8D; B = 8'h5; #100;
A = 8'h8D; B = 8'h6; #100;
A = 8'h8D; B = 8'h7; #100;
A = 8'h8D; B = 8'h8; #100;
A = 8'h8D; B = 8'h9; #100;
A = 8'h8D; B = 8'hA; #100;
A = 8'h8D; B = 8'hB; #100;
A = 8'h8D; B = 8'hC; #100;
A = 8'h8D; B = 8'hD; #100;
A = 8'h8D; B = 8'hE; #100;
A = 8'h8D; B = 8'hF; #100;
A = 8'h8D; B = 8'h10; #100;
A = 8'h8D; B = 8'h11; #100;
A = 8'h8D; B = 8'h12; #100;
A = 8'h8D; B = 8'h13; #100;
A = 8'h8D; B = 8'h14; #100;
A = 8'h8D; B = 8'h15; #100;
A = 8'h8D; B = 8'h16; #100;
A = 8'h8D; B = 8'h17; #100;
A = 8'h8D; B = 8'h18; #100;
A = 8'h8D; B = 8'h19; #100;
A = 8'h8D; B = 8'h1A; #100;
A = 8'h8D; B = 8'h1B; #100;
A = 8'h8D; B = 8'h1C; #100;
A = 8'h8D; B = 8'h1D; #100;
A = 8'h8D; B = 8'h1E; #100;
A = 8'h8D; B = 8'h1F; #100;
A = 8'h8D; B = 8'h20; #100;
A = 8'h8D; B = 8'h21; #100;
A = 8'h8D; B = 8'h22; #100;
A = 8'h8D; B = 8'h23; #100;
A = 8'h8D; B = 8'h24; #100;
A = 8'h8D; B = 8'h25; #100;
A = 8'h8D; B = 8'h26; #100;
A = 8'h8D; B = 8'h27; #100;
A = 8'h8D; B = 8'h28; #100;
A = 8'h8D; B = 8'h29; #100;
A = 8'h8D; B = 8'h2A; #100;
A = 8'h8D; B = 8'h2B; #100;
A = 8'h8D; B = 8'h2C; #100;
A = 8'h8D; B = 8'h2D; #100;
A = 8'h8D; B = 8'h2E; #100;
A = 8'h8D; B = 8'h2F; #100;
A = 8'h8D; B = 8'h30; #100;
A = 8'h8D; B = 8'h31; #100;
A = 8'h8D; B = 8'h32; #100;
A = 8'h8D; B = 8'h33; #100;
A = 8'h8D; B = 8'h34; #100;
A = 8'h8D; B = 8'h35; #100;
A = 8'h8D; B = 8'h36; #100;
A = 8'h8D; B = 8'h37; #100;
A = 8'h8D; B = 8'h38; #100;
A = 8'h8D; B = 8'h39; #100;
A = 8'h8D; B = 8'h3A; #100;
A = 8'h8D; B = 8'h3B; #100;
A = 8'h8D; B = 8'h3C; #100;
A = 8'h8D; B = 8'h3D; #100;
A = 8'h8D; B = 8'h3E; #100;
A = 8'h8D; B = 8'h3F; #100;
A = 8'h8D; B = 8'h40; #100;
A = 8'h8D; B = 8'h41; #100;
A = 8'h8D; B = 8'h42; #100;
A = 8'h8D; B = 8'h43; #100;
A = 8'h8D; B = 8'h44; #100;
A = 8'h8D; B = 8'h45; #100;
A = 8'h8D; B = 8'h46; #100;
A = 8'h8D; B = 8'h47; #100;
A = 8'h8D; B = 8'h48; #100;
A = 8'h8D; B = 8'h49; #100;
A = 8'h8D; B = 8'h4A; #100;
A = 8'h8D; B = 8'h4B; #100;
A = 8'h8D; B = 8'h4C; #100;
A = 8'h8D; B = 8'h4D; #100;
A = 8'h8D; B = 8'h4E; #100;
A = 8'h8D; B = 8'h4F; #100;
A = 8'h8D; B = 8'h50; #100;
A = 8'h8D; B = 8'h51; #100;
A = 8'h8D; B = 8'h52; #100;
A = 8'h8D; B = 8'h53; #100;
A = 8'h8D; B = 8'h54; #100;
A = 8'h8D; B = 8'h55; #100;
A = 8'h8D; B = 8'h56; #100;
A = 8'h8D; B = 8'h57; #100;
A = 8'h8D; B = 8'h58; #100;
A = 8'h8D; B = 8'h59; #100;
A = 8'h8D; B = 8'h5A; #100;
A = 8'h8D; B = 8'h5B; #100;
A = 8'h8D; B = 8'h5C; #100;
A = 8'h8D; B = 8'h5D; #100;
A = 8'h8D; B = 8'h5E; #100;
A = 8'h8D; B = 8'h5F; #100;
A = 8'h8D; B = 8'h60; #100;
A = 8'h8D; B = 8'h61; #100;
A = 8'h8D; B = 8'h62; #100;
A = 8'h8D; B = 8'h63; #100;
A = 8'h8D; B = 8'h64; #100;
A = 8'h8D; B = 8'h65; #100;
A = 8'h8D; B = 8'h66; #100;
A = 8'h8D; B = 8'h67; #100;
A = 8'h8D; B = 8'h68; #100;
A = 8'h8D; B = 8'h69; #100;
A = 8'h8D; B = 8'h6A; #100;
A = 8'h8D; B = 8'h6B; #100;
A = 8'h8D; B = 8'h6C; #100;
A = 8'h8D; B = 8'h6D; #100;
A = 8'h8D; B = 8'h6E; #100;
A = 8'h8D; B = 8'h6F; #100;
A = 8'h8D; B = 8'h70; #100;
A = 8'h8D; B = 8'h71; #100;
A = 8'h8D; B = 8'h72; #100;
A = 8'h8D; B = 8'h73; #100;
A = 8'h8D; B = 8'h74; #100;
A = 8'h8D; B = 8'h75; #100;
A = 8'h8D; B = 8'h76; #100;
A = 8'h8D; B = 8'h77; #100;
A = 8'h8D; B = 8'h78; #100;
A = 8'h8D; B = 8'h79; #100;
A = 8'h8D; B = 8'h7A; #100;
A = 8'h8D; B = 8'h7B; #100;
A = 8'h8D; B = 8'h7C; #100;
A = 8'h8D; B = 8'h7D; #100;
A = 8'h8D; B = 8'h7E; #100;
A = 8'h8D; B = 8'h7F; #100;
A = 8'h8D; B = 8'h80; #100;
A = 8'h8D; B = 8'h81; #100;
A = 8'h8D; B = 8'h82; #100;
A = 8'h8D; B = 8'h83; #100;
A = 8'h8D; B = 8'h84; #100;
A = 8'h8D; B = 8'h85; #100;
A = 8'h8D; B = 8'h86; #100;
A = 8'h8D; B = 8'h87; #100;
A = 8'h8D; B = 8'h88; #100;
A = 8'h8D; B = 8'h89; #100;
A = 8'h8D; B = 8'h8A; #100;
A = 8'h8D; B = 8'h8B; #100;
A = 8'h8D; B = 8'h8C; #100;
A = 8'h8D; B = 8'h8D; #100;
A = 8'h8D; B = 8'h8E; #100;
A = 8'h8D; B = 8'h8F; #100;
A = 8'h8D; B = 8'h90; #100;
A = 8'h8D; B = 8'h91; #100;
A = 8'h8D; B = 8'h92; #100;
A = 8'h8D; B = 8'h93; #100;
A = 8'h8D; B = 8'h94; #100;
A = 8'h8D; B = 8'h95; #100;
A = 8'h8D; B = 8'h96; #100;
A = 8'h8D; B = 8'h97; #100;
A = 8'h8D; B = 8'h98; #100;
A = 8'h8D; B = 8'h99; #100;
A = 8'h8D; B = 8'h9A; #100;
A = 8'h8D; B = 8'h9B; #100;
A = 8'h8D; B = 8'h9C; #100;
A = 8'h8D; B = 8'h9D; #100;
A = 8'h8D; B = 8'h9E; #100;
A = 8'h8D; B = 8'h9F; #100;
A = 8'h8D; B = 8'hA0; #100;
A = 8'h8D; B = 8'hA1; #100;
A = 8'h8D; B = 8'hA2; #100;
A = 8'h8D; B = 8'hA3; #100;
A = 8'h8D; B = 8'hA4; #100;
A = 8'h8D; B = 8'hA5; #100;
A = 8'h8D; B = 8'hA6; #100;
A = 8'h8D; B = 8'hA7; #100;
A = 8'h8D; B = 8'hA8; #100;
A = 8'h8D; B = 8'hA9; #100;
A = 8'h8D; B = 8'hAA; #100;
A = 8'h8D; B = 8'hAB; #100;
A = 8'h8D; B = 8'hAC; #100;
A = 8'h8D; B = 8'hAD; #100;
A = 8'h8D; B = 8'hAE; #100;
A = 8'h8D; B = 8'hAF; #100;
A = 8'h8D; B = 8'hB0; #100;
A = 8'h8D; B = 8'hB1; #100;
A = 8'h8D; B = 8'hB2; #100;
A = 8'h8D; B = 8'hB3; #100;
A = 8'h8D; B = 8'hB4; #100;
A = 8'h8D; B = 8'hB5; #100;
A = 8'h8D; B = 8'hB6; #100;
A = 8'h8D; B = 8'hB7; #100;
A = 8'h8D; B = 8'hB8; #100;
A = 8'h8D; B = 8'hB9; #100;
A = 8'h8D; B = 8'hBA; #100;
A = 8'h8D; B = 8'hBB; #100;
A = 8'h8D; B = 8'hBC; #100;
A = 8'h8D; B = 8'hBD; #100;
A = 8'h8D; B = 8'hBE; #100;
A = 8'h8D; B = 8'hBF; #100;
A = 8'h8D; B = 8'hC0; #100;
A = 8'h8D; B = 8'hC1; #100;
A = 8'h8D; B = 8'hC2; #100;
A = 8'h8D; B = 8'hC3; #100;
A = 8'h8D; B = 8'hC4; #100;
A = 8'h8D; B = 8'hC5; #100;
A = 8'h8D; B = 8'hC6; #100;
A = 8'h8D; B = 8'hC7; #100;
A = 8'h8D; B = 8'hC8; #100;
A = 8'h8D; B = 8'hC9; #100;
A = 8'h8D; B = 8'hCA; #100;
A = 8'h8D; B = 8'hCB; #100;
A = 8'h8D; B = 8'hCC; #100;
A = 8'h8D; B = 8'hCD; #100;
A = 8'h8D; B = 8'hCE; #100;
A = 8'h8D; B = 8'hCF; #100;
A = 8'h8D; B = 8'hD0; #100;
A = 8'h8D; B = 8'hD1; #100;
A = 8'h8D; B = 8'hD2; #100;
A = 8'h8D; B = 8'hD3; #100;
A = 8'h8D; B = 8'hD4; #100;
A = 8'h8D; B = 8'hD5; #100;
A = 8'h8D; B = 8'hD6; #100;
A = 8'h8D; B = 8'hD7; #100;
A = 8'h8D; B = 8'hD8; #100;
A = 8'h8D; B = 8'hD9; #100;
A = 8'h8D; B = 8'hDA; #100;
A = 8'h8D; B = 8'hDB; #100;
A = 8'h8D; B = 8'hDC; #100;
A = 8'h8D; B = 8'hDD; #100;
A = 8'h8D; B = 8'hDE; #100;
A = 8'h8D; B = 8'hDF; #100;
A = 8'h8D; B = 8'hE0; #100;
A = 8'h8D; B = 8'hE1; #100;
A = 8'h8D; B = 8'hE2; #100;
A = 8'h8D; B = 8'hE3; #100;
A = 8'h8D; B = 8'hE4; #100;
A = 8'h8D; B = 8'hE5; #100;
A = 8'h8D; B = 8'hE6; #100;
A = 8'h8D; B = 8'hE7; #100;
A = 8'h8D; B = 8'hE8; #100;
A = 8'h8D; B = 8'hE9; #100;
A = 8'h8D; B = 8'hEA; #100;
A = 8'h8D; B = 8'hEB; #100;
A = 8'h8D; B = 8'hEC; #100;
A = 8'h8D; B = 8'hED; #100;
A = 8'h8D; B = 8'hEE; #100;
A = 8'h8D; B = 8'hEF; #100;
A = 8'h8D; B = 8'hF0; #100;
A = 8'h8D; B = 8'hF1; #100;
A = 8'h8D; B = 8'hF2; #100;
A = 8'h8D; B = 8'hF3; #100;
A = 8'h8D; B = 8'hF4; #100;
A = 8'h8D; B = 8'hF5; #100;
A = 8'h8D; B = 8'hF6; #100;
A = 8'h8D; B = 8'hF7; #100;
A = 8'h8D; B = 8'hF8; #100;
A = 8'h8D; B = 8'hF9; #100;
A = 8'h8D; B = 8'hFA; #100;
A = 8'h8D; B = 8'hFB; #100;
A = 8'h8D; B = 8'hFC; #100;
A = 8'h8D; B = 8'hFD; #100;
A = 8'h8D; B = 8'hFE; #100;
A = 8'h8D; B = 8'hFF; #100;
A = 8'h8E; B = 8'h0; #100;
A = 8'h8E; B = 8'h1; #100;
A = 8'h8E; B = 8'h2; #100;
A = 8'h8E; B = 8'h3; #100;
A = 8'h8E; B = 8'h4; #100;
A = 8'h8E; B = 8'h5; #100;
A = 8'h8E; B = 8'h6; #100;
A = 8'h8E; B = 8'h7; #100;
A = 8'h8E; B = 8'h8; #100;
A = 8'h8E; B = 8'h9; #100;
A = 8'h8E; B = 8'hA; #100;
A = 8'h8E; B = 8'hB; #100;
A = 8'h8E; B = 8'hC; #100;
A = 8'h8E; B = 8'hD; #100;
A = 8'h8E; B = 8'hE; #100;
A = 8'h8E; B = 8'hF; #100;
A = 8'h8E; B = 8'h10; #100;
A = 8'h8E; B = 8'h11; #100;
A = 8'h8E; B = 8'h12; #100;
A = 8'h8E; B = 8'h13; #100;
A = 8'h8E; B = 8'h14; #100;
A = 8'h8E; B = 8'h15; #100;
A = 8'h8E; B = 8'h16; #100;
A = 8'h8E; B = 8'h17; #100;
A = 8'h8E; B = 8'h18; #100;
A = 8'h8E; B = 8'h19; #100;
A = 8'h8E; B = 8'h1A; #100;
A = 8'h8E; B = 8'h1B; #100;
A = 8'h8E; B = 8'h1C; #100;
A = 8'h8E; B = 8'h1D; #100;
A = 8'h8E; B = 8'h1E; #100;
A = 8'h8E; B = 8'h1F; #100;
A = 8'h8E; B = 8'h20; #100;
A = 8'h8E; B = 8'h21; #100;
A = 8'h8E; B = 8'h22; #100;
A = 8'h8E; B = 8'h23; #100;
A = 8'h8E; B = 8'h24; #100;
A = 8'h8E; B = 8'h25; #100;
A = 8'h8E; B = 8'h26; #100;
A = 8'h8E; B = 8'h27; #100;
A = 8'h8E; B = 8'h28; #100;
A = 8'h8E; B = 8'h29; #100;
A = 8'h8E; B = 8'h2A; #100;
A = 8'h8E; B = 8'h2B; #100;
A = 8'h8E; B = 8'h2C; #100;
A = 8'h8E; B = 8'h2D; #100;
A = 8'h8E; B = 8'h2E; #100;
A = 8'h8E; B = 8'h2F; #100;
A = 8'h8E; B = 8'h30; #100;
A = 8'h8E; B = 8'h31; #100;
A = 8'h8E; B = 8'h32; #100;
A = 8'h8E; B = 8'h33; #100;
A = 8'h8E; B = 8'h34; #100;
A = 8'h8E; B = 8'h35; #100;
A = 8'h8E; B = 8'h36; #100;
A = 8'h8E; B = 8'h37; #100;
A = 8'h8E; B = 8'h38; #100;
A = 8'h8E; B = 8'h39; #100;
A = 8'h8E; B = 8'h3A; #100;
A = 8'h8E; B = 8'h3B; #100;
A = 8'h8E; B = 8'h3C; #100;
A = 8'h8E; B = 8'h3D; #100;
A = 8'h8E; B = 8'h3E; #100;
A = 8'h8E; B = 8'h3F; #100;
A = 8'h8E; B = 8'h40; #100;
A = 8'h8E; B = 8'h41; #100;
A = 8'h8E; B = 8'h42; #100;
A = 8'h8E; B = 8'h43; #100;
A = 8'h8E; B = 8'h44; #100;
A = 8'h8E; B = 8'h45; #100;
A = 8'h8E; B = 8'h46; #100;
A = 8'h8E; B = 8'h47; #100;
A = 8'h8E; B = 8'h48; #100;
A = 8'h8E; B = 8'h49; #100;
A = 8'h8E; B = 8'h4A; #100;
A = 8'h8E; B = 8'h4B; #100;
A = 8'h8E; B = 8'h4C; #100;
A = 8'h8E; B = 8'h4D; #100;
A = 8'h8E; B = 8'h4E; #100;
A = 8'h8E; B = 8'h4F; #100;
A = 8'h8E; B = 8'h50; #100;
A = 8'h8E; B = 8'h51; #100;
A = 8'h8E; B = 8'h52; #100;
A = 8'h8E; B = 8'h53; #100;
A = 8'h8E; B = 8'h54; #100;
A = 8'h8E; B = 8'h55; #100;
A = 8'h8E; B = 8'h56; #100;
A = 8'h8E; B = 8'h57; #100;
A = 8'h8E; B = 8'h58; #100;
A = 8'h8E; B = 8'h59; #100;
A = 8'h8E; B = 8'h5A; #100;
A = 8'h8E; B = 8'h5B; #100;
A = 8'h8E; B = 8'h5C; #100;
A = 8'h8E; B = 8'h5D; #100;
A = 8'h8E; B = 8'h5E; #100;
A = 8'h8E; B = 8'h5F; #100;
A = 8'h8E; B = 8'h60; #100;
A = 8'h8E; B = 8'h61; #100;
A = 8'h8E; B = 8'h62; #100;
A = 8'h8E; B = 8'h63; #100;
A = 8'h8E; B = 8'h64; #100;
A = 8'h8E; B = 8'h65; #100;
A = 8'h8E; B = 8'h66; #100;
A = 8'h8E; B = 8'h67; #100;
A = 8'h8E; B = 8'h68; #100;
A = 8'h8E; B = 8'h69; #100;
A = 8'h8E; B = 8'h6A; #100;
A = 8'h8E; B = 8'h6B; #100;
A = 8'h8E; B = 8'h6C; #100;
A = 8'h8E; B = 8'h6D; #100;
A = 8'h8E; B = 8'h6E; #100;
A = 8'h8E; B = 8'h6F; #100;
A = 8'h8E; B = 8'h70; #100;
A = 8'h8E; B = 8'h71; #100;
A = 8'h8E; B = 8'h72; #100;
A = 8'h8E; B = 8'h73; #100;
A = 8'h8E; B = 8'h74; #100;
A = 8'h8E; B = 8'h75; #100;
A = 8'h8E; B = 8'h76; #100;
A = 8'h8E; B = 8'h77; #100;
A = 8'h8E; B = 8'h78; #100;
A = 8'h8E; B = 8'h79; #100;
A = 8'h8E; B = 8'h7A; #100;
A = 8'h8E; B = 8'h7B; #100;
A = 8'h8E; B = 8'h7C; #100;
A = 8'h8E; B = 8'h7D; #100;
A = 8'h8E; B = 8'h7E; #100;
A = 8'h8E; B = 8'h7F; #100;
A = 8'h8E; B = 8'h80; #100;
A = 8'h8E; B = 8'h81; #100;
A = 8'h8E; B = 8'h82; #100;
A = 8'h8E; B = 8'h83; #100;
A = 8'h8E; B = 8'h84; #100;
A = 8'h8E; B = 8'h85; #100;
A = 8'h8E; B = 8'h86; #100;
A = 8'h8E; B = 8'h87; #100;
A = 8'h8E; B = 8'h88; #100;
A = 8'h8E; B = 8'h89; #100;
A = 8'h8E; B = 8'h8A; #100;
A = 8'h8E; B = 8'h8B; #100;
A = 8'h8E; B = 8'h8C; #100;
A = 8'h8E; B = 8'h8D; #100;
A = 8'h8E; B = 8'h8E; #100;
A = 8'h8E; B = 8'h8F; #100;
A = 8'h8E; B = 8'h90; #100;
A = 8'h8E; B = 8'h91; #100;
A = 8'h8E; B = 8'h92; #100;
A = 8'h8E; B = 8'h93; #100;
A = 8'h8E; B = 8'h94; #100;
A = 8'h8E; B = 8'h95; #100;
A = 8'h8E; B = 8'h96; #100;
A = 8'h8E; B = 8'h97; #100;
A = 8'h8E; B = 8'h98; #100;
A = 8'h8E; B = 8'h99; #100;
A = 8'h8E; B = 8'h9A; #100;
A = 8'h8E; B = 8'h9B; #100;
A = 8'h8E; B = 8'h9C; #100;
A = 8'h8E; B = 8'h9D; #100;
A = 8'h8E; B = 8'h9E; #100;
A = 8'h8E; B = 8'h9F; #100;
A = 8'h8E; B = 8'hA0; #100;
A = 8'h8E; B = 8'hA1; #100;
A = 8'h8E; B = 8'hA2; #100;
A = 8'h8E; B = 8'hA3; #100;
A = 8'h8E; B = 8'hA4; #100;
A = 8'h8E; B = 8'hA5; #100;
A = 8'h8E; B = 8'hA6; #100;
A = 8'h8E; B = 8'hA7; #100;
A = 8'h8E; B = 8'hA8; #100;
A = 8'h8E; B = 8'hA9; #100;
A = 8'h8E; B = 8'hAA; #100;
A = 8'h8E; B = 8'hAB; #100;
A = 8'h8E; B = 8'hAC; #100;
A = 8'h8E; B = 8'hAD; #100;
A = 8'h8E; B = 8'hAE; #100;
A = 8'h8E; B = 8'hAF; #100;
A = 8'h8E; B = 8'hB0; #100;
A = 8'h8E; B = 8'hB1; #100;
A = 8'h8E; B = 8'hB2; #100;
A = 8'h8E; B = 8'hB3; #100;
A = 8'h8E; B = 8'hB4; #100;
A = 8'h8E; B = 8'hB5; #100;
A = 8'h8E; B = 8'hB6; #100;
A = 8'h8E; B = 8'hB7; #100;
A = 8'h8E; B = 8'hB8; #100;
A = 8'h8E; B = 8'hB9; #100;
A = 8'h8E; B = 8'hBA; #100;
A = 8'h8E; B = 8'hBB; #100;
A = 8'h8E; B = 8'hBC; #100;
A = 8'h8E; B = 8'hBD; #100;
A = 8'h8E; B = 8'hBE; #100;
A = 8'h8E; B = 8'hBF; #100;
A = 8'h8E; B = 8'hC0; #100;
A = 8'h8E; B = 8'hC1; #100;
A = 8'h8E; B = 8'hC2; #100;
A = 8'h8E; B = 8'hC3; #100;
A = 8'h8E; B = 8'hC4; #100;
A = 8'h8E; B = 8'hC5; #100;
A = 8'h8E; B = 8'hC6; #100;
A = 8'h8E; B = 8'hC7; #100;
A = 8'h8E; B = 8'hC8; #100;
A = 8'h8E; B = 8'hC9; #100;
A = 8'h8E; B = 8'hCA; #100;
A = 8'h8E; B = 8'hCB; #100;
A = 8'h8E; B = 8'hCC; #100;
A = 8'h8E; B = 8'hCD; #100;
A = 8'h8E; B = 8'hCE; #100;
A = 8'h8E; B = 8'hCF; #100;
A = 8'h8E; B = 8'hD0; #100;
A = 8'h8E; B = 8'hD1; #100;
A = 8'h8E; B = 8'hD2; #100;
A = 8'h8E; B = 8'hD3; #100;
A = 8'h8E; B = 8'hD4; #100;
A = 8'h8E; B = 8'hD5; #100;
A = 8'h8E; B = 8'hD6; #100;
A = 8'h8E; B = 8'hD7; #100;
A = 8'h8E; B = 8'hD8; #100;
A = 8'h8E; B = 8'hD9; #100;
A = 8'h8E; B = 8'hDA; #100;
A = 8'h8E; B = 8'hDB; #100;
A = 8'h8E; B = 8'hDC; #100;
A = 8'h8E; B = 8'hDD; #100;
A = 8'h8E; B = 8'hDE; #100;
A = 8'h8E; B = 8'hDF; #100;
A = 8'h8E; B = 8'hE0; #100;
A = 8'h8E; B = 8'hE1; #100;
A = 8'h8E; B = 8'hE2; #100;
A = 8'h8E; B = 8'hE3; #100;
A = 8'h8E; B = 8'hE4; #100;
A = 8'h8E; B = 8'hE5; #100;
A = 8'h8E; B = 8'hE6; #100;
A = 8'h8E; B = 8'hE7; #100;
A = 8'h8E; B = 8'hE8; #100;
A = 8'h8E; B = 8'hE9; #100;
A = 8'h8E; B = 8'hEA; #100;
A = 8'h8E; B = 8'hEB; #100;
A = 8'h8E; B = 8'hEC; #100;
A = 8'h8E; B = 8'hED; #100;
A = 8'h8E; B = 8'hEE; #100;
A = 8'h8E; B = 8'hEF; #100;
A = 8'h8E; B = 8'hF0; #100;
A = 8'h8E; B = 8'hF1; #100;
A = 8'h8E; B = 8'hF2; #100;
A = 8'h8E; B = 8'hF3; #100;
A = 8'h8E; B = 8'hF4; #100;
A = 8'h8E; B = 8'hF5; #100;
A = 8'h8E; B = 8'hF6; #100;
A = 8'h8E; B = 8'hF7; #100;
A = 8'h8E; B = 8'hF8; #100;
A = 8'h8E; B = 8'hF9; #100;
A = 8'h8E; B = 8'hFA; #100;
A = 8'h8E; B = 8'hFB; #100;
A = 8'h8E; B = 8'hFC; #100;
A = 8'h8E; B = 8'hFD; #100;
A = 8'h8E; B = 8'hFE; #100;
A = 8'h8E; B = 8'hFF; #100;
A = 8'h8F; B = 8'h0; #100;
A = 8'h8F; B = 8'h1; #100;
A = 8'h8F; B = 8'h2; #100;
A = 8'h8F; B = 8'h3; #100;
A = 8'h8F; B = 8'h4; #100;
A = 8'h8F; B = 8'h5; #100;
A = 8'h8F; B = 8'h6; #100;
A = 8'h8F; B = 8'h7; #100;
A = 8'h8F; B = 8'h8; #100;
A = 8'h8F; B = 8'h9; #100;
A = 8'h8F; B = 8'hA; #100;
A = 8'h8F; B = 8'hB; #100;
A = 8'h8F; B = 8'hC; #100;
A = 8'h8F; B = 8'hD; #100;
A = 8'h8F; B = 8'hE; #100;
A = 8'h8F; B = 8'hF; #100;
A = 8'h8F; B = 8'h10; #100;
A = 8'h8F; B = 8'h11; #100;
A = 8'h8F; B = 8'h12; #100;
A = 8'h8F; B = 8'h13; #100;
A = 8'h8F; B = 8'h14; #100;
A = 8'h8F; B = 8'h15; #100;
A = 8'h8F; B = 8'h16; #100;
A = 8'h8F; B = 8'h17; #100;
A = 8'h8F; B = 8'h18; #100;
A = 8'h8F; B = 8'h19; #100;
A = 8'h8F; B = 8'h1A; #100;
A = 8'h8F; B = 8'h1B; #100;
A = 8'h8F; B = 8'h1C; #100;
A = 8'h8F; B = 8'h1D; #100;
A = 8'h8F; B = 8'h1E; #100;
A = 8'h8F; B = 8'h1F; #100;
A = 8'h8F; B = 8'h20; #100;
A = 8'h8F; B = 8'h21; #100;
A = 8'h8F; B = 8'h22; #100;
A = 8'h8F; B = 8'h23; #100;
A = 8'h8F; B = 8'h24; #100;
A = 8'h8F; B = 8'h25; #100;
A = 8'h8F; B = 8'h26; #100;
A = 8'h8F; B = 8'h27; #100;
A = 8'h8F; B = 8'h28; #100;
A = 8'h8F; B = 8'h29; #100;
A = 8'h8F; B = 8'h2A; #100;
A = 8'h8F; B = 8'h2B; #100;
A = 8'h8F; B = 8'h2C; #100;
A = 8'h8F; B = 8'h2D; #100;
A = 8'h8F; B = 8'h2E; #100;
A = 8'h8F; B = 8'h2F; #100;
A = 8'h8F; B = 8'h30; #100;
A = 8'h8F; B = 8'h31; #100;
A = 8'h8F; B = 8'h32; #100;
A = 8'h8F; B = 8'h33; #100;
A = 8'h8F; B = 8'h34; #100;
A = 8'h8F; B = 8'h35; #100;
A = 8'h8F; B = 8'h36; #100;
A = 8'h8F; B = 8'h37; #100;
A = 8'h8F; B = 8'h38; #100;
A = 8'h8F; B = 8'h39; #100;
A = 8'h8F; B = 8'h3A; #100;
A = 8'h8F; B = 8'h3B; #100;
A = 8'h8F; B = 8'h3C; #100;
A = 8'h8F; B = 8'h3D; #100;
A = 8'h8F; B = 8'h3E; #100;
A = 8'h8F; B = 8'h3F; #100;
A = 8'h8F; B = 8'h40; #100;
A = 8'h8F; B = 8'h41; #100;
A = 8'h8F; B = 8'h42; #100;
A = 8'h8F; B = 8'h43; #100;
A = 8'h8F; B = 8'h44; #100;
A = 8'h8F; B = 8'h45; #100;
A = 8'h8F; B = 8'h46; #100;
A = 8'h8F; B = 8'h47; #100;
A = 8'h8F; B = 8'h48; #100;
A = 8'h8F; B = 8'h49; #100;
A = 8'h8F; B = 8'h4A; #100;
A = 8'h8F; B = 8'h4B; #100;
A = 8'h8F; B = 8'h4C; #100;
A = 8'h8F; B = 8'h4D; #100;
A = 8'h8F; B = 8'h4E; #100;
A = 8'h8F; B = 8'h4F; #100;
A = 8'h8F; B = 8'h50; #100;
A = 8'h8F; B = 8'h51; #100;
A = 8'h8F; B = 8'h52; #100;
A = 8'h8F; B = 8'h53; #100;
A = 8'h8F; B = 8'h54; #100;
A = 8'h8F; B = 8'h55; #100;
A = 8'h8F; B = 8'h56; #100;
A = 8'h8F; B = 8'h57; #100;
A = 8'h8F; B = 8'h58; #100;
A = 8'h8F; B = 8'h59; #100;
A = 8'h8F; B = 8'h5A; #100;
A = 8'h8F; B = 8'h5B; #100;
A = 8'h8F; B = 8'h5C; #100;
A = 8'h8F; B = 8'h5D; #100;
A = 8'h8F; B = 8'h5E; #100;
A = 8'h8F; B = 8'h5F; #100;
A = 8'h8F; B = 8'h60; #100;
A = 8'h8F; B = 8'h61; #100;
A = 8'h8F; B = 8'h62; #100;
A = 8'h8F; B = 8'h63; #100;
A = 8'h8F; B = 8'h64; #100;
A = 8'h8F; B = 8'h65; #100;
A = 8'h8F; B = 8'h66; #100;
A = 8'h8F; B = 8'h67; #100;
A = 8'h8F; B = 8'h68; #100;
A = 8'h8F; B = 8'h69; #100;
A = 8'h8F; B = 8'h6A; #100;
A = 8'h8F; B = 8'h6B; #100;
A = 8'h8F; B = 8'h6C; #100;
A = 8'h8F; B = 8'h6D; #100;
A = 8'h8F; B = 8'h6E; #100;
A = 8'h8F; B = 8'h6F; #100;
A = 8'h8F; B = 8'h70; #100;
A = 8'h8F; B = 8'h71; #100;
A = 8'h8F; B = 8'h72; #100;
A = 8'h8F; B = 8'h73; #100;
A = 8'h8F; B = 8'h74; #100;
A = 8'h8F; B = 8'h75; #100;
A = 8'h8F; B = 8'h76; #100;
A = 8'h8F; B = 8'h77; #100;
A = 8'h8F; B = 8'h78; #100;
A = 8'h8F; B = 8'h79; #100;
A = 8'h8F; B = 8'h7A; #100;
A = 8'h8F; B = 8'h7B; #100;
A = 8'h8F; B = 8'h7C; #100;
A = 8'h8F; B = 8'h7D; #100;
A = 8'h8F; B = 8'h7E; #100;
A = 8'h8F; B = 8'h7F; #100;
A = 8'h8F; B = 8'h80; #100;
A = 8'h8F; B = 8'h81; #100;
A = 8'h8F; B = 8'h82; #100;
A = 8'h8F; B = 8'h83; #100;
A = 8'h8F; B = 8'h84; #100;
A = 8'h8F; B = 8'h85; #100;
A = 8'h8F; B = 8'h86; #100;
A = 8'h8F; B = 8'h87; #100;
A = 8'h8F; B = 8'h88; #100;
A = 8'h8F; B = 8'h89; #100;
A = 8'h8F; B = 8'h8A; #100;
A = 8'h8F; B = 8'h8B; #100;
A = 8'h8F; B = 8'h8C; #100;
A = 8'h8F; B = 8'h8D; #100;
A = 8'h8F; B = 8'h8E; #100;
A = 8'h8F; B = 8'h8F; #100;
A = 8'h8F; B = 8'h90; #100;
A = 8'h8F; B = 8'h91; #100;
A = 8'h8F; B = 8'h92; #100;
A = 8'h8F; B = 8'h93; #100;
A = 8'h8F; B = 8'h94; #100;
A = 8'h8F; B = 8'h95; #100;
A = 8'h8F; B = 8'h96; #100;
A = 8'h8F; B = 8'h97; #100;
A = 8'h8F; B = 8'h98; #100;
A = 8'h8F; B = 8'h99; #100;
A = 8'h8F; B = 8'h9A; #100;
A = 8'h8F; B = 8'h9B; #100;
A = 8'h8F; B = 8'h9C; #100;
A = 8'h8F; B = 8'h9D; #100;
A = 8'h8F; B = 8'h9E; #100;
A = 8'h8F; B = 8'h9F; #100;
A = 8'h8F; B = 8'hA0; #100;
A = 8'h8F; B = 8'hA1; #100;
A = 8'h8F; B = 8'hA2; #100;
A = 8'h8F; B = 8'hA3; #100;
A = 8'h8F; B = 8'hA4; #100;
A = 8'h8F; B = 8'hA5; #100;
A = 8'h8F; B = 8'hA6; #100;
A = 8'h8F; B = 8'hA7; #100;
A = 8'h8F; B = 8'hA8; #100;
A = 8'h8F; B = 8'hA9; #100;
A = 8'h8F; B = 8'hAA; #100;
A = 8'h8F; B = 8'hAB; #100;
A = 8'h8F; B = 8'hAC; #100;
A = 8'h8F; B = 8'hAD; #100;
A = 8'h8F; B = 8'hAE; #100;
A = 8'h8F; B = 8'hAF; #100;
A = 8'h8F; B = 8'hB0; #100;
A = 8'h8F; B = 8'hB1; #100;
A = 8'h8F; B = 8'hB2; #100;
A = 8'h8F; B = 8'hB3; #100;
A = 8'h8F; B = 8'hB4; #100;
A = 8'h8F; B = 8'hB5; #100;
A = 8'h8F; B = 8'hB6; #100;
A = 8'h8F; B = 8'hB7; #100;
A = 8'h8F; B = 8'hB8; #100;
A = 8'h8F; B = 8'hB9; #100;
A = 8'h8F; B = 8'hBA; #100;
A = 8'h8F; B = 8'hBB; #100;
A = 8'h8F; B = 8'hBC; #100;
A = 8'h8F; B = 8'hBD; #100;
A = 8'h8F; B = 8'hBE; #100;
A = 8'h8F; B = 8'hBF; #100;
A = 8'h8F; B = 8'hC0; #100;
A = 8'h8F; B = 8'hC1; #100;
A = 8'h8F; B = 8'hC2; #100;
A = 8'h8F; B = 8'hC3; #100;
A = 8'h8F; B = 8'hC4; #100;
A = 8'h8F; B = 8'hC5; #100;
A = 8'h8F; B = 8'hC6; #100;
A = 8'h8F; B = 8'hC7; #100;
A = 8'h8F; B = 8'hC8; #100;
A = 8'h8F; B = 8'hC9; #100;
A = 8'h8F; B = 8'hCA; #100;
A = 8'h8F; B = 8'hCB; #100;
A = 8'h8F; B = 8'hCC; #100;
A = 8'h8F; B = 8'hCD; #100;
A = 8'h8F; B = 8'hCE; #100;
A = 8'h8F; B = 8'hCF; #100;
A = 8'h8F; B = 8'hD0; #100;
A = 8'h8F; B = 8'hD1; #100;
A = 8'h8F; B = 8'hD2; #100;
A = 8'h8F; B = 8'hD3; #100;
A = 8'h8F; B = 8'hD4; #100;
A = 8'h8F; B = 8'hD5; #100;
A = 8'h8F; B = 8'hD6; #100;
A = 8'h8F; B = 8'hD7; #100;
A = 8'h8F; B = 8'hD8; #100;
A = 8'h8F; B = 8'hD9; #100;
A = 8'h8F; B = 8'hDA; #100;
A = 8'h8F; B = 8'hDB; #100;
A = 8'h8F; B = 8'hDC; #100;
A = 8'h8F; B = 8'hDD; #100;
A = 8'h8F; B = 8'hDE; #100;
A = 8'h8F; B = 8'hDF; #100;
A = 8'h8F; B = 8'hE0; #100;
A = 8'h8F; B = 8'hE1; #100;
A = 8'h8F; B = 8'hE2; #100;
A = 8'h8F; B = 8'hE3; #100;
A = 8'h8F; B = 8'hE4; #100;
A = 8'h8F; B = 8'hE5; #100;
A = 8'h8F; B = 8'hE6; #100;
A = 8'h8F; B = 8'hE7; #100;
A = 8'h8F; B = 8'hE8; #100;
A = 8'h8F; B = 8'hE9; #100;
A = 8'h8F; B = 8'hEA; #100;
A = 8'h8F; B = 8'hEB; #100;
A = 8'h8F; B = 8'hEC; #100;
A = 8'h8F; B = 8'hED; #100;
A = 8'h8F; B = 8'hEE; #100;
A = 8'h8F; B = 8'hEF; #100;
A = 8'h8F; B = 8'hF0; #100;
A = 8'h8F; B = 8'hF1; #100;
A = 8'h8F; B = 8'hF2; #100;
A = 8'h8F; B = 8'hF3; #100;
A = 8'h8F; B = 8'hF4; #100;
A = 8'h8F; B = 8'hF5; #100;
A = 8'h8F; B = 8'hF6; #100;
A = 8'h8F; B = 8'hF7; #100;
A = 8'h8F; B = 8'hF8; #100;
A = 8'h8F; B = 8'hF9; #100;
A = 8'h8F; B = 8'hFA; #100;
A = 8'h8F; B = 8'hFB; #100;
A = 8'h8F; B = 8'hFC; #100;
A = 8'h8F; B = 8'hFD; #100;
A = 8'h8F; B = 8'hFE; #100;
A = 8'h8F; B = 8'hFF; #100;
A = 8'h90; B = 8'h0; #100;
A = 8'h90; B = 8'h1; #100;
A = 8'h90; B = 8'h2; #100;
A = 8'h90; B = 8'h3; #100;
A = 8'h90; B = 8'h4; #100;
A = 8'h90; B = 8'h5; #100;
A = 8'h90; B = 8'h6; #100;
A = 8'h90; B = 8'h7; #100;
A = 8'h90; B = 8'h8; #100;
A = 8'h90; B = 8'h9; #100;
A = 8'h90; B = 8'hA; #100;
A = 8'h90; B = 8'hB; #100;
A = 8'h90; B = 8'hC; #100;
A = 8'h90; B = 8'hD; #100;
A = 8'h90; B = 8'hE; #100;
A = 8'h90; B = 8'hF; #100;
A = 8'h90; B = 8'h10; #100;
A = 8'h90; B = 8'h11; #100;
A = 8'h90; B = 8'h12; #100;
A = 8'h90; B = 8'h13; #100;
A = 8'h90; B = 8'h14; #100;
A = 8'h90; B = 8'h15; #100;
A = 8'h90; B = 8'h16; #100;
A = 8'h90; B = 8'h17; #100;
A = 8'h90; B = 8'h18; #100;
A = 8'h90; B = 8'h19; #100;
A = 8'h90; B = 8'h1A; #100;
A = 8'h90; B = 8'h1B; #100;
A = 8'h90; B = 8'h1C; #100;
A = 8'h90; B = 8'h1D; #100;
A = 8'h90; B = 8'h1E; #100;
A = 8'h90; B = 8'h1F; #100;
A = 8'h90; B = 8'h20; #100;
A = 8'h90; B = 8'h21; #100;
A = 8'h90; B = 8'h22; #100;
A = 8'h90; B = 8'h23; #100;
A = 8'h90; B = 8'h24; #100;
A = 8'h90; B = 8'h25; #100;
A = 8'h90; B = 8'h26; #100;
A = 8'h90; B = 8'h27; #100;
A = 8'h90; B = 8'h28; #100;
A = 8'h90; B = 8'h29; #100;
A = 8'h90; B = 8'h2A; #100;
A = 8'h90; B = 8'h2B; #100;
A = 8'h90; B = 8'h2C; #100;
A = 8'h90; B = 8'h2D; #100;
A = 8'h90; B = 8'h2E; #100;
A = 8'h90; B = 8'h2F; #100;
A = 8'h90; B = 8'h30; #100;
A = 8'h90; B = 8'h31; #100;
A = 8'h90; B = 8'h32; #100;
A = 8'h90; B = 8'h33; #100;
A = 8'h90; B = 8'h34; #100;
A = 8'h90; B = 8'h35; #100;
A = 8'h90; B = 8'h36; #100;
A = 8'h90; B = 8'h37; #100;
A = 8'h90; B = 8'h38; #100;
A = 8'h90; B = 8'h39; #100;
A = 8'h90; B = 8'h3A; #100;
A = 8'h90; B = 8'h3B; #100;
A = 8'h90; B = 8'h3C; #100;
A = 8'h90; B = 8'h3D; #100;
A = 8'h90; B = 8'h3E; #100;
A = 8'h90; B = 8'h3F; #100;
A = 8'h90; B = 8'h40; #100;
A = 8'h90; B = 8'h41; #100;
A = 8'h90; B = 8'h42; #100;
A = 8'h90; B = 8'h43; #100;
A = 8'h90; B = 8'h44; #100;
A = 8'h90; B = 8'h45; #100;
A = 8'h90; B = 8'h46; #100;
A = 8'h90; B = 8'h47; #100;
A = 8'h90; B = 8'h48; #100;
A = 8'h90; B = 8'h49; #100;
A = 8'h90; B = 8'h4A; #100;
A = 8'h90; B = 8'h4B; #100;
A = 8'h90; B = 8'h4C; #100;
A = 8'h90; B = 8'h4D; #100;
A = 8'h90; B = 8'h4E; #100;
A = 8'h90; B = 8'h4F; #100;
A = 8'h90; B = 8'h50; #100;
A = 8'h90; B = 8'h51; #100;
A = 8'h90; B = 8'h52; #100;
A = 8'h90; B = 8'h53; #100;
A = 8'h90; B = 8'h54; #100;
A = 8'h90; B = 8'h55; #100;
A = 8'h90; B = 8'h56; #100;
A = 8'h90; B = 8'h57; #100;
A = 8'h90; B = 8'h58; #100;
A = 8'h90; B = 8'h59; #100;
A = 8'h90; B = 8'h5A; #100;
A = 8'h90; B = 8'h5B; #100;
A = 8'h90; B = 8'h5C; #100;
A = 8'h90; B = 8'h5D; #100;
A = 8'h90; B = 8'h5E; #100;
A = 8'h90; B = 8'h5F; #100;
A = 8'h90; B = 8'h60; #100;
A = 8'h90; B = 8'h61; #100;
A = 8'h90; B = 8'h62; #100;
A = 8'h90; B = 8'h63; #100;
A = 8'h90; B = 8'h64; #100;
A = 8'h90; B = 8'h65; #100;
A = 8'h90; B = 8'h66; #100;
A = 8'h90; B = 8'h67; #100;
A = 8'h90; B = 8'h68; #100;
A = 8'h90; B = 8'h69; #100;
A = 8'h90; B = 8'h6A; #100;
A = 8'h90; B = 8'h6B; #100;
A = 8'h90; B = 8'h6C; #100;
A = 8'h90; B = 8'h6D; #100;
A = 8'h90; B = 8'h6E; #100;
A = 8'h90; B = 8'h6F; #100;
A = 8'h90; B = 8'h70; #100;
A = 8'h90; B = 8'h71; #100;
A = 8'h90; B = 8'h72; #100;
A = 8'h90; B = 8'h73; #100;
A = 8'h90; B = 8'h74; #100;
A = 8'h90; B = 8'h75; #100;
A = 8'h90; B = 8'h76; #100;
A = 8'h90; B = 8'h77; #100;
A = 8'h90; B = 8'h78; #100;
A = 8'h90; B = 8'h79; #100;
A = 8'h90; B = 8'h7A; #100;
A = 8'h90; B = 8'h7B; #100;
A = 8'h90; B = 8'h7C; #100;
A = 8'h90; B = 8'h7D; #100;
A = 8'h90; B = 8'h7E; #100;
A = 8'h90; B = 8'h7F; #100;
A = 8'h90; B = 8'h80; #100;
A = 8'h90; B = 8'h81; #100;
A = 8'h90; B = 8'h82; #100;
A = 8'h90; B = 8'h83; #100;
A = 8'h90; B = 8'h84; #100;
A = 8'h90; B = 8'h85; #100;
A = 8'h90; B = 8'h86; #100;
A = 8'h90; B = 8'h87; #100;
A = 8'h90; B = 8'h88; #100;
A = 8'h90; B = 8'h89; #100;
A = 8'h90; B = 8'h8A; #100;
A = 8'h90; B = 8'h8B; #100;
A = 8'h90; B = 8'h8C; #100;
A = 8'h90; B = 8'h8D; #100;
A = 8'h90; B = 8'h8E; #100;
A = 8'h90; B = 8'h8F; #100;
A = 8'h90; B = 8'h90; #100;
A = 8'h90; B = 8'h91; #100;
A = 8'h90; B = 8'h92; #100;
A = 8'h90; B = 8'h93; #100;
A = 8'h90; B = 8'h94; #100;
A = 8'h90; B = 8'h95; #100;
A = 8'h90; B = 8'h96; #100;
A = 8'h90; B = 8'h97; #100;
A = 8'h90; B = 8'h98; #100;
A = 8'h90; B = 8'h99; #100;
A = 8'h90; B = 8'h9A; #100;
A = 8'h90; B = 8'h9B; #100;
A = 8'h90; B = 8'h9C; #100;
A = 8'h90; B = 8'h9D; #100;
A = 8'h90; B = 8'h9E; #100;
A = 8'h90; B = 8'h9F; #100;
A = 8'h90; B = 8'hA0; #100;
A = 8'h90; B = 8'hA1; #100;
A = 8'h90; B = 8'hA2; #100;
A = 8'h90; B = 8'hA3; #100;
A = 8'h90; B = 8'hA4; #100;
A = 8'h90; B = 8'hA5; #100;
A = 8'h90; B = 8'hA6; #100;
A = 8'h90; B = 8'hA7; #100;
A = 8'h90; B = 8'hA8; #100;
A = 8'h90; B = 8'hA9; #100;
A = 8'h90; B = 8'hAA; #100;
A = 8'h90; B = 8'hAB; #100;
A = 8'h90; B = 8'hAC; #100;
A = 8'h90; B = 8'hAD; #100;
A = 8'h90; B = 8'hAE; #100;
A = 8'h90; B = 8'hAF; #100;
A = 8'h90; B = 8'hB0; #100;
A = 8'h90; B = 8'hB1; #100;
A = 8'h90; B = 8'hB2; #100;
A = 8'h90; B = 8'hB3; #100;
A = 8'h90; B = 8'hB4; #100;
A = 8'h90; B = 8'hB5; #100;
A = 8'h90; B = 8'hB6; #100;
A = 8'h90; B = 8'hB7; #100;
A = 8'h90; B = 8'hB8; #100;
A = 8'h90; B = 8'hB9; #100;
A = 8'h90; B = 8'hBA; #100;
A = 8'h90; B = 8'hBB; #100;
A = 8'h90; B = 8'hBC; #100;
A = 8'h90; B = 8'hBD; #100;
A = 8'h90; B = 8'hBE; #100;
A = 8'h90; B = 8'hBF; #100;
A = 8'h90; B = 8'hC0; #100;
A = 8'h90; B = 8'hC1; #100;
A = 8'h90; B = 8'hC2; #100;
A = 8'h90; B = 8'hC3; #100;
A = 8'h90; B = 8'hC4; #100;
A = 8'h90; B = 8'hC5; #100;
A = 8'h90; B = 8'hC6; #100;
A = 8'h90; B = 8'hC7; #100;
A = 8'h90; B = 8'hC8; #100;
A = 8'h90; B = 8'hC9; #100;
A = 8'h90; B = 8'hCA; #100;
A = 8'h90; B = 8'hCB; #100;
A = 8'h90; B = 8'hCC; #100;
A = 8'h90; B = 8'hCD; #100;
A = 8'h90; B = 8'hCE; #100;
A = 8'h90; B = 8'hCF; #100;
A = 8'h90; B = 8'hD0; #100;
A = 8'h90; B = 8'hD1; #100;
A = 8'h90; B = 8'hD2; #100;
A = 8'h90; B = 8'hD3; #100;
A = 8'h90; B = 8'hD4; #100;
A = 8'h90; B = 8'hD5; #100;
A = 8'h90; B = 8'hD6; #100;
A = 8'h90; B = 8'hD7; #100;
A = 8'h90; B = 8'hD8; #100;
A = 8'h90; B = 8'hD9; #100;
A = 8'h90; B = 8'hDA; #100;
A = 8'h90; B = 8'hDB; #100;
A = 8'h90; B = 8'hDC; #100;
A = 8'h90; B = 8'hDD; #100;
A = 8'h90; B = 8'hDE; #100;
A = 8'h90; B = 8'hDF; #100;
A = 8'h90; B = 8'hE0; #100;
A = 8'h90; B = 8'hE1; #100;
A = 8'h90; B = 8'hE2; #100;
A = 8'h90; B = 8'hE3; #100;
A = 8'h90; B = 8'hE4; #100;
A = 8'h90; B = 8'hE5; #100;
A = 8'h90; B = 8'hE6; #100;
A = 8'h90; B = 8'hE7; #100;
A = 8'h90; B = 8'hE8; #100;
A = 8'h90; B = 8'hE9; #100;
A = 8'h90; B = 8'hEA; #100;
A = 8'h90; B = 8'hEB; #100;
A = 8'h90; B = 8'hEC; #100;
A = 8'h90; B = 8'hED; #100;
A = 8'h90; B = 8'hEE; #100;
A = 8'h90; B = 8'hEF; #100;
A = 8'h90; B = 8'hF0; #100;
A = 8'h90; B = 8'hF1; #100;
A = 8'h90; B = 8'hF2; #100;
A = 8'h90; B = 8'hF3; #100;
A = 8'h90; B = 8'hF4; #100;
A = 8'h90; B = 8'hF5; #100;
A = 8'h90; B = 8'hF6; #100;
A = 8'h90; B = 8'hF7; #100;
A = 8'h90; B = 8'hF8; #100;
A = 8'h90; B = 8'hF9; #100;
A = 8'h90; B = 8'hFA; #100;
A = 8'h90; B = 8'hFB; #100;
A = 8'h90; B = 8'hFC; #100;
A = 8'h90; B = 8'hFD; #100;
A = 8'h90; B = 8'hFE; #100;
A = 8'h90; B = 8'hFF; #100;
A = 8'h91; B = 8'h0; #100;
A = 8'h91; B = 8'h1; #100;
A = 8'h91; B = 8'h2; #100;
A = 8'h91; B = 8'h3; #100;
A = 8'h91; B = 8'h4; #100;
A = 8'h91; B = 8'h5; #100;
A = 8'h91; B = 8'h6; #100;
A = 8'h91; B = 8'h7; #100;
A = 8'h91; B = 8'h8; #100;
A = 8'h91; B = 8'h9; #100;
A = 8'h91; B = 8'hA; #100;
A = 8'h91; B = 8'hB; #100;
A = 8'h91; B = 8'hC; #100;
A = 8'h91; B = 8'hD; #100;
A = 8'h91; B = 8'hE; #100;
A = 8'h91; B = 8'hF; #100;
A = 8'h91; B = 8'h10; #100;
A = 8'h91; B = 8'h11; #100;
A = 8'h91; B = 8'h12; #100;
A = 8'h91; B = 8'h13; #100;
A = 8'h91; B = 8'h14; #100;
A = 8'h91; B = 8'h15; #100;
A = 8'h91; B = 8'h16; #100;
A = 8'h91; B = 8'h17; #100;
A = 8'h91; B = 8'h18; #100;
A = 8'h91; B = 8'h19; #100;
A = 8'h91; B = 8'h1A; #100;
A = 8'h91; B = 8'h1B; #100;
A = 8'h91; B = 8'h1C; #100;
A = 8'h91; B = 8'h1D; #100;
A = 8'h91; B = 8'h1E; #100;
A = 8'h91; B = 8'h1F; #100;
A = 8'h91; B = 8'h20; #100;
A = 8'h91; B = 8'h21; #100;
A = 8'h91; B = 8'h22; #100;
A = 8'h91; B = 8'h23; #100;
A = 8'h91; B = 8'h24; #100;
A = 8'h91; B = 8'h25; #100;
A = 8'h91; B = 8'h26; #100;
A = 8'h91; B = 8'h27; #100;
A = 8'h91; B = 8'h28; #100;
A = 8'h91; B = 8'h29; #100;
A = 8'h91; B = 8'h2A; #100;
A = 8'h91; B = 8'h2B; #100;
A = 8'h91; B = 8'h2C; #100;
A = 8'h91; B = 8'h2D; #100;
A = 8'h91; B = 8'h2E; #100;
A = 8'h91; B = 8'h2F; #100;
A = 8'h91; B = 8'h30; #100;
A = 8'h91; B = 8'h31; #100;
A = 8'h91; B = 8'h32; #100;
A = 8'h91; B = 8'h33; #100;
A = 8'h91; B = 8'h34; #100;
A = 8'h91; B = 8'h35; #100;
A = 8'h91; B = 8'h36; #100;
A = 8'h91; B = 8'h37; #100;
A = 8'h91; B = 8'h38; #100;
A = 8'h91; B = 8'h39; #100;
A = 8'h91; B = 8'h3A; #100;
A = 8'h91; B = 8'h3B; #100;
A = 8'h91; B = 8'h3C; #100;
A = 8'h91; B = 8'h3D; #100;
A = 8'h91; B = 8'h3E; #100;
A = 8'h91; B = 8'h3F; #100;
A = 8'h91; B = 8'h40; #100;
A = 8'h91; B = 8'h41; #100;
A = 8'h91; B = 8'h42; #100;
A = 8'h91; B = 8'h43; #100;
A = 8'h91; B = 8'h44; #100;
A = 8'h91; B = 8'h45; #100;
A = 8'h91; B = 8'h46; #100;
A = 8'h91; B = 8'h47; #100;
A = 8'h91; B = 8'h48; #100;
A = 8'h91; B = 8'h49; #100;
A = 8'h91; B = 8'h4A; #100;
A = 8'h91; B = 8'h4B; #100;
A = 8'h91; B = 8'h4C; #100;
A = 8'h91; B = 8'h4D; #100;
A = 8'h91; B = 8'h4E; #100;
A = 8'h91; B = 8'h4F; #100;
A = 8'h91; B = 8'h50; #100;
A = 8'h91; B = 8'h51; #100;
A = 8'h91; B = 8'h52; #100;
A = 8'h91; B = 8'h53; #100;
A = 8'h91; B = 8'h54; #100;
A = 8'h91; B = 8'h55; #100;
A = 8'h91; B = 8'h56; #100;
A = 8'h91; B = 8'h57; #100;
A = 8'h91; B = 8'h58; #100;
A = 8'h91; B = 8'h59; #100;
A = 8'h91; B = 8'h5A; #100;
A = 8'h91; B = 8'h5B; #100;
A = 8'h91; B = 8'h5C; #100;
A = 8'h91; B = 8'h5D; #100;
A = 8'h91; B = 8'h5E; #100;
A = 8'h91; B = 8'h5F; #100;
A = 8'h91; B = 8'h60; #100;
A = 8'h91; B = 8'h61; #100;
A = 8'h91; B = 8'h62; #100;
A = 8'h91; B = 8'h63; #100;
A = 8'h91; B = 8'h64; #100;
A = 8'h91; B = 8'h65; #100;
A = 8'h91; B = 8'h66; #100;
A = 8'h91; B = 8'h67; #100;
A = 8'h91; B = 8'h68; #100;
A = 8'h91; B = 8'h69; #100;
A = 8'h91; B = 8'h6A; #100;
A = 8'h91; B = 8'h6B; #100;
A = 8'h91; B = 8'h6C; #100;
A = 8'h91; B = 8'h6D; #100;
A = 8'h91; B = 8'h6E; #100;
A = 8'h91; B = 8'h6F; #100;
A = 8'h91; B = 8'h70; #100;
A = 8'h91; B = 8'h71; #100;
A = 8'h91; B = 8'h72; #100;
A = 8'h91; B = 8'h73; #100;
A = 8'h91; B = 8'h74; #100;
A = 8'h91; B = 8'h75; #100;
A = 8'h91; B = 8'h76; #100;
A = 8'h91; B = 8'h77; #100;
A = 8'h91; B = 8'h78; #100;
A = 8'h91; B = 8'h79; #100;
A = 8'h91; B = 8'h7A; #100;
A = 8'h91; B = 8'h7B; #100;
A = 8'h91; B = 8'h7C; #100;
A = 8'h91; B = 8'h7D; #100;
A = 8'h91; B = 8'h7E; #100;
A = 8'h91; B = 8'h7F; #100;
A = 8'h91; B = 8'h80; #100;
A = 8'h91; B = 8'h81; #100;
A = 8'h91; B = 8'h82; #100;
A = 8'h91; B = 8'h83; #100;
A = 8'h91; B = 8'h84; #100;
A = 8'h91; B = 8'h85; #100;
A = 8'h91; B = 8'h86; #100;
A = 8'h91; B = 8'h87; #100;
A = 8'h91; B = 8'h88; #100;
A = 8'h91; B = 8'h89; #100;
A = 8'h91; B = 8'h8A; #100;
A = 8'h91; B = 8'h8B; #100;
A = 8'h91; B = 8'h8C; #100;
A = 8'h91; B = 8'h8D; #100;
A = 8'h91; B = 8'h8E; #100;
A = 8'h91; B = 8'h8F; #100;
A = 8'h91; B = 8'h90; #100;
A = 8'h91; B = 8'h91; #100;
A = 8'h91; B = 8'h92; #100;
A = 8'h91; B = 8'h93; #100;
A = 8'h91; B = 8'h94; #100;
A = 8'h91; B = 8'h95; #100;
A = 8'h91; B = 8'h96; #100;
A = 8'h91; B = 8'h97; #100;
A = 8'h91; B = 8'h98; #100;
A = 8'h91; B = 8'h99; #100;
A = 8'h91; B = 8'h9A; #100;
A = 8'h91; B = 8'h9B; #100;
A = 8'h91; B = 8'h9C; #100;
A = 8'h91; B = 8'h9D; #100;
A = 8'h91; B = 8'h9E; #100;
A = 8'h91; B = 8'h9F; #100;
A = 8'h91; B = 8'hA0; #100;
A = 8'h91; B = 8'hA1; #100;
A = 8'h91; B = 8'hA2; #100;
A = 8'h91; B = 8'hA3; #100;
A = 8'h91; B = 8'hA4; #100;
A = 8'h91; B = 8'hA5; #100;
A = 8'h91; B = 8'hA6; #100;
A = 8'h91; B = 8'hA7; #100;
A = 8'h91; B = 8'hA8; #100;
A = 8'h91; B = 8'hA9; #100;
A = 8'h91; B = 8'hAA; #100;
A = 8'h91; B = 8'hAB; #100;
A = 8'h91; B = 8'hAC; #100;
A = 8'h91; B = 8'hAD; #100;
A = 8'h91; B = 8'hAE; #100;
A = 8'h91; B = 8'hAF; #100;
A = 8'h91; B = 8'hB0; #100;
A = 8'h91; B = 8'hB1; #100;
A = 8'h91; B = 8'hB2; #100;
A = 8'h91; B = 8'hB3; #100;
A = 8'h91; B = 8'hB4; #100;
A = 8'h91; B = 8'hB5; #100;
A = 8'h91; B = 8'hB6; #100;
A = 8'h91; B = 8'hB7; #100;
A = 8'h91; B = 8'hB8; #100;
A = 8'h91; B = 8'hB9; #100;
A = 8'h91; B = 8'hBA; #100;
A = 8'h91; B = 8'hBB; #100;
A = 8'h91; B = 8'hBC; #100;
A = 8'h91; B = 8'hBD; #100;
A = 8'h91; B = 8'hBE; #100;
A = 8'h91; B = 8'hBF; #100;
A = 8'h91; B = 8'hC0; #100;
A = 8'h91; B = 8'hC1; #100;
A = 8'h91; B = 8'hC2; #100;
A = 8'h91; B = 8'hC3; #100;
A = 8'h91; B = 8'hC4; #100;
A = 8'h91; B = 8'hC5; #100;
A = 8'h91; B = 8'hC6; #100;
A = 8'h91; B = 8'hC7; #100;
A = 8'h91; B = 8'hC8; #100;
A = 8'h91; B = 8'hC9; #100;
A = 8'h91; B = 8'hCA; #100;
A = 8'h91; B = 8'hCB; #100;
A = 8'h91; B = 8'hCC; #100;
A = 8'h91; B = 8'hCD; #100;
A = 8'h91; B = 8'hCE; #100;
A = 8'h91; B = 8'hCF; #100;
A = 8'h91; B = 8'hD0; #100;
A = 8'h91; B = 8'hD1; #100;
A = 8'h91; B = 8'hD2; #100;
A = 8'h91; B = 8'hD3; #100;
A = 8'h91; B = 8'hD4; #100;
A = 8'h91; B = 8'hD5; #100;
A = 8'h91; B = 8'hD6; #100;
A = 8'h91; B = 8'hD7; #100;
A = 8'h91; B = 8'hD8; #100;
A = 8'h91; B = 8'hD9; #100;
A = 8'h91; B = 8'hDA; #100;
A = 8'h91; B = 8'hDB; #100;
A = 8'h91; B = 8'hDC; #100;
A = 8'h91; B = 8'hDD; #100;
A = 8'h91; B = 8'hDE; #100;
A = 8'h91; B = 8'hDF; #100;
A = 8'h91; B = 8'hE0; #100;
A = 8'h91; B = 8'hE1; #100;
A = 8'h91; B = 8'hE2; #100;
A = 8'h91; B = 8'hE3; #100;
A = 8'h91; B = 8'hE4; #100;
A = 8'h91; B = 8'hE5; #100;
A = 8'h91; B = 8'hE6; #100;
A = 8'h91; B = 8'hE7; #100;
A = 8'h91; B = 8'hE8; #100;
A = 8'h91; B = 8'hE9; #100;
A = 8'h91; B = 8'hEA; #100;
A = 8'h91; B = 8'hEB; #100;
A = 8'h91; B = 8'hEC; #100;
A = 8'h91; B = 8'hED; #100;
A = 8'h91; B = 8'hEE; #100;
A = 8'h91; B = 8'hEF; #100;
A = 8'h91; B = 8'hF0; #100;
A = 8'h91; B = 8'hF1; #100;
A = 8'h91; B = 8'hF2; #100;
A = 8'h91; B = 8'hF3; #100;
A = 8'h91; B = 8'hF4; #100;
A = 8'h91; B = 8'hF5; #100;
A = 8'h91; B = 8'hF6; #100;
A = 8'h91; B = 8'hF7; #100;
A = 8'h91; B = 8'hF8; #100;
A = 8'h91; B = 8'hF9; #100;
A = 8'h91; B = 8'hFA; #100;
A = 8'h91; B = 8'hFB; #100;
A = 8'h91; B = 8'hFC; #100;
A = 8'h91; B = 8'hFD; #100;
A = 8'h91; B = 8'hFE; #100;
A = 8'h91; B = 8'hFF; #100;
A = 8'h92; B = 8'h0; #100;
A = 8'h92; B = 8'h1; #100;
A = 8'h92; B = 8'h2; #100;
A = 8'h92; B = 8'h3; #100;
A = 8'h92; B = 8'h4; #100;
A = 8'h92; B = 8'h5; #100;
A = 8'h92; B = 8'h6; #100;
A = 8'h92; B = 8'h7; #100;
A = 8'h92; B = 8'h8; #100;
A = 8'h92; B = 8'h9; #100;
A = 8'h92; B = 8'hA; #100;
A = 8'h92; B = 8'hB; #100;
A = 8'h92; B = 8'hC; #100;
A = 8'h92; B = 8'hD; #100;
A = 8'h92; B = 8'hE; #100;
A = 8'h92; B = 8'hF; #100;
A = 8'h92; B = 8'h10; #100;
A = 8'h92; B = 8'h11; #100;
A = 8'h92; B = 8'h12; #100;
A = 8'h92; B = 8'h13; #100;
A = 8'h92; B = 8'h14; #100;
A = 8'h92; B = 8'h15; #100;
A = 8'h92; B = 8'h16; #100;
A = 8'h92; B = 8'h17; #100;
A = 8'h92; B = 8'h18; #100;
A = 8'h92; B = 8'h19; #100;
A = 8'h92; B = 8'h1A; #100;
A = 8'h92; B = 8'h1B; #100;
A = 8'h92; B = 8'h1C; #100;
A = 8'h92; B = 8'h1D; #100;
A = 8'h92; B = 8'h1E; #100;
A = 8'h92; B = 8'h1F; #100;
A = 8'h92; B = 8'h20; #100;
A = 8'h92; B = 8'h21; #100;
A = 8'h92; B = 8'h22; #100;
A = 8'h92; B = 8'h23; #100;
A = 8'h92; B = 8'h24; #100;
A = 8'h92; B = 8'h25; #100;
A = 8'h92; B = 8'h26; #100;
A = 8'h92; B = 8'h27; #100;
A = 8'h92; B = 8'h28; #100;
A = 8'h92; B = 8'h29; #100;
A = 8'h92; B = 8'h2A; #100;
A = 8'h92; B = 8'h2B; #100;
A = 8'h92; B = 8'h2C; #100;
A = 8'h92; B = 8'h2D; #100;
A = 8'h92; B = 8'h2E; #100;
A = 8'h92; B = 8'h2F; #100;
A = 8'h92; B = 8'h30; #100;
A = 8'h92; B = 8'h31; #100;
A = 8'h92; B = 8'h32; #100;
A = 8'h92; B = 8'h33; #100;
A = 8'h92; B = 8'h34; #100;
A = 8'h92; B = 8'h35; #100;
A = 8'h92; B = 8'h36; #100;
A = 8'h92; B = 8'h37; #100;
A = 8'h92; B = 8'h38; #100;
A = 8'h92; B = 8'h39; #100;
A = 8'h92; B = 8'h3A; #100;
A = 8'h92; B = 8'h3B; #100;
A = 8'h92; B = 8'h3C; #100;
A = 8'h92; B = 8'h3D; #100;
A = 8'h92; B = 8'h3E; #100;
A = 8'h92; B = 8'h3F; #100;
A = 8'h92; B = 8'h40; #100;
A = 8'h92; B = 8'h41; #100;
A = 8'h92; B = 8'h42; #100;
A = 8'h92; B = 8'h43; #100;
A = 8'h92; B = 8'h44; #100;
A = 8'h92; B = 8'h45; #100;
A = 8'h92; B = 8'h46; #100;
A = 8'h92; B = 8'h47; #100;
A = 8'h92; B = 8'h48; #100;
A = 8'h92; B = 8'h49; #100;
A = 8'h92; B = 8'h4A; #100;
A = 8'h92; B = 8'h4B; #100;
A = 8'h92; B = 8'h4C; #100;
A = 8'h92; B = 8'h4D; #100;
A = 8'h92; B = 8'h4E; #100;
A = 8'h92; B = 8'h4F; #100;
A = 8'h92; B = 8'h50; #100;
A = 8'h92; B = 8'h51; #100;
A = 8'h92; B = 8'h52; #100;
A = 8'h92; B = 8'h53; #100;
A = 8'h92; B = 8'h54; #100;
A = 8'h92; B = 8'h55; #100;
A = 8'h92; B = 8'h56; #100;
A = 8'h92; B = 8'h57; #100;
A = 8'h92; B = 8'h58; #100;
A = 8'h92; B = 8'h59; #100;
A = 8'h92; B = 8'h5A; #100;
A = 8'h92; B = 8'h5B; #100;
A = 8'h92; B = 8'h5C; #100;
A = 8'h92; B = 8'h5D; #100;
A = 8'h92; B = 8'h5E; #100;
A = 8'h92; B = 8'h5F; #100;
A = 8'h92; B = 8'h60; #100;
A = 8'h92; B = 8'h61; #100;
A = 8'h92; B = 8'h62; #100;
A = 8'h92; B = 8'h63; #100;
A = 8'h92; B = 8'h64; #100;
A = 8'h92; B = 8'h65; #100;
A = 8'h92; B = 8'h66; #100;
A = 8'h92; B = 8'h67; #100;
A = 8'h92; B = 8'h68; #100;
A = 8'h92; B = 8'h69; #100;
A = 8'h92; B = 8'h6A; #100;
A = 8'h92; B = 8'h6B; #100;
A = 8'h92; B = 8'h6C; #100;
A = 8'h92; B = 8'h6D; #100;
A = 8'h92; B = 8'h6E; #100;
A = 8'h92; B = 8'h6F; #100;
A = 8'h92; B = 8'h70; #100;
A = 8'h92; B = 8'h71; #100;
A = 8'h92; B = 8'h72; #100;
A = 8'h92; B = 8'h73; #100;
A = 8'h92; B = 8'h74; #100;
A = 8'h92; B = 8'h75; #100;
A = 8'h92; B = 8'h76; #100;
A = 8'h92; B = 8'h77; #100;
A = 8'h92; B = 8'h78; #100;
A = 8'h92; B = 8'h79; #100;
A = 8'h92; B = 8'h7A; #100;
A = 8'h92; B = 8'h7B; #100;
A = 8'h92; B = 8'h7C; #100;
A = 8'h92; B = 8'h7D; #100;
A = 8'h92; B = 8'h7E; #100;
A = 8'h92; B = 8'h7F; #100;
A = 8'h92; B = 8'h80; #100;
A = 8'h92; B = 8'h81; #100;
A = 8'h92; B = 8'h82; #100;
A = 8'h92; B = 8'h83; #100;
A = 8'h92; B = 8'h84; #100;
A = 8'h92; B = 8'h85; #100;
A = 8'h92; B = 8'h86; #100;
A = 8'h92; B = 8'h87; #100;
A = 8'h92; B = 8'h88; #100;
A = 8'h92; B = 8'h89; #100;
A = 8'h92; B = 8'h8A; #100;
A = 8'h92; B = 8'h8B; #100;
A = 8'h92; B = 8'h8C; #100;
A = 8'h92; B = 8'h8D; #100;
A = 8'h92; B = 8'h8E; #100;
A = 8'h92; B = 8'h8F; #100;
A = 8'h92; B = 8'h90; #100;
A = 8'h92; B = 8'h91; #100;
A = 8'h92; B = 8'h92; #100;
A = 8'h92; B = 8'h93; #100;
A = 8'h92; B = 8'h94; #100;
A = 8'h92; B = 8'h95; #100;
A = 8'h92; B = 8'h96; #100;
A = 8'h92; B = 8'h97; #100;
A = 8'h92; B = 8'h98; #100;
A = 8'h92; B = 8'h99; #100;
A = 8'h92; B = 8'h9A; #100;
A = 8'h92; B = 8'h9B; #100;
A = 8'h92; B = 8'h9C; #100;
A = 8'h92; B = 8'h9D; #100;
A = 8'h92; B = 8'h9E; #100;
A = 8'h92; B = 8'h9F; #100;
A = 8'h92; B = 8'hA0; #100;
A = 8'h92; B = 8'hA1; #100;
A = 8'h92; B = 8'hA2; #100;
A = 8'h92; B = 8'hA3; #100;
A = 8'h92; B = 8'hA4; #100;
A = 8'h92; B = 8'hA5; #100;
A = 8'h92; B = 8'hA6; #100;
A = 8'h92; B = 8'hA7; #100;
A = 8'h92; B = 8'hA8; #100;
A = 8'h92; B = 8'hA9; #100;
A = 8'h92; B = 8'hAA; #100;
A = 8'h92; B = 8'hAB; #100;
A = 8'h92; B = 8'hAC; #100;
A = 8'h92; B = 8'hAD; #100;
A = 8'h92; B = 8'hAE; #100;
A = 8'h92; B = 8'hAF; #100;
A = 8'h92; B = 8'hB0; #100;
A = 8'h92; B = 8'hB1; #100;
A = 8'h92; B = 8'hB2; #100;
A = 8'h92; B = 8'hB3; #100;
A = 8'h92; B = 8'hB4; #100;
A = 8'h92; B = 8'hB5; #100;
A = 8'h92; B = 8'hB6; #100;
A = 8'h92; B = 8'hB7; #100;
A = 8'h92; B = 8'hB8; #100;
A = 8'h92; B = 8'hB9; #100;
A = 8'h92; B = 8'hBA; #100;
A = 8'h92; B = 8'hBB; #100;
A = 8'h92; B = 8'hBC; #100;
A = 8'h92; B = 8'hBD; #100;
A = 8'h92; B = 8'hBE; #100;
A = 8'h92; B = 8'hBF; #100;
A = 8'h92; B = 8'hC0; #100;
A = 8'h92; B = 8'hC1; #100;
A = 8'h92; B = 8'hC2; #100;
A = 8'h92; B = 8'hC3; #100;
A = 8'h92; B = 8'hC4; #100;
A = 8'h92; B = 8'hC5; #100;
A = 8'h92; B = 8'hC6; #100;
A = 8'h92; B = 8'hC7; #100;
A = 8'h92; B = 8'hC8; #100;
A = 8'h92; B = 8'hC9; #100;
A = 8'h92; B = 8'hCA; #100;
A = 8'h92; B = 8'hCB; #100;
A = 8'h92; B = 8'hCC; #100;
A = 8'h92; B = 8'hCD; #100;
A = 8'h92; B = 8'hCE; #100;
A = 8'h92; B = 8'hCF; #100;
A = 8'h92; B = 8'hD0; #100;
A = 8'h92; B = 8'hD1; #100;
A = 8'h92; B = 8'hD2; #100;
A = 8'h92; B = 8'hD3; #100;
A = 8'h92; B = 8'hD4; #100;
A = 8'h92; B = 8'hD5; #100;
A = 8'h92; B = 8'hD6; #100;
A = 8'h92; B = 8'hD7; #100;
A = 8'h92; B = 8'hD8; #100;
A = 8'h92; B = 8'hD9; #100;
A = 8'h92; B = 8'hDA; #100;
A = 8'h92; B = 8'hDB; #100;
A = 8'h92; B = 8'hDC; #100;
A = 8'h92; B = 8'hDD; #100;
A = 8'h92; B = 8'hDE; #100;
A = 8'h92; B = 8'hDF; #100;
A = 8'h92; B = 8'hE0; #100;
A = 8'h92; B = 8'hE1; #100;
A = 8'h92; B = 8'hE2; #100;
A = 8'h92; B = 8'hE3; #100;
A = 8'h92; B = 8'hE4; #100;
A = 8'h92; B = 8'hE5; #100;
A = 8'h92; B = 8'hE6; #100;
A = 8'h92; B = 8'hE7; #100;
A = 8'h92; B = 8'hE8; #100;
A = 8'h92; B = 8'hE9; #100;
A = 8'h92; B = 8'hEA; #100;
A = 8'h92; B = 8'hEB; #100;
A = 8'h92; B = 8'hEC; #100;
A = 8'h92; B = 8'hED; #100;
A = 8'h92; B = 8'hEE; #100;
A = 8'h92; B = 8'hEF; #100;
A = 8'h92; B = 8'hF0; #100;
A = 8'h92; B = 8'hF1; #100;
A = 8'h92; B = 8'hF2; #100;
A = 8'h92; B = 8'hF3; #100;
A = 8'h92; B = 8'hF4; #100;
A = 8'h92; B = 8'hF5; #100;
A = 8'h92; B = 8'hF6; #100;
A = 8'h92; B = 8'hF7; #100;
A = 8'h92; B = 8'hF8; #100;
A = 8'h92; B = 8'hF9; #100;
A = 8'h92; B = 8'hFA; #100;
A = 8'h92; B = 8'hFB; #100;
A = 8'h92; B = 8'hFC; #100;
A = 8'h92; B = 8'hFD; #100;
A = 8'h92; B = 8'hFE; #100;
A = 8'h92; B = 8'hFF; #100;
A = 8'h93; B = 8'h0; #100;
A = 8'h93; B = 8'h1; #100;
A = 8'h93; B = 8'h2; #100;
A = 8'h93; B = 8'h3; #100;
A = 8'h93; B = 8'h4; #100;
A = 8'h93; B = 8'h5; #100;
A = 8'h93; B = 8'h6; #100;
A = 8'h93; B = 8'h7; #100;
A = 8'h93; B = 8'h8; #100;
A = 8'h93; B = 8'h9; #100;
A = 8'h93; B = 8'hA; #100;
A = 8'h93; B = 8'hB; #100;
A = 8'h93; B = 8'hC; #100;
A = 8'h93; B = 8'hD; #100;
A = 8'h93; B = 8'hE; #100;
A = 8'h93; B = 8'hF; #100;
A = 8'h93; B = 8'h10; #100;
A = 8'h93; B = 8'h11; #100;
A = 8'h93; B = 8'h12; #100;
A = 8'h93; B = 8'h13; #100;
A = 8'h93; B = 8'h14; #100;
A = 8'h93; B = 8'h15; #100;
A = 8'h93; B = 8'h16; #100;
A = 8'h93; B = 8'h17; #100;
A = 8'h93; B = 8'h18; #100;
A = 8'h93; B = 8'h19; #100;
A = 8'h93; B = 8'h1A; #100;
A = 8'h93; B = 8'h1B; #100;
A = 8'h93; B = 8'h1C; #100;
A = 8'h93; B = 8'h1D; #100;
A = 8'h93; B = 8'h1E; #100;
A = 8'h93; B = 8'h1F; #100;
A = 8'h93; B = 8'h20; #100;
A = 8'h93; B = 8'h21; #100;
A = 8'h93; B = 8'h22; #100;
A = 8'h93; B = 8'h23; #100;
A = 8'h93; B = 8'h24; #100;
A = 8'h93; B = 8'h25; #100;
A = 8'h93; B = 8'h26; #100;
A = 8'h93; B = 8'h27; #100;
A = 8'h93; B = 8'h28; #100;
A = 8'h93; B = 8'h29; #100;
A = 8'h93; B = 8'h2A; #100;
A = 8'h93; B = 8'h2B; #100;
A = 8'h93; B = 8'h2C; #100;
A = 8'h93; B = 8'h2D; #100;
A = 8'h93; B = 8'h2E; #100;
A = 8'h93; B = 8'h2F; #100;
A = 8'h93; B = 8'h30; #100;
A = 8'h93; B = 8'h31; #100;
A = 8'h93; B = 8'h32; #100;
A = 8'h93; B = 8'h33; #100;
A = 8'h93; B = 8'h34; #100;
A = 8'h93; B = 8'h35; #100;
A = 8'h93; B = 8'h36; #100;
A = 8'h93; B = 8'h37; #100;
A = 8'h93; B = 8'h38; #100;
A = 8'h93; B = 8'h39; #100;
A = 8'h93; B = 8'h3A; #100;
A = 8'h93; B = 8'h3B; #100;
A = 8'h93; B = 8'h3C; #100;
A = 8'h93; B = 8'h3D; #100;
A = 8'h93; B = 8'h3E; #100;
A = 8'h93; B = 8'h3F; #100;
A = 8'h93; B = 8'h40; #100;
A = 8'h93; B = 8'h41; #100;
A = 8'h93; B = 8'h42; #100;
A = 8'h93; B = 8'h43; #100;
A = 8'h93; B = 8'h44; #100;
A = 8'h93; B = 8'h45; #100;
A = 8'h93; B = 8'h46; #100;
A = 8'h93; B = 8'h47; #100;
A = 8'h93; B = 8'h48; #100;
A = 8'h93; B = 8'h49; #100;
A = 8'h93; B = 8'h4A; #100;
A = 8'h93; B = 8'h4B; #100;
A = 8'h93; B = 8'h4C; #100;
A = 8'h93; B = 8'h4D; #100;
A = 8'h93; B = 8'h4E; #100;
A = 8'h93; B = 8'h4F; #100;
A = 8'h93; B = 8'h50; #100;
A = 8'h93; B = 8'h51; #100;
A = 8'h93; B = 8'h52; #100;
A = 8'h93; B = 8'h53; #100;
A = 8'h93; B = 8'h54; #100;
A = 8'h93; B = 8'h55; #100;
A = 8'h93; B = 8'h56; #100;
A = 8'h93; B = 8'h57; #100;
A = 8'h93; B = 8'h58; #100;
A = 8'h93; B = 8'h59; #100;
A = 8'h93; B = 8'h5A; #100;
A = 8'h93; B = 8'h5B; #100;
A = 8'h93; B = 8'h5C; #100;
A = 8'h93; B = 8'h5D; #100;
A = 8'h93; B = 8'h5E; #100;
A = 8'h93; B = 8'h5F; #100;
A = 8'h93; B = 8'h60; #100;
A = 8'h93; B = 8'h61; #100;
A = 8'h93; B = 8'h62; #100;
A = 8'h93; B = 8'h63; #100;
A = 8'h93; B = 8'h64; #100;
A = 8'h93; B = 8'h65; #100;
A = 8'h93; B = 8'h66; #100;
A = 8'h93; B = 8'h67; #100;
A = 8'h93; B = 8'h68; #100;
A = 8'h93; B = 8'h69; #100;
A = 8'h93; B = 8'h6A; #100;
A = 8'h93; B = 8'h6B; #100;
A = 8'h93; B = 8'h6C; #100;
A = 8'h93; B = 8'h6D; #100;
A = 8'h93; B = 8'h6E; #100;
A = 8'h93; B = 8'h6F; #100;
A = 8'h93; B = 8'h70; #100;
A = 8'h93; B = 8'h71; #100;
A = 8'h93; B = 8'h72; #100;
A = 8'h93; B = 8'h73; #100;
A = 8'h93; B = 8'h74; #100;
A = 8'h93; B = 8'h75; #100;
A = 8'h93; B = 8'h76; #100;
A = 8'h93; B = 8'h77; #100;
A = 8'h93; B = 8'h78; #100;
A = 8'h93; B = 8'h79; #100;
A = 8'h93; B = 8'h7A; #100;
A = 8'h93; B = 8'h7B; #100;
A = 8'h93; B = 8'h7C; #100;
A = 8'h93; B = 8'h7D; #100;
A = 8'h93; B = 8'h7E; #100;
A = 8'h93; B = 8'h7F; #100;
A = 8'h93; B = 8'h80; #100;
A = 8'h93; B = 8'h81; #100;
A = 8'h93; B = 8'h82; #100;
A = 8'h93; B = 8'h83; #100;
A = 8'h93; B = 8'h84; #100;
A = 8'h93; B = 8'h85; #100;
A = 8'h93; B = 8'h86; #100;
A = 8'h93; B = 8'h87; #100;
A = 8'h93; B = 8'h88; #100;
A = 8'h93; B = 8'h89; #100;
A = 8'h93; B = 8'h8A; #100;
A = 8'h93; B = 8'h8B; #100;
A = 8'h93; B = 8'h8C; #100;
A = 8'h93; B = 8'h8D; #100;
A = 8'h93; B = 8'h8E; #100;
A = 8'h93; B = 8'h8F; #100;
A = 8'h93; B = 8'h90; #100;
A = 8'h93; B = 8'h91; #100;
A = 8'h93; B = 8'h92; #100;
A = 8'h93; B = 8'h93; #100;
A = 8'h93; B = 8'h94; #100;
A = 8'h93; B = 8'h95; #100;
A = 8'h93; B = 8'h96; #100;
A = 8'h93; B = 8'h97; #100;
A = 8'h93; B = 8'h98; #100;
A = 8'h93; B = 8'h99; #100;
A = 8'h93; B = 8'h9A; #100;
A = 8'h93; B = 8'h9B; #100;
A = 8'h93; B = 8'h9C; #100;
A = 8'h93; B = 8'h9D; #100;
A = 8'h93; B = 8'h9E; #100;
A = 8'h93; B = 8'h9F; #100;
A = 8'h93; B = 8'hA0; #100;
A = 8'h93; B = 8'hA1; #100;
A = 8'h93; B = 8'hA2; #100;
A = 8'h93; B = 8'hA3; #100;
A = 8'h93; B = 8'hA4; #100;
A = 8'h93; B = 8'hA5; #100;
A = 8'h93; B = 8'hA6; #100;
A = 8'h93; B = 8'hA7; #100;
A = 8'h93; B = 8'hA8; #100;
A = 8'h93; B = 8'hA9; #100;
A = 8'h93; B = 8'hAA; #100;
A = 8'h93; B = 8'hAB; #100;
A = 8'h93; B = 8'hAC; #100;
A = 8'h93; B = 8'hAD; #100;
A = 8'h93; B = 8'hAE; #100;
A = 8'h93; B = 8'hAF; #100;
A = 8'h93; B = 8'hB0; #100;
A = 8'h93; B = 8'hB1; #100;
A = 8'h93; B = 8'hB2; #100;
A = 8'h93; B = 8'hB3; #100;
A = 8'h93; B = 8'hB4; #100;
A = 8'h93; B = 8'hB5; #100;
A = 8'h93; B = 8'hB6; #100;
A = 8'h93; B = 8'hB7; #100;
A = 8'h93; B = 8'hB8; #100;
A = 8'h93; B = 8'hB9; #100;
A = 8'h93; B = 8'hBA; #100;
A = 8'h93; B = 8'hBB; #100;
A = 8'h93; B = 8'hBC; #100;
A = 8'h93; B = 8'hBD; #100;
A = 8'h93; B = 8'hBE; #100;
A = 8'h93; B = 8'hBF; #100;
A = 8'h93; B = 8'hC0; #100;
A = 8'h93; B = 8'hC1; #100;
A = 8'h93; B = 8'hC2; #100;
A = 8'h93; B = 8'hC3; #100;
A = 8'h93; B = 8'hC4; #100;
A = 8'h93; B = 8'hC5; #100;
A = 8'h93; B = 8'hC6; #100;
A = 8'h93; B = 8'hC7; #100;
A = 8'h93; B = 8'hC8; #100;
A = 8'h93; B = 8'hC9; #100;
A = 8'h93; B = 8'hCA; #100;
A = 8'h93; B = 8'hCB; #100;
A = 8'h93; B = 8'hCC; #100;
A = 8'h93; B = 8'hCD; #100;
A = 8'h93; B = 8'hCE; #100;
A = 8'h93; B = 8'hCF; #100;
A = 8'h93; B = 8'hD0; #100;
A = 8'h93; B = 8'hD1; #100;
A = 8'h93; B = 8'hD2; #100;
A = 8'h93; B = 8'hD3; #100;
A = 8'h93; B = 8'hD4; #100;
A = 8'h93; B = 8'hD5; #100;
A = 8'h93; B = 8'hD6; #100;
A = 8'h93; B = 8'hD7; #100;
A = 8'h93; B = 8'hD8; #100;
A = 8'h93; B = 8'hD9; #100;
A = 8'h93; B = 8'hDA; #100;
A = 8'h93; B = 8'hDB; #100;
A = 8'h93; B = 8'hDC; #100;
A = 8'h93; B = 8'hDD; #100;
A = 8'h93; B = 8'hDE; #100;
A = 8'h93; B = 8'hDF; #100;
A = 8'h93; B = 8'hE0; #100;
A = 8'h93; B = 8'hE1; #100;
A = 8'h93; B = 8'hE2; #100;
A = 8'h93; B = 8'hE3; #100;
A = 8'h93; B = 8'hE4; #100;
A = 8'h93; B = 8'hE5; #100;
A = 8'h93; B = 8'hE6; #100;
A = 8'h93; B = 8'hE7; #100;
A = 8'h93; B = 8'hE8; #100;
A = 8'h93; B = 8'hE9; #100;
A = 8'h93; B = 8'hEA; #100;
A = 8'h93; B = 8'hEB; #100;
A = 8'h93; B = 8'hEC; #100;
A = 8'h93; B = 8'hED; #100;
A = 8'h93; B = 8'hEE; #100;
A = 8'h93; B = 8'hEF; #100;
A = 8'h93; B = 8'hF0; #100;
A = 8'h93; B = 8'hF1; #100;
A = 8'h93; B = 8'hF2; #100;
A = 8'h93; B = 8'hF3; #100;
A = 8'h93; B = 8'hF4; #100;
A = 8'h93; B = 8'hF5; #100;
A = 8'h93; B = 8'hF6; #100;
A = 8'h93; B = 8'hF7; #100;
A = 8'h93; B = 8'hF8; #100;
A = 8'h93; B = 8'hF9; #100;
A = 8'h93; B = 8'hFA; #100;
A = 8'h93; B = 8'hFB; #100;
A = 8'h93; B = 8'hFC; #100;
A = 8'h93; B = 8'hFD; #100;
A = 8'h93; B = 8'hFE; #100;
A = 8'h93; B = 8'hFF; #100;
A = 8'h94; B = 8'h0; #100;
A = 8'h94; B = 8'h1; #100;
A = 8'h94; B = 8'h2; #100;
A = 8'h94; B = 8'h3; #100;
A = 8'h94; B = 8'h4; #100;
A = 8'h94; B = 8'h5; #100;
A = 8'h94; B = 8'h6; #100;
A = 8'h94; B = 8'h7; #100;
A = 8'h94; B = 8'h8; #100;
A = 8'h94; B = 8'h9; #100;
A = 8'h94; B = 8'hA; #100;
A = 8'h94; B = 8'hB; #100;
A = 8'h94; B = 8'hC; #100;
A = 8'h94; B = 8'hD; #100;
A = 8'h94; B = 8'hE; #100;
A = 8'h94; B = 8'hF; #100;
A = 8'h94; B = 8'h10; #100;
A = 8'h94; B = 8'h11; #100;
A = 8'h94; B = 8'h12; #100;
A = 8'h94; B = 8'h13; #100;
A = 8'h94; B = 8'h14; #100;
A = 8'h94; B = 8'h15; #100;
A = 8'h94; B = 8'h16; #100;
A = 8'h94; B = 8'h17; #100;
A = 8'h94; B = 8'h18; #100;
A = 8'h94; B = 8'h19; #100;
A = 8'h94; B = 8'h1A; #100;
A = 8'h94; B = 8'h1B; #100;
A = 8'h94; B = 8'h1C; #100;
A = 8'h94; B = 8'h1D; #100;
A = 8'h94; B = 8'h1E; #100;
A = 8'h94; B = 8'h1F; #100;
A = 8'h94; B = 8'h20; #100;
A = 8'h94; B = 8'h21; #100;
A = 8'h94; B = 8'h22; #100;
A = 8'h94; B = 8'h23; #100;
A = 8'h94; B = 8'h24; #100;
A = 8'h94; B = 8'h25; #100;
A = 8'h94; B = 8'h26; #100;
A = 8'h94; B = 8'h27; #100;
A = 8'h94; B = 8'h28; #100;
A = 8'h94; B = 8'h29; #100;
A = 8'h94; B = 8'h2A; #100;
A = 8'h94; B = 8'h2B; #100;
A = 8'h94; B = 8'h2C; #100;
A = 8'h94; B = 8'h2D; #100;
A = 8'h94; B = 8'h2E; #100;
A = 8'h94; B = 8'h2F; #100;
A = 8'h94; B = 8'h30; #100;
A = 8'h94; B = 8'h31; #100;
A = 8'h94; B = 8'h32; #100;
A = 8'h94; B = 8'h33; #100;
A = 8'h94; B = 8'h34; #100;
A = 8'h94; B = 8'h35; #100;
A = 8'h94; B = 8'h36; #100;
A = 8'h94; B = 8'h37; #100;
A = 8'h94; B = 8'h38; #100;
A = 8'h94; B = 8'h39; #100;
A = 8'h94; B = 8'h3A; #100;
A = 8'h94; B = 8'h3B; #100;
A = 8'h94; B = 8'h3C; #100;
A = 8'h94; B = 8'h3D; #100;
A = 8'h94; B = 8'h3E; #100;
A = 8'h94; B = 8'h3F; #100;
A = 8'h94; B = 8'h40; #100;
A = 8'h94; B = 8'h41; #100;
A = 8'h94; B = 8'h42; #100;
A = 8'h94; B = 8'h43; #100;
A = 8'h94; B = 8'h44; #100;
A = 8'h94; B = 8'h45; #100;
A = 8'h94; B = 8'h46; #100;
A = 8'h94; B = 8'h47; #100;
A = 8'h94; B = 8'h48; #100;
A = 8'h94; B = 8'h49; #100;
A = 8'h94; B = 8'h4A; #100;
A = 8'h94; B = 8'h4B; #100;
A = 8'h94; B = 8'h4C; #100;
A = 8'h94; B = 8'h4D; #100;
A = 8'h94; B = 8'h4E; #100;
A = 8'h94; B = 8'h4F; #100;
A = 8'h94; B = 8'h50; #100;
A = 8'h94; B = 8'h51; #100;
A = 8'h94; B = 8'h52; #100;
A = 8'h94; B = 8'h53; #100;
A = 8'h94; B = 8'h54; #100;
A = 8'h94; B = 8'h55; #100;
A = 8'h94; B = 8'h56; #100;
A = 8'h94; B = 8'h57; #100;
A = 8'h94; B = 8'h58; #100;
A = 8'h94; B = 8'h59; #100;
A = 8'h94; B = 8'h5A; #100;
A = 8'h94; B = 8'h5B; #100;
A = 8'h94; B = 8'h5C; #100;
A = 8'h94; B = 8'h5D; #100;
A = 8'h94; B = 8'h5E; #100;
A = 8'h94; B = 8'h5F; #100;
A = 8'h94; B = 8'h60; #100;
A = 8'h94; B = 8'h61; #100;
A = 8'h94; B = 8'h62; #100;
A = 8'h94; B = 8'h63; #100;
A = 8'h94; B = 8'h64; #100;
A = 8'h94; B = 8'h65; #100;
A = 8'h94; B = 8'h66; #100;
A = 8'h94; B = 8'h67; #100;
A = 8'h94; B = 8'h68; #100;
A = 8'h94; B = 8'h69; #100;
A = 8'h94; B = 8'h6A; #100;
A = 8'h94; B = 8'h6B; #100;
A = 8'h94; B = 8'h6C; #100;
A = 8'h94; B = 8'h6D; #100;
A = 8'h94; B = 8'h6E; #100;
A = 8'h94; B = 8'h6F; #100;
A = 8'h94; B = 8'h70; #100;
A = 8'h94; B = 8'h71; #100;
A = 8'h94; B = 8'h72; #100;
A = 8'h94; B = 8'h73; #100;
A = 8'h94; B = 8'h74; #100;
A = 8'h94; B = 8'h75; #100;
A = 8'h94; B = 8'h76; #100;
A = 8'h94; B = 8'h77; #100;
A = 8'h94; B = 8'h78; #100;
A = 8'h94; B = 8'h79; #100;
A = 8'h94; B = 8'h7A; #100;
A = 8'h94; B = 8'h7B; #100;
A = 8'h94; B = 8'h7C; #100;
A = 8'h94; B = 8'h7D; #100;
A = 8'h94; B = 8'h7E; #100;
A = 8'h94; B = 8'h7F; #100;
A = 8'h94; B = 8'h80; #100;
A = 8'h94; B = 8'h81; #100;
A = 8'h94; B = 8'h82; #100;
A = 8'h94; B = 8'h83; #100;
A = 8'h94; B = 8'h84; #100;
A = 8'h94; B = 8'h85; #100;
A = 8'h94; B = 8'h86; #100;
A = 8'h94; B = 8'h87; #100;
A = 8'h94; B = 8'h88; #100;
A = 8'h94; B = 8'h89; #100;
A = 8'h94; B = 8'h8A; #100;
A = 8'h94; B = 8'h8B; #100;
A = 8'h94; B = 8'h8C; #100;
A = 8'h94; B = 8'h8D; #100;
A = 8'h94; B = 8'h8E; #100;
A = 8'h94; B = 8'h8F; #100;
A = 8'h94; B = 8'h90; #100;
A = 8'h94; B = 8'h91; #100;
A = 8'h94; B = 8'h92; #100;
A = 8'h94; B = 8'h93; #100;
A = 8'h94; B = 8'h94; #100;
A = 8'h94; B = 8'h95; #100;
A = 8'h94; B = 8'h96; #100;
A = 8'h94; B = 8'h97; #100;
A = 8'h94; B = 8'h98; #100;
A = 8'h94; B = 8'h99; #100;
A = 8'h94; B = 8'h9A; #100;
A = 8'h94; B = 8'h9B; #100;
A = 8'h94; B = 8'h9C; #100;
A = 8'h94; B = 8'h9D; #100;
A = 8'h94; B = 8'h9E; #100;
A = 8'h94; B = 8'h9F; #100;
A = 8'h94; B = 8'hA0; #100;
A = 8'h94; B = 8'hA1; #100;
A = 8'h94; B = 8'hA2; #100;
A = 8'h94; B = 8'hA3; #100;
A = 8'h94; B = 8'hA4; #100;
A = 8'h94; B = 8'hA5; #100;
A = 8'h94; B = 8'hA6; #100;
A = 8'h94; B = 8'hA7; #100;
A = 8'h94; B = 8'hA8; #100;
A = 8'h94; B = 8'hA9; #100;
A = 8'h94; B = 8'hAA; #100;
A = 8'h94; B = 8'hAB; #100;
A = 8'h94; B = 8'hAC; #100;
A = 8'h94; B = 8'hAD; #100;
A = 8'h94; B = 8'hAE; #100;
A = 8'h94; B = 8'hAF; #100;
A = 8'h94; B = 8'hB0; #100;
A = 8'h94; B = 8'hB1; #100;
A = 8'h94; B = 8'hB2; #100;
A = 8'h94; B = 8'hB3; #100;
A = 8'h94; B = 8'hB4; #100;
A = 8'h94; B = 8'hB5; #100;
A = 8'h94; B = 8'hB6; #100;
A = 8'h94; B = 8'hB7; #100;
A = 8'h94; B = 8'hB8; #100;
A = 8'h94; B = 8'hB9; #100;
A = 8'h94; B = 8'hBA; #100;
A = 8'h94; B = 8'hBB; #100;
A = 8'h94; B = 8'hBC; #100;
A = 8'h94; B = 8'hBD; #100;
A = 8'h94; B = 8'hBE; #100;
A = 8'h94; B = 8'hBF; #100;
A = 8'h94; B = 8'hC0; #100;
A = 8'h94; B = 8'hC1; #100;
A = 8'h94; B = 8'hC2; #100;
A = 8'h94; B = 8'hC3; #100;
A = 8'h94; B = 8'hC4; #100;
A = 8'h94; B = 8'hC5; #100;
A = 8'h94; B = 8'hC6; #100;
A = 8'h94; B = 8'hC7; #100;
A = 8'h94; B = 8'hC8; #100;
A = 8'h94; B = 8'hC9; #100;
A = 8'h94; B = 8'hCA; #100;
A = 8'h94; B = 8'hCB; #100;
A = 8'h94; B = 8'hCC; #100;
A = 8'h94; B = 8'hCD; #100;
A = 8'h94; B = 8'hCE; #100;
A = 8'h94; B = 8'hCF; #100;
A = 8'h94; B = 8'hD0; #100;
A = 8'h94; B = 8'hD1; #100;
A = 8'h94; B = 8'hD2; #100;
A = 8'h94; B = 8'hD3; #100;
A = 8'h94; B = 8'hD4; #100;
A = 8'h94; B = 8'hD5; #100;
A = 8'h94; B = 8'hD6; #100;
A = 8'h94; B = 8'hD7; #100;
A = 8'h94; B = 8'hD8; #100;
A = 8'h94; B = 8'hD9; #100;
A = 8'h94; B = 8'hDA; #100;
A = 8'h94; B = 8'hDB; #100;
A = 8'h94; B = 8'hDC; #100;
A = 8'h94; B = 8'hDD; #100;
A = 8'h94; B = 8'hDE; #100;
A = 8'h94; B = 8'hDF; #100;
A = 8'h94; B = 8'hE0; #100;
A = 8'h94; B = 8'hE1; #100;
A = 8'h94; B = 8'hE2; #100;
A = 8'h94; B = 8'hE3; #100;
A = 8'h94; B = 8'hE4; #100;
A = 8'h94; B = 8'hE5; #100;
A = 8'h94; B = 8'hE6; #100;
A = 8'h94; B = 8'hE7; #100;
A = 8'h94; B = 8'hE8; #100;
A = 8'h94; B = 8'hE9; #100;
A = 8'h94; B = 8'hEA; #100;
A = 8'h94; B = 8'hEB; #100;
A = 8'h94; B = 8'hEC; #100;
A = 8'h94; B = 8'hED; #100;
A = 8'h94; B = 8'hEE; #100;
A = 8'h94; B = 8'hEF; #100;
A = 8'h94; B = 8'hF0; #100;
A = 8'h94; B = 8'hF1; #100;
A = 8'h94; B = 8'hF2; #100;
A = 8'h94; B = 8'hF3; #100;
A = 8'h94; B = 8'hF4; #100;
A = 8'h94; B = 8'hF5; #100;
A = 8'h94; B = 8'hF6; #100;
A = 8'h94; B = 8'hF7; #100;
A = 8'h94; B = 8'hF8; #100;
A = 8'h94; B = 8'hF9; #100;
A = 8'h94; B = 8'hFA; #100;
A = 8'h94; B = 8'hFB; #100;
A = 8'h94; B = 8'hFC; #100;
A = 8'h94; B = 8'hFD; #100;
A = 8'h94; B = 8'hFE; #100;
A = 8'h94; B = 8'hFF; #100;
A = 8'h95; B = 8'h0; #100;
A = 8'h95; B = 8'h1; #100;
A = 8'h95; B = 8'h2; #100;
A = 8'h95; B = 8'h3; #100;
A = 8'h95; B = 8'h4; #100;
A = 8'h95; B = 8'h5; #100;
A = 8'h95; B = 8'h6; #100;
A = 8'h95; B = 8'h7; #100;
A = 8'h95; B = 8'h8; #100;
A = 8'h95; B = 8'h9; #100;
A = 8'h95; B = 8'hA; #100;
A = 8'h95; B = 8'hB; #100;
A = 8'h95; B = 8'hC; #100;
A = 8'h95; B = 8'hD; #100;
A = 8'h95; B = 8'hE; #100;
A = 8'h95; B = 8'hF; #100;
A = 8'h95; B = 8'h10; #100;
A = 8'h95; B = 8'h11; #100;
A = 8'h95; B = 8'h12; #100;
A = 8'h95; B = 8'h13; #100;
A = 8'h95; B = 8'h14; #100;
A = 8'h95; B = 8'h15; #100;
A = 8'h95; B = 8'h16; #100;
A = 8'h95; B = 8'h17; #100;
A = 8'h95; B = 8'h18; #100;
A = 8'h95; B = 8'h19; #100;
A = 8'h95; B = 8'h1A; #100;
A = 8'h95; B = 8'h1B; #100;
A = 8'h95; B = 8'h1C; #100;
A = 8'h95; B = 8'h1D; #100;
A = 8'h95; B = 8'h1E; #100;
A = 8'h95; B = 8'h1F; #100;
A = 8'h95; B = 8'h20; #100;
A = 8'h95; B = 8'h21; #100;
A = 8'h95; B = 8'h22; #100;
A = 8'h95; B = 8'h23; #100;
A = 8'h95; B = 8'h24; #100;
A = 8'h95; B = 8'h25; #100;
A = 8'h95; B = 8'h26; #100;
A = 8'h95; B = 8'h27; #100;
A = 8'h95; B = 8'h28; #100;
A = 8'h95; B = 8'h29; #100;
A = 8'h95; B = 8'h2A; #100;
A = 8'h95; B = 8'h2B; #100;
A = 8'h95; B = 8'h2C; #100;
A = 8'h95; B = 8'h2D; #100;
A = 8'h95; B = 8'h2E; #100;
A = 8'h95; B = 8'h2F; #100;
A = 8'h95; B = 8'h30; #100;
A = 8'h95; B = 8'h31; #100;
A = 8'h95; B = 8'h32; #100;
A = 8'h95; B = 8'h33; #100;
A = 8'h95; B = 8'h34; #100;
A = 8'h95; B = 8'h35; #100;
A = 8'h95; B = 8'h36; #100;
A = 8'h95; B = 8'h37; #100;
A = 8'h95; B = 8'h38; #100;
A = 8'h95; B = 8'h39; #100;
A = 8'h95; B = 8'h3A; #100;
A = 8'h95; B = 8'h3B; #100;
A = 8'h95; B = 8'h3C; #100;
A = 8'h95; B = 8'h3D; #100;
A = 8'h95; B = 8'h3E; #100;
A = 8'h95; B = 8'h3F; #100;
A = 8'h95; B = 8'h40; #100;
A = 8'h95; B = 8'h41; #100;
A = 8'h95; B = 8'h42; #100;
A = 8'h95; B = 8'h43; #100;
A = 8'h95; B = 8'h44; #100;
A = 8'h95; B = 8'h45; #100;
A = 8'h95; B = 8'h46; #100;
A = 8'h95; B = 8'h47; #100;
A = 8'h95; B = 8'h48; #100;
A = 8'h95; B = 8'h49; #100;
A = 8'h95; B = 8'h4A; #100;
A = 8'h95; B = 8'h4B; #100;
A = 8'h95; B = 8'h4C; #100;
A = 8'h95; B = 8'h4D; #100;
A = 8'h95; B = 8'h4E; #100;
A = 8'h95; B = 8'h4F; #100;
A = 8'h95; B = 8'h50; #100;
A = 8'h95; B = 8'h51; #100;
A = 8'h95; B = 8'h52; #100;
A = 8'h95; B = 8'h53; #100;
A = 8'h95; B = 8'h54; #100;
A = 8'h95; B = 8'h55; #100;
A = 8'h95; B = 8'h56; #100;
A = 8'h95; B = 8'h57; #100;
A = 8'h95; B = 8'h58; #100;
A = 8'h95; B = 8'h59; #100;
A = 8'h95; B = 8'h5A; #100;
A = 8'h95; B = 8'h5B; #100;
A = 8'h95; B = 8'h5C; #100;
A = 8'h95; B = 8'h5D; #100;
A = 8'h95; B = 8'h5E; #100;
A = 8'h95; B = 8'h5F; #100;
A = 8'h95; B = 8'h60; #100;
A = 8'h95; B = 8'h61; #100;
A = 8'h95; B = 8'h62; #100;
A = 8'h95; B = 8'h63; #100;
A = 8'h95; B = 8'h64; #100;
A = 8'h95; B = 8'h65; #100;
A = 8'h95; B = 8'h66; #100;
A = 8'h95; B = 8'h67; #100;
A = 8'h95; B = 8'h68; #100;
A = 8'h95; B = 8'h69; #100;
A = 8'h95; B = 8'h6A; #100;
A = 8'h95; B = 8'h6B; #100;
A = 8'h95; B = 8'h6C; #100;
A = 8'h95; B = 8'h6D; #100;
A = 8'h95; B = 8'h6E; #100;
A = 8'h95; B = 8'h6F; #100;
A = 8'h95; B = 8'h70; #100;
A = 8'h95; B = 8'h71; #100;
A = 8'h95; B = 8'h72; #100;
A = 8'h95; B = 8'h73; #100;
A = 8'h95; B = 8'h74; #100;
A = 8'h95; B = 8'h75; #100;
A = 8'h95; B = 8'h76; #100;
A = 8'h95; B = 8'h77; #100;
A = 8'h95; B = 8'h78; #100;
A = 8'h95; B = 8'h79; #100;
A = 8'h95; B = 8'h7A; #100;
A = 8'h95; B = 8'h7B; #100;
A = 8'h95; B = 8'h7C; #100;
A = 8'h95; B = 8'h7D; #100;
A = 8'h95; B = 8'h7E; #100;
A = 8'h95; B = 8'h7F; #100;
A = 8'h95; B = 8'h80; #100;
A = 8'h95; B = 8'h81; #100;
A = 8'h95; B = 8'h82; #100;
A = 8'h95; B = 8'h83; #100;
A = 8'h95; B = 8'h84; #100;
A = 8'h95; B = 8'h85; #100;
A = 8'h95; B = 8'h86; #100;
A = 8'h95; B = 8'h87; #100;
A = 8'h95; B = 8'h88; #100;
A = 8'h95; B = 8'h89; #100;
A = 8'h95; B = 8'h8A; #100;
A = 8'h95; B = 8'h8B; #100;
A = 8'h95; B = 8'h8C; #100;
A = 8'h95; B = 8'h8D; #100;
A = 8'h95; B = 8'h8E; #100;
A = 8'h95; B = 8'h8F; #100;
A = 8'h95; B = 8'h90; #100;
A = 8'h95; B = 8'h91; #100;
A = 8'h95; B = 8'h92; #100;
A = 8'h95; B = 8'h93; #100;
A = 8'h95; B = 8'h94; #100;
A = 8'h95; B = 8'h95; #100;
A = 8'h95; B = 8'h96; #100;
A = 8'h95; B = 8'h97; #100;
A = 8'h95; B = 8'h98; #100;
A = 8'h95; B = 8'h99; #100;
A = 8'h95; B = 8'h9A; #100;
A = 8'h95; B = 8'h9B; #100;
A = 8'h95; B = 8'h9C; #100;
A = 8'h95; B = 8'h9D; #100;
A = 8'h95; B = 8'h9E; #100;
A = 8'h95; B = 8'h9F; #100;
A = 8'h95; B = 8'hA0; #100;
A = 8'h95; B = 8'hA1; #100;
A = 8'h95; B = 8'hA2; #100;
A = 8'h95; B = 8'hA3; #100;
A = 8'h95; B = 8'hA4; #100;
A = 8'h95; B = 8'hA5; #100;
A = 8'h95; B = 8'hA6; #100;
A = 8'h95; B = 8'hA7; #100;
A = 8'h95; B = 8'hA8; #100;
A = 8'h95; B = 8'hA9; #100;
A = 8'h95; B = 8'hAA; #100;
A = 8'h95; B = 8'hAB; #100;
A = 8'h95; B = 8'hAC; #100;
A = 8'h95; B = 8'hAD; #100;
A = 8'h95; B = 8'hAE; #100;
A = 8'h95; B = 8'hAF; #100;
A = 8'h95; B = 8'hB0; #100;
A = 8'h95; B = 8'hB1; #100;
A = 8'h95; B = 8'hB2; #100;
A = 8'h95; B = 8'hB3; #100;
A = 8'h95; B = 8'hB4; #100;
A = 8'h95; B = 8'hB5; #100;
A = 8'h95; B = 8'hB6; #100;
A = 8'h95; B = 8'hB7; #100;
A = 8'h95; B = 8'hB8; #100;
A = 8'h95; B = 8'hB9; #100;
A = 8'h95; B = 8'hBA; #100;
A = 8'h95; B = 8'hBB; #100;
A = 8'h95; B = 8'hBC; #100;
A = 8'h95; B = 8'hBD; #100;
A = 8'h95; B = 8'hBE; #100;
A = 8'h95; B = 8'hBF; #100;
A = 8'h95; B = 8'hC0; #100;
A = 8'h95; B = 8'hC1; #100;
A = 8'h95; B = 8'hC2; #100;
A = 8'h95; B = 8'hC3; #100;
A = 8'h95; B = 8'hC4; #100;
A = 8'h95; B = 8'hC5; #100;
A = 8'h95; B = 8'hC6; #100;
A = 8'h95; B = 8'hC7; #100;
A = 8'h95; B = 8'hC8; #100;
A = 8'h95; B = 8'hC9; #100;
A = 8'h95; B = 8'hCA; #100;
A = 8'h95; B = 8'hCB; #100;
A = 8'h95; B = 8'hCC; #100;
A = 8'h95; B = 8'hCD; #100;
A = 8'h95; B = 8'hCE; #100;
A = 8'h95; B = 8'hCF; #100;
A = 8'h95; B = 8'hD0; #100;
A = 8'h95; B = 8'hD1; #100;
A = 8'h95; B = 8'hD2; #100;
A = 8'h95; B = 8'hD3; #100;
A = 8'h95; B = 8'hD4; #100;
A = 8'h95; B = 8'hD5; #100;
A = 8'h95; B = 8'hD6; #100;
A = 8'h95; B = 8'hD7; #100;
A = 8'h95; B = 8'hD8; #100;
A = 8'h95; B = 8'hD9; #100;
A = 8'h95; B = 8'hDA; #100;
A = 8'h95; B = 8'hDB; #100;
A = 8'h95; B = 8'hDC; #100;
A = 8'h95; B = 8'hDD; #100;
A = 8'h95; B = 8'hDE; #100;
A = 8'h95; B = 8'hDF; #100;
A = 8'h95; B = 8'hE0; #100;
A = 8'h95; B = 8'hE1; #100;
A = 8'h95; B = 8'hE2; #100;
A = 8'h95; B = 8'hE3; #100;
A = 8'h95; B = 8'hE4; #100;
A = 8'h95; B = 8'hE5; #100;
A = 8'h95; B = 8'hE6; #100;
A = 8'h95; B = 8'hE7; #100;
A = 8'h95; B = 8'hE8; #100;
A = 8'h95; B = 8'hE9; #100;
A = 8'h95; B = 8'hEA; #100;
A = 8'h95; B = 8'hEB; #100;
A = 8'h95; B = 8'hEC; #100;
A = 8'h95; B = 8'hED; #100;
A = 8'h95; B = 8'hEE; #100;
A = 8'h95; B = 8'hEF; #100;
A = 8'h95; B = 8'hF0; #100;
A = 8'h95; B = 8'hF1; #100;
A = 8'h95; B = 8'hF2; #100;
A = 8'h95; B = 8'hF3; #100;
A = 8'h95; B = 8'hF4; #100;
A = 8'h95; B = 8'hF5; #100;
A = 8'h95; B = 8'hF6; #100;
A = 8'h95; B = 8'hF7; #100;
A = 8'h95; B = 8'hF8; #100;
A = 8'h95; B = 8'hF9; #100;
A = 8'h95; B = 8'hFA; #100;
A = 8'h95; B = 8'hFB; #100;
A = 8'h95; B = 8'hFC; #100;
A = 8'h95; B = 8'hFD; #100;
A = 8'h95; B = 8'hFE; #100;
A = 8'h95; B = 8'hFF; #100;
A = 8'h96; B = 8'h0; #100;
A = 8'h96; B = 8'h1; #100;
A = 8'h96; B = 8'h2; #100;
A = 8'h96; B = 8'h3; #100;
A = 8'h96; B = 8'h4; #100;
A = 8'h96; B = 8'h5; #100;
A = 8'h96; B = 8'h6; #100;
A = 8'h96; B = 8'h7; #100;
A = 8'h96; B = 8'h8; #100;
A = 8'h96; B = 8'h9; #100;
A = 8'h96; B = 8'hA; #100;
A = 8'h96; B = 8'hB; #100;
A = 8'h96; B = 8'hC; #100;
A = 8'h96; B = 8'hD; #100;
A = 8'h96; B = 8'hE; #100;
A = 8'h96; B = 8'hF; #100;
A = 8'h96; B = 8'h10; #100;
A = 8'h96; B = 8'h11; #100;
A = 8'h96; B = 8'h12; #100;
A = 8'h96; B = 8'h13; #100;
A = 8'h96; B = 8'h14; #100;
A = 8'h96; B = 8'h15; #100;
A = 8'h96; B = 8'h16; #100;
A = 8'h96; B = 8'h17; #100;
A = 8'h96; B = 8'h18; #100;
A = 8'h96; B = 8'h19; #100;
A = 8'h96; B = 8'h1A; #100;
A = 8'h96; B = 8'h1B; #100;
A = 8'h96; B = 8'h1C; #100;
A = 8'h96; B = 8'h1D; #100;
A = 8'h96; B = 8'h1E; #100;
A = 8'h96; B = 8'h1F; #100;
A = 8'h96; B = 8'h20; #100;
A = 8'h96; B = 8'h21; #100;
A = 8'h96; B = 8'h22; #100;
A = 8'h96; B = 8'h23; #100;
A = 8'h96; B = 8'h24; #100;
A = 8'h96; B = 8'h25; #100;
A = 8'h96; B = 8'h26; #100;
A = 8'h96; B = 8'h27; #100;
A = 8'h96; B = 8'h28; #100;
A = 8'h96; B = 8'h29; #100;
A = 8'h96; B = 8'h2A; #100;
A = 8'h96; B = 8'h2B; #100;
A = 8'h96; B = 8'h2C; #100;
A = 8'h96; B = 8'h2D; #100;
A = 8'h96; B = 8'h2E; #100;
A = 8'h96; B = 8'h2F; #100;
A = 8'h96; B = 8'h30; #100;
A = 8'h96; B = 8'h31; #100;
A = 8'h96; B = 8'h32; #100;
A = 8'h96; B = 8'h33; #100;
A = 8'h96; B = 8'h34; #100;
A = 8'h96; B = 8'h35; #100;
A = 8'h96; B = 8'h36; #100;
A = 8'h96; B = 8'h37; #100;
A = 8'h96; B = 8'h38; #100;
A = 8'h96; B = 8'h39; #100;
A = 8'h96; B = 8'h3A; #100;
A = 8'h96; B = 8'h3B; #100;
A = 8'h96; B = 8'h3C; #100;
A = 8'h96; B = 8'h3D; #100;
A = 8'h96; B = 8'h3E; #100;
A = 8'h96; B = 8'h3F; #100;
A = 8'h96; B = 8'h40; #100;
A = 8'h96; B = 8'h41; #100;
A = 8'h96; B = 8'h42; #100;
A = 8'h96; B = 8'h43; #100;
A = 8'h96; B = 8'h44; #100;
A = 8'h96; B = 8'h45; #100;
A = 8'h96; B = 8'h46; #100;
A = 8'h96; B = 8'h47; #100;
A = 8'h96; B = 8'h48; #100;
A = 8'h96; B = 8'h49; #100;
A = 8'h96; B = 8'h4A; #100;
A = 8'h96; B = 8'h4B; #100;
A = 8'h96; B = 8'h4C; #100;
A = 8'h96; B = 8'h4D; #100;
A = 8'h96; B = 8'h4E; #100;
A = 8'h96; B = 8'h4F; #100;
A = 8'h96; B = 8'h50; #100;
A = 8'h96; B = 8'h51; #100;
A = 8'h96; B = 8'h52; #100;
A = 8'h96; B = 8'h53; #100;
A = 8'h96; B = 8'h54; #100;
A = 8'h96; B = 8'h55; #100;
A = 8'h96; B = 8'h56; #100;
A = 8'h96; B = 8'h57; #100;
A = 8'h96; B = 8'h58; #100;
A = 8'h96; B = 8'h59; #100;
A = 8'h96; B = 8'h5A; #100;
A = 8'h96; B = 8'h5B; #100;
A = 8'h96; B = 8'h5C; #100;
A = 8'h96; B = 8'h5D; #100;
A = 8'h96; B = 8'h5E; #100;
A = 8'h96; B = 8'h5F; #100;
A = 8'h96; B = 8'h60; #100;
A = 8'h96; B = 8'h61; #100;
A = 8'h96; B = 8'h62; #100;
A = 8'h96; B = 8'h63; #100;
A = 8'h96; B = 8'h64; #100;
A = 8'h96; B = 8'h65; #100;
A = 8'h96; B = 8'h66; #100;
A = 8'h96; B = 8'h67; #100;
A = 8'h96; B = 8'h68; #100;
A = 8'h96; B = 8'h69; #100;
A = 8'h96; B = 8'h6A; #100;
A = 8'h96; B = 8'h6B; #100;
A = 8'h96; B = 8'h6C; #100;
A = 8'h96; B = 8'h6D; #100;
A = 8'h96; B = 8'h6E; #100;
A = 8'h96; B = 8'h6F; #100;
A = 8'h96; B = 8'h70; #100;
A = 8'h96; B = 8'h71; #100;
A = 8'h96; B = 8'h72; #100;
A = 8'h96; B = 8'h73; #100;
A = 8'h96; B = 8'h74; #100;
A = 8'h96; B = 8'h75; #100;
A = 8'h96; B = 8'h76; #100;
A = 8'h96; B = 8'h77; #100;
A = 8'h96; B = 8'h78; #100;
A = 8'h96; B = 8'h79; #100;
A = 8'h96; B = 8'h7A; #100;
A = 8'h96; B = 8'h7B; #100;
A = 8'h96; B = 8'h7C; #100;
A = 8'h96; B = 8'h7D; #100;
A = 8'h96; B = 8'h7E; #100;
A = 8'h96; B = 8'h7F; #100;
A = 8'h96; B = 8'h80; #100;
A = 8'h96; B = 8'h81; #100;
A = 8'h96; B = 8'h82; #100;
A = 8'h96; B = 8'h83; #100;
A = 8'h96; B = 8'h84; #100;
A = 8'h96; B = 8'h85; #100;
A = 8'h96; B = 8'h86; #100;
A = 8'h96; B = 8'h87; #100;
A = 8'h96; B = 8'h88; #100;
A = 8'h96; B = 8'h89; #100;
A = 8'h96; B = 8'h8A; #100;
A = 8'h96; B = 8'h8B; #100;
A = 8'h96; B = 8'h8C; #100;
A = 8'h96; B = 8'h8D; #100;
A = 8'h96; B = 8'h8E; #100;
A = 8'h96; B = 8'h8F; #100;
A = 8'h96; B = 8'h90; #100;
A = 8'h96; B = 8'h91; #100;
A = 8'h96; B = 8'h92; #100;
A = 8'h96; B = 8'h93; #100;
A = 8'h96; B = 8'h94; #100;
A = 8'h96; B = 8'h95; #100;
A = 8'h96; B = 8'h96; #100;
A = 8'h96; B = 8'h97; #100;
A = 8'h96; B = 8'h98; #100;
A = 8'h96; B = 8'h99; #100;
A = 8'h96; B = 8'h9A; #100;
A = 8'h96; B = 8'h9B; #100;
A = 8'h96; B = 8'h9C; #100;
A = 8'h96; B = 8'h9D; #100;
A = 8'h96; B = 8'h9E; #100;
A = 8'h96; B = 8'h9F; #100;
A = 8'h96; B = 8'hA0; #100;
A = 8'h96; B = 8'hA1; #100;
A = 8'h96; B = 8'hA2; #100;
A = 8'h96; B = 8'hA3; #100;
A = 8'h96; B = 8'hA4; #100;
A = 8'h96; B = 8'hA5; #100;
A = 8'h96; B = 8'hA6; #100;
A = 8'h96; B = 8'hA7; #100;
A = 8'h96; B = 8'hA8; #100;
A = 8'h96; B = 8'hA9; #100;
A = 8'h96; B = 8'hAA; #100;
A = 8'h96; B = 8'hAB; #100;
A = 8'h96; B = 8'hAC; #100;
A = 8'h96; B = 8'hAD; #100;
A = 8'h96; B = 8'hAE; #100;
A = 8'h96; B = 8'hAF; #100;
A = 8'h96; B = 8'hB0; #100;
A = 8'h96; B = 8'hB1; #100;
A = 8'h96; B = 8'hB2; #100;
A = 8'h96; B = 8'hB3; #100;
A = 8'h96; B = 8'hB4; #100;
A = 8'h96; B = 8'hB5; #100;
A = 8'h96; B = 8'hB6; #100;
A = 8'h96; B = 8'hB7; #100;
A = 8'h96; B = 8'hB8; #100;
A = 8'h96; B = 8'hB9; #100;
A = 8'h96; B = 8'hBA; #100;
A = 8'h96; B = 8'hBB; #100;
A = 8'h96; B = 8'hBC; #100;
A = 8'h96; B = 8'hBD; #100;
A = 8'h96; B = 8'hBE; #100;
A = 8'h96; B = 8'hBF; #100;
A = 8'h96; B = 8'hC0; #100;
A = 8'h96; B = 8'hC1; #100;
A = 8'h96; B = 8'hC2; #100;
A = 8'h96; B = 8'hC3; #100;
A = 8'h96; B = 8'hC4; #100;
A = 8'h96; B = 8'hC5; #100;
A = 8'h96; B = 8'hC6; #100;
A = 8'h96; B = 8'hC7; #100;
A = 8'h96; B = 8'hC8; #100;
A = 8'h96; B = 8'hC9; #100;
A = 8'h96; B = 8'hCA; #100;
A = 8'h96; B = 8'hCB; #100;
A = 8'h96; B = 8'hCC; #100;
A = 8'h96; B = 8'hCD; #100;
A = 8'h96; B = 8'hCE; #100;
A = 8'h96; B = 8'hCF; #100;
A = 8'h96; B = 8'hD0; #100;
A = 8'h96; B = 8'hD1; #100;
A = 8'h96; B = 8'hD2; #100;
A = 8'h96; B = 8'hD3; #100;
A = 8'h96; B = 8'hD4; #100;
A = 8'h96; B = 8'hD5; #100;
A = 8'h96; B = 8'hD6; #100;
A = 8'h96; B = 8'hD7; #100;
A = 8'h96; B = 8'hD8; #100;
A = 8'h96; B = 8'hD9; #100;
A = 8'h96; B = 8'hDA; #100;
A = 8'h96; B = 8'hDB; #100;
A = 8'h96; B = 8'hDC; #100;
A = 8'h96; B = 8'hDD; #100;
A = 8'h96; B = 8'hDE; #100;
A = 8'h96; B = 8'hDF; #100;
A = 8'h96; B = 8'hE0; #100;
A = 8'h96; B = 8'hE1; #100;
A = 8'h96; B = 8'hE2; #100;
A = 8'h96; B = 8'hE3; #100;
A = 8'h96; B = 8'hE4; #100;
A = 8'h96; B = 8'hE5; #100;
A = 8'h96; B = 8'hE6; #100;
A = 8'h96; B = 8'hE7; #100;
A = 8'h96; B = 8'hE8; #100;
A = 8'h96; B = 8'hE9; #100;
A = 8'h96; B = 8'hEA; #100;
A = 8'h96; B = 8'hEB; #100;
A = 8'h96; B = 8'hEC; #100;
A = 8'h96; B = 8'hED; #100;
A = 8'h96; B = 8'hEE; #100;
A = 8'h96; B = 8'hEF; #100;
A = 8'h96; B = 8'hF0; #100;
A = 8'h96; B = 8'hF1; #100;
A = 8'h96; B = 8'hF2; #100;
A = 8'h96; B = 8'hF3; #100;
A = 8'h96; B = 8'hF4; #100;
A = 8'h96; B = 8'hF5; #100;
A = 8'h96; B = 8'hF6; #100;
A = 8'h96; B = 8'hF7; #100;
A = 8'h96; B = 8'hF8; #100;
A = 8'h96; B = 8'hF9; #100;
A = 8'h96; B = 8'hFA; #100;
A = 8'h96; B = 8'hFB; #100;
A = 8'h96; B = 8'hFC; #100;
A = 8'h96; B = 8'hFD; #100;
A = 8'h96; B = 8'hFE; #100;
A = 8'h96; B = 8'hFF; #100;
A = 8'h97; B = 8'h0; #100;
A = 8'h97; B = 8'h1; #100;
A = 8'h97; B = 8'h2; #100;
A = 8'h97; B = 8'h3; #100;
A = 8'h97; B = 8'h4; #100;
A = 8'h97; B = 8'h5; #100;
A = 8'h97; B = 8'h6; #100;
A = 8'h97; B = 8'h7; #100;
A = 8'h97; B = 8'h8; #100;
A = 8'h97; B = 8'h9; #100;
A = 8'h97; B = 8'hA; #100;
A = 8'h97; B = 8'hB; #100;
A = 8'h97; B = 8'hC; #100;
A = 8'h97; B = 8'hD; #100;
A = 8'h97; B = 8'hE; #100;
A = 8'h97; B = 8'hF; #100;
A = 8'h97; B = 8'h10; #100;
A = 8'h97; B = 8'h11; #100;
A = 8'h97; B = 8'h12; #100;
A = 8'h97; B = 8'h13; #100;
A = 8'h97; B = 8'h14; #100;
A = 8'h97; B = 8'h15; #100;
A = 8'h97; B = 8'h16; #100;
A = 8'h97; B = 8'h17; #100;
A = 8'h97; B = 8'h18; #100;
A = 8'h97; B = 8'h19; #100;
A = 8'h97; B = 8'h1A; #100;
A = 8'h97; B = 8'h1B; #100;
A = 8'h97; B = 8'h1C; #100;
A = 8'h97; B = 8'h1D; #100;
A = 8'h97; B = 8'h1E; #100;
A = 8'h97; B = 8'h1F; #100;
A = 8'h97; B = 8'h20; #100;
A = 8'h97; B = 8'h21; #100;
A = 8'h97; B = 8'h22; #100;
A = 8'h97; B = 8'h23; #100;
A = 8'h97; B = 8'h24; #100;
A = 8'h97; B = 8'h25; #100;
A = 8'h97; B = 8'h26; #100;
A = 8'h97; B = 8'h27; #100;
A = 8'h97; B = 8'h28; #100;
A = 8'h97; B = 8'h29; #100;
A = 8'h97; B = 8'h2A; #100;
A = 8'h97; B = 8'h2B; #100;
A = 8'h97; B = 8'h2C; #100;
A = 8'h97; B = 8'h2D; #100;
A = 8'h97; B = 8'h2E; #100;
A = 8'h97; B = 8'h2F; #100;
A = 8'h97; B = 8'h30; #100;
A = 8'h97; B = 8'h31; #100;
A = 8'h97; B = 8'h32; #100;
A = 8'h97; B = 8'h33; #100;
A = 8'h97; B = 8'h34; #100;
A = 8'h97; B = 8'h35; #100;
A = 8'h97; B = 8'h36; #100;
A = 8'h97; B = 8'h37; #100;
A = 8'h97; B = 8'h38; #100;
A = 8'h97; B = 8'h39; #100;
A = 8'h97; B = 8'h3A; #100;
A = 8'h97; B = 8'h3B; #100;
A = 8'h97; B = 8'h3C; #100;
A = 8'h97; B = 8'h3D; #100;
A = 8'h97; B = 8'h3E; #100;
A = 8'h97; B = 8'h3F; #100;
A = 8'h97; B = 8'h40; #100;
A = 8'h97; B = 8'h41; #100;
A = 8'h97; B = 8'h42; #100;
A = 8'h97; B = 8'h43; #100;
A = 8'h97; B = 8'h44; #100;
A = 8'h97; B = 8'h45; #100;
A = 8'h97; B = 8'h46; #100;
A = 8'h97; B = 8'h47; #100;
A = 8'h97; B = 8'h48; #100;
A = 8'h97; B = 8'h49; #100;
A = 8'h97; B = 8'h4A; #100;
A = 8'h97; B = 8'h4B; #100;
A = 8'h97; B = 8'h4C; #100;
A = 8'h97; B = 8'h4D; #100;
A = 8'h97; B = 8'h4E; #100;
A = 8'h97; B = 8'h4F; #100;
A = 8'h97; B = 8'h50; #100;
A = 8'h97; B = 8'h51; #100;
A = 8'h97; B = 8'h52; #100;
A = 8'h97; B = 8'h53; #100;
A = 8'h97; B = 8'h54; #100;
A = 8'h97; B = 8'h55; #100;
A = 8'h97; B = 8'h56; #100;
A = 8'h97; B = 8'h57; #100;
A = 8'h97; B = 8'h58; #100;
A = 8'h97; B = 8'h59; #100;
A = 8'h97; B = 8'h5A; #100;
A = 8'h97; B = 8'h5B; #100;
A = 8'h97; B = 8'h5C; #100;
A = 8'h97; B = 8'h5D; #100;
A = 8'h97; B = 8'h5E; #100;
A = 8'h97; B = 8'h5F; #100;
A = 8'h97; B = 8'h60; #100;
A = 8'h97; B = 8'h61; #100;
A = 8'h97; B = 8'h62; #100;
A = 8'h97; B = 8'h63; #100;
A = 8'h97; B = 8'h64; #100;
A = 8'h97; B = 8'h65; #100;
A = 8'h97; B = 8'h66; #100;
A = 8'h97; B = 8'h67; #100;
A = 8'h97; B = 8'h68; #100;
A = 8'h97; B = 8'h69; #100;
A = 8'h97; B = 8'h6A; #100;
A = 8'h97; B = 8'h6B; #100;
A = 8'h97; B = 8'h6C; #100;
A = 8'h97; B = 8'h6D; #100;
A = 8'h97; B = 8'h6E; #100;
A = 8'h97; B = 8'h6F; #100;
A = 8'h97; B = 8'h70; #100;
A = 8'h97; B = 8'h71; #100;
A = 8'h97; B = 8'h72; #100;
A = 8'h97; B = 8'h73; #100;
A = 8'h97; B = 8'h74; #100;
A = 8'h97; B = 8'h75; #100;
A = 8'h97; B = 8'h76; #100;
A = 8'h97; B = 8'h77; #100;
A = 8'h97; B = 8'h78; #100;
A = 8'h97; B = 8'h79; #100;
A = 8'h97; B = 8'h7A; #100;
A = 8'h97; B = 8'h7B; #100;
A = 8'h97; B = 8'h7C; #100;
A = 8'h97; B = 8'h7D; #100;
A = 8'h97; B = 8'h7E; #100;
A = 8'h97; B = 8'h7F; #100;
A = 8'h97; B = 8'h80; #100;
A = 8'h97; B = 8'h81; #100;
A = 8'h97; B = 8'h82; #100;
A = 8'h97; B = 8'h83; #100;
A = 8'h97; B = 8'h84; #100;
A = 8'h97; B = 8'h85; #100;
A = 8'h97; B = 8'h86; #100;
A = 8'h97; B = 8'h87; #100;
A = 8'h97; B = 8'h88; #100;
A = 8'h97; B = 8'h89; #100;
A = 8'h97; B = 8'h8A; #100;
A = 8'h97; B = 8'h8B; #100;
A = 8'h97; B = 8'h8C; #100;
A = 8'h97; B = 8'h8D; #100;
A = 8'h97; B = 8'h8E; #100;
A = 8'h97; B = 8'h8F; #100;
A = 8'h97; B = 8'h90; #100;
A = 8'h97; B = 8'h91; #100;
A = 8'h97; B = 8'h92; #100;
A = 8'h97; B = 8'h93; #100;
A = 8'h97; B = 8'h94; #100;
A = 8'h97; B = 8'h95; #100;
A = 8'h97; B = 8'h96; #100;
A = 8'h97; B = 8'h97; #100;
A = 8'h97; B = 8'h98; #100;
A = 8'h97; B = 8'h99; #100;
A = 8'h97; B = 8'h9A; #100;
A = 8'h97; B = 8'h9B; #100;
A = 8'h97; B = 8'h9C; #100;
A = 8'h97; B = 8'h9D; #100;
A = 8'h97; B = 8'h9E; #100;
A = 8'h97; B = 8'h9F; #100;
A = 8'h97; B = 8'hA0; #100;
A = 8'h97; B = 8'hA1; #100;
A = 8'h97; B = 8'hA2; #100;
A = 8'h97; B = 8'hA3; #100;
A = 8'h97; B = 8'hA4; #100;
A = 8'h97; B = 8'hA5; #100;
A = 8'h97; B = 8'hA6; #100;
A = 8'h97; B = 8'hA7; #100;
A = 8'h97; B = 8'hA8; #100;
A = 8'h97; B = 8'hA9; #100;
A = 8'h97; B = 8'hAA; #100;
A = 8'h97; B = 8'hAB; #100;
A = 8'h97; B = 8'hAC; #100;
A = 8'h97; B = 8'hAD; #100;
A = 8'h97; B = 8'hAE; #100;
A = 8'h97; B = 8'hAF; #100;
A = 8'h97; B = 8'hB0; #100;
A = 8'h97; B = 8'hB1; #100;
A = 8'h97; B = 8'hB2; #100;
A = 8'h97; B = 8'hB3; #100;
A = 8'h97; B = 8'hB4; #100;
A = 8'h97; B = 8'hB5; #100;
A = 8'h97; B = 8'hB6; #100;
A = 8'h97; B = 8'hB7; #100;
A = 8'h97; B = 8'hB8; #100;
A = 8'h97; B = 8'hB9; #100;
A = 8'h97; B = 8'hBA; #100;
A = 8'h97; B = 8'hBB; #100;
A = 8'h97; B = 8'hBC; #100;
A = 8'h97; B = 8'hBD; #100;
A = 8'h97; B = 8'hBE; #100;
A = 8'h97; B = 8'hBF; #100;
A = 8'h97; B = 8'hC0; #100;
A = 8'h97; B = 8'hC1; #100;
A = 8'h97; B = 8'hC2; #100;
A = 8'h97; B = 8'hC3; #100;
A = 8'h97; B = 8'hC4; #100;
A = 8'h97; B = 8'hC5; #100;
A = 8'h97; B = 8'hC6; #100;
A = 8'h97; B = 8'hC7; #100;
A = 8'h97; B = 8'hC8; #100;
A = 8'h97; B = 8'hC9; #100;
A = 8'h97; B = 8'hCA; #100;
A = 8'h97; B = 8'hCB; #100;
A = 8'h97; B = 8'hCC; #100;
A = 8'h97; B = 8'hCD; #100;
A = 8'h97; B = 8'hCE; #100;
A = 8'h97; B = 8'hCF; #100;
A = 8'h97; B = 8'hD0; #100;
A = 8'h97; B = 8'hD1; #100;
A = 8'h97; B = 8'hD2; #100;
A = 8'h97; B = 8'hD3; #100;
A = 8'h97; B = 8'hD4; #100;
A = 8'h97; B = 8'hD5; #100;
A = 8'h97; B = 8'hD6; #100;
A = 8'h97; B = 8'hD7; #100;
A = 8'h97; B = 8'hD8; #100;
A = 8'h97; B = 8'hD9; #100;
A = 8'h97; B = 8'hDA; #100;
A = 8'h97; B = 8'hDB; #100;
A = 8'h97; B = 8'hDC; #100;
A = 8'h97; B = 8'hDD; #100;
A = 8'h97; B = 8'hDE; #100;
A = 8'h97; B = 8'hDF; #100;
A = 8'h97; B = 8'hE0; #100;
A = 8'h97; B = 8'hE1; #100;
A = 8'h97; B = 8'hE2; #100;
A = 8'h97; B = 8'hE3; #100;
A = 8'h97; B = 8'hE4; #100;
A = 8'h97; B = 8'hE5; #100;
A = 8'h97; B = 8'hE6; #100;
A = 8'h97; B = 8'hE7; #100;
A = 8'h97; B = 8'hE8; #100;
A = 8'h97; B = 8'hE9; #100;
A = 8'h97; B = 8'hEA; #100;
A = 8'h97; B = 8'hEB; #100;
A = 8'h97; B = 8'hEC; #100;
A = 8'h97; B = 8'hED; #100;
A = 8'h97; B = 8'hEE; #100;
A = 8'h97; B = 8'hEF; #100;
A = 8'h97; B = 8'hF0; #100;
A = 8'h97; B = 8'hF1; #100;
A = 8'h97; B = 8'hF2; #100;
A = 8'h97; B = 8'hF3; #100;
A = 8'h97; B = 8'hF4; #100;
A = 8'h97; B = 8'hF5; #100;
A = 8'h97; B = 8'hF6; #100;
A = 8'h97; B = 8'hF7; #100;
A = 8'h97; B = 8'hF8; #100;
A = 8'h97; B = 8'hF9; #100;
A = 8'h97; B = 8'hFA; #100;
A = 8'h97; B = 8'hFB; #100;
A = 8'h97; B = 8'hFC; #100;
A = 8'h97; B = 8'hFD; #100;
A = 8'h97; B = 8'hFE; #100;
A = 8'h97; B = 8'hFF; #100;
A = 8'h98; B = 8'h0; #100;
A = 8'h98; B = 8'h1; #100;
A = 8'h98; B = 8'h2; #100;
A = 8'h98; B = 8'h3; #100;
A = 8'h98; B = 8'h4; #100;
A = 8'h98; B = 8'h5; #100;
A = 8'h98; B = 8'h6; #100;
A = 8'h98; B = 8'h7; #100;
A = 8'h98; B = 8'h8; #100;
A = 8'h98; B = 8'h9; #100;
A = 8'h98; B = 8'hA; #100;
A = 8'h98; B = 8'hB; #100;
A = 8'h98; B = 8'hC; #100;
A = 8'h98; B = 8'hD; #100;
A = 8'h98; B = 8'hE; #100;
A = 8'h98; B = 8'hF; #100;
A = 8'h98; B = 8'h10; #100;
A = 8'h98; B = 8'h11; #100;
A = 8'h98; B = 8'h12; #100;
A = 8'h98; B = 8'h13; #100;
A = 8'h98; B = 8'h14; #100;
A = 8'h98; B = 8'h15; #100;
A = 8'h98; B = 8'h16; #100;
A = 8'h98; B = 8'h17; #100;
A = 8'h98; B = 8'h18; #100;
A = 8'h98; B = 8'h19; #100;
A = 8'h98; B = 8'h1A; #100;
A = 8'h98; B = 8'h1B; #100;
A = 8'h98; B = 8'h1C; #100;
A = 8'h98; B = 8'h1D; #100;
A = 8'h98; B = 8'h1E; #100;
A = 8'h98; B = 8'h1F; #100;
A = 8'h98; B = 8'h20; #100;
A = 8'h98; B = 8'h21; #100;
A = 8'h98; B = 8'h22; #100;
A = 8'h98; B = 8'h23; #100;
A = 8'h98; B = 8'h24; #100;
A = 8'h98; B = 8'h25; #100;
A = 8'h98; B = 8'h26; #100;
A = 8'h98; B = 8'h27; #100;
A = 8'h98; B = 8'h28; #100;
A = 8'h98; B = 8'h29; #100;
A = 8'h98; B = 8'h2A; #100;
A = 8'h98; B = 8'h2B; #100;
A = 8'h98; B = 8'h2C; #100;
A = 8'h98; B = 8'h2D; #100;
A = 8'h98; B = 8'h2E; #100;
A = 8'h98; B = 8'h2F; #100;
A = 8'h98; B = 8'h30; #100;
A = 8'h98; B = 8'h31; #100;
A = 8'h98; B = 8'h32; #100;
A = 8'h98; B = 8'h33; #100;
A = 8'h98; B = 8'h34; #100;
A = 8'h98; B = 8'h35; #100;
A = 8'h98; B = 8'h36; #100;
A = 8'h98; B = 8'h37; #100;
A = 8'h98; B = 8'h38; #100;
A = 8'h98; B = 8'h39; #100;
A = 8'h98; B = 8'h3A; #100;
A = 8'h98; B = 8'h3B; #100;
A = 8'h98; B = 8'h3C; #100;
A = 8'h98; B = 8'h3D; #100;
A = 8'h98; B = 8'h3E; #100;
A = 8'h98; B = 8'h3F; #100;
A = 8'h98; B = 8'h40; #100;
A = 8'h98; B = 8'h41; #100;
A = 8'h98; B = 8'h42; #100;
A = 8'h98; B = 8'h43; #100;
A = 8'h98; B = 8'h44; #100;
A = 8'h98; B = 8'h45; #100;
A = 8'h98; B = 8'h46; #100;
A = 8'h98; B = 8'h47; #100;
A = 8'h98; B = 8'h48; #100;
A = 8'h98; B = 8'h49; #100;
A = 8'h98; B = 8'h4A; #100;
A = 8'h98; B = 8'h4B; #100;
A = 8'h98; B = 8'h4C; #100;
A = 8'h98; B = 8'h4D; #100;
A = 8'h98; B = 8'h4E; #100;
A = 8'h98; B = 8'h4F; #100;
A = 8'h98; B = 8'h50; #100;
A = 8'h98; B = 8'h51; #100;
A = 8'h98; B = 8'h52; #100;
A = 8'h98; B = 8'h53; #100;
A = 8'h98; B = 8'h54; #100;
A = 8'h98; B = 8'h55; #100;
A = 8'h98; B = 8'h56; #100;
A = 8'h98; B = 8'h57; #100;
A = 8'h98; B = 8'h58; #100;
A = 8'h98; B = 8'h59; #100;
A = 8'h98; B = 8'h5A; #100;
A = 8'h98; B = 8'h5B; #100;
A = 8'h98; B = 8'h5C; #100;
A = 8'h98; B = 8'h5D; #100;
A = 8'h98; B = 8'h5E; #100;
A = 8'h98; B = 8'h5F; #100;
A = 8'h98; B = 8'h60; #100;
A = 8'h98; B = 8'h61; #100;
A = 8'h98; B = 8'h62; #100;
A = 8'h98; B = 8'h63; #100;
A = 8'h98; B = 8'h64; #100;
A = 8'h98; B = 8'h65; #100;
A = 8'h98; B = 8'h66; #100;
A = 8'h98; B = 8'h67; #100;
A = 8'h98; B = 8'h68; #100;
A = 8'h98; B = 8'h69; #100;
A = 8'h98; B = 8'h6A; #100;
A = 8'h98; B = 8'h6B; #100;
A = 8'h98; B = 8'h6C; #100;
A = 8'h98; B = 8'h6D; #100;
A = 8'h98; B = 8'h6E; #100;
A = 8'h98; B = 8'h6F; #100;
A = 8'h98; B = 8'h70; #100;
A = 8'h98; B = 8'h71; #100;
A = 8'h98; B = 8'h72; #100;
A = 8'h98; B = 8'h73; #100;
A = 8'h98; B = 8'h74; #100;
A = 8'h98; B = 8'h75; #100;
A = 8'h98; B = 8'h76; #100;
A = 8'h98; B = 8'h77; #100;
A = 8'h98; B = 8'h78; #100;
A = 8'h98; B = 8'h79; #100;
A = 8'h98; B = 8'h7A; #100;
A = 8'h98; B = 8'h7B; #100;
A = 8'h98; B = 8'h7C; #100;
A = 8'h98; B = 8'h7D; #100;
A = 8'h98; B = 8'h7E; #100;
A = 8'h98; B = 8'h7F; #100;
A = 8'h98; B = 8'h80; #100;
A = 8'h98; B = 8'h81; #100;
A = 8'h98; B = 8'h82; #100;
A = 8'h98; B = 8'h83; #100;
A = 8'h98; B = 8'h84; #100;
A = 8'h98; B = 8'h85; #100;
A = 8'h98; B = 8'h86; #100;
A = 8'h98; B = 8'h87; #100;
A = 8'h98; B = 8'h88; #100;
A = 8'h98; B = 8'h89; #100;
A = 8'h98; B = 8'h8A; #100;
A = 8'h98; B = 8'h8B; #100;
A = 8'h98; B = 8'h8C; #100;
A = 8'h98; B = 8'h8D; #100;
A = 8'h98; B = 8'h8E; #100;
A = 8'h98; B = 8'h8F; #100;
A = 8'h98; B = 8'h90; #100;
A = 8'h98; B = 8'h91; #100;
A = 8'h98; B = 8'h92; #100;
A = 8'h98; B = 8'h93; #100;
A = 8'h98; B = 8'h94; #100;
A = 8'h98; B = 8'h95; #100;
A = 8'h98; B = 8'h96; #100;
A = 8'h98; B = 8'h97; #100;
A = 8'h98; B = 8'h98; #100;
A = 8'h98; B = 8'h99; #100;
A = 8'h98; B = 8'h9A; #100;
A = 8'h98; B = 8'h9B; #100;
A = 8'h98; B = 8'h9C; #100;
A = 8'h98; B = 8'h9D; #100;
A = 8'h98; B = 8'h9E; #100;
A = 8'h98; B = 8'h9F; #100;
A = 8'h98; B = 8'hA0; #100;
A = 8'h98; B = 8'hA1; #100;
A = 8'h98; B = 8'hA2; #100;
A = 8'h98; B = 8'hA3; #100;
A = 8'h98; B = 8'hA4; #100;
A = 8'h98; B = 8'hA5; #100;
A = 8'h98; B = 8'hA6; #100;
A = 8'h98; B = 8'hA7; #100;
A = 8'h98; B = 8'hA8; #100;
A = 8'h98; B = 8'hA9; #100;
A = 8'h98; B = 8'hAA; #100;
A = 8'h98; B = 8'hAB; #100;
A = 8'h98; B = 8'hAC; #100;
A = 8'h98; B = 8'hAD; #100;
A = 8'h98; B = 8'hAE; #100;
A = 8'h98; B = 8'hAF; #100;
A = 8'h98; B = 8'hB0; #100;
A = 8'h98; B = 8'hB1; #100;
A = 8'h98; B = 8'hB2; #100;
A = 8'h98; B = 8'hB3; #100;
A = 8'h98; B = 8'hB4; #100;
A = 8'h98; B = 8'hB5; #100;
A = 8'h98; B = 8'hB6; #100;
A = 8'h98; B = 8'hB7; #100;
A = 8'h98; B = 8'hB8; #100;
A = 8'h98; B = 8'hB9; #100;
A = 8'h98; B = 8'hBA; #100;
A = 8'h98; B = 8'hBB; #100;
A = 8'h98; B = 8'hBC; #100;
A = 8'h98; B = 8'hBD; #100;
A = 8'h98; B = 8'hBE; #100;
A = 8'h98; B = 8'hBF; #100;
A = 8'h98; B = 8'hC0; #100;
A = 8'h98; B = 8'hC1; #100;
A = 8'h98; B = 8'hC2; #100;
A = 8'h98; B = 8'hC3; #100;
A = 8'h98; B = 8'hC4; #100;
A = 8'h98; B = 8'hC5; #100;
A = 8'h98; B = 8'hC6; #100;
A = 8'h98; B = 8'hC7; #100;
A = 8'h98; B = 8'hC8; #100;
A = 8'h98; B = 8'hC9; #100;
A = 8'h98; B = 8'hCA; #100;
A = 8'h98; B = 8'hCB; #100;
A = 8'h98; B = 8'hCC; #100;
A = 8'h98; B = 8'hCD; #100;
A = 8'h98; B = 8'hCE; #100;
A = 8'h98; B = 8'hCF; #100;
A = 8'h98; B = 8'hD0; #100;
A = 8'h98; B = 8'hD1; #100;
A = 8'h98; B = 8'hD2; #100;
A = 8'h98; B = 8'hD3; #100;
A = 8'h98; B = 8'hD4; #100;
A = 8'h98; B = 8'hD5; #100;
A = 8'h98; B = 8'hD6; #100;
A = 8'h98; B = 8'hD7; #100;
A = 8'h98; B = 8'hD8; #100;
A = 8'h98; B = 8'hD9; #100;
A = 8'h98; B = 8'hDA; #100;
A = 8'h98; B = 8'hDB; #100;
A = 8'h98; B = 8'hDC; #100;
A = 8'h98; B = 8'hDD; #100;
A = 8'h98; B = 8'hDE; #100;
A = 8'h98; B = 8'hDF; #100;
A = 8'h98; B = 8'hE0; #100;
A = 8'h98; B = 8'hE1; #100;
A = 8'h98; B = 8'hE2; #100;
A = 8'h98; B = 8'hE3; #100;
A = 8'h98; B = 8'hE4; #100;
A = 8'h98; B = 8'hE5; #100;
A = 8'h98; B = 8'hE6; #100;
A = 8'h98; B = 8'hE7; #100;
A = 8'h98; B = 8'hE8; #100;
A = 8'h98; B = 8'hE9; #100;
A = 8'h98; B = 8'hEA; #100;
A = 8'h98; B = 8'hEB; #100;
A = 8'h98; B = 8'hEC; #100;
A = 8'h98; B = 8'hED; #100;
A = 8'h98; B = 8'hEE; #100;
A = 8'h98; B = 8'hEF; #100;
A = 8'h98; B = 8'hF0; #100;
A = 8'h98; B = 8'hF1; #100;
A = 8'h98; B = 8'hF2; #100;
A = 8'h98; B = 8'hF3; #100;
A = 8'h98; B = 8'hF4; #100;
A = 8'h98; B = 8'hF5; #100;
A = 8'h98; B = 8'hF6; #100;
A = 8'h98; B = 8'hF7; #100;
A = 8'h98; B = 8'hF8; #100;
A = 8'h98; B = 8'hF9; #100;
A = 8'h98; B = 8'hFA; #100;
A = 8'h98; B = 8'hFB; #100;
A = 8'h98; B = 8'hFC; #100;
A = 8'h98; B = 8'hFD; #100;
A = 8'h98; B = 8'hFE; #100;
A = 8'h98; B = 8'hFF; #100;
A = 8'h99; B = 8'h0; #100;
A = 8'h99; B = 8'h1; #100;
A = 8'h99; B = 8'h2; #100;
A = 8'h99; B = 8'h3; #100;
A = 8'h99; B = 8'h4; #100;
A = 8'h99; B = 8'h5; #100;
A = 8'h99; B = 8'h6; #100;
A = 8'h99; B = 8'h7; #100;
A = 8'h99; B = 8'h8; #100;
A = 8'h99; B = 8'h9; #100;
A = 8'h99; B = 8'hA; #100;
A = 8'h99; B = 8'hB; #100;
A = 8'h99; B = 8'hC; #100;
A = 8'h99; B = 8'hD; #100;
A = 8'h99; B = 8'hE; #100;
A = 8'h99; B = 8'hF; #100;
A = 8'h99; B = 8'h10; #100;
A = 8'h99; B = 8'h11; #100;
A = 8'h99; B = 8'h12; #100;
A = 8'h99; B = 8'h13; #100;
A = 8'h99; B = 8'h14; #100;
A = 8'h99; B = 8'h15; #100;
A = 8'h99; B = 8'h16; #100;
A = 8'h99; B = 8'h17; #100;
A = 8'h99; B = 8'h18; #100;
A = 8'h99; B = 8'h19; #100;
A = 8'h99; B = 8'h1A; #100;
A = 8'h99; B = 8'h1B; #100;
A = 8'h99; B = 8'h1C; #100;
A = 8'h99; B = 8'h1D; #100;
A = 8'h99; B = 8'h1E; #100;
A = 8'h99; B = 8'h1F; #100;
A = 8'h99; B = 8'h20; #100;
A = 8'h99; B = 8'h21; #100;
A = 8'h99; B = 8'h22; #100;
A = 8'h99; B = 8'h23; #100;
A = 8'h99; B = 8'h24; #100;
A = 8'h99; B = 8'h25; #100;
A = 8'h99; B = 8'h26; #100;
A = 8'h99; B = 8'h27; #100;
A = 8'h99; B = 8'h28; #100;
A = 8'h99; B = 8'h29; #100;
A = 8'h99; B = 8'h2A; #100;
A = 8'h99; B = 8'h2B; #100;
A = 8'h99; B = 8'h2C; #100;
A = 8'h99; B = 8'h2D; #100;
A = 8'h99; B = 8'h2E; #100;
A = 8'h99; B = 8'h2F; #100;
A = 8'h99; B = 8'h30; #100;
A = 8'h99; B = 8'h31; #100;
A = 8'h99; B = 8'h32; #100;
A = 8'h99; B = 8'h33; #100;
A = 8'h99; B = 8'h34; #100;
A = 8'h99; B = 8'h35; #100;
A = 8'h99; B = 8'h36; #100;
A = 8'h99; B = 8'h37; #100;
A = 8'h99; B = 8'h38; #100;
A = 8'h99; B = 8'h39; #100;
A = 8'h99; B = 8'h3A; #100;
A = 8'h99; B = 8'h3B; #100;
A = 8'h99; B = 8'h3C; #100;
A = 8'h99; B = 8'h3D; #100;
A = 8'h99; B = 8'h3E; #100;
A = 8'h99; B = 8'h3F; #100;
A = 8'h99; B = 8'h40; #100;
A = 8'h99; B = 8'h41; #100;
A = 8'h99; B = 8'h42; #100;
A = 8'h99; B = 8'h43; #100;
A = 8'h99; B = 8'h44; #100;
A = 8'h99; B = 8'h45; #100;
A = 8'h99; B = 8'h46; #100;
A = 8'h99; B = 8'h47; #100;
A = 8'h99; B = 8'h48; #100;
A = 8'h99; B = 8'h49; #100;
A = 8'h99; B = 8'h4A; #100;
A = 8'h99; B = 8'h4B; #100;
A = 8'h99; B = 8'h4C; #100;
A = 8'h99; B = 8'h4D; #100;
A = 8'h99; B = 8'h4E; #100;
A = 8'h99; B = 8'h4F; #100;
A = 8'h99; B = 8'h50; #100;
A = 8'h99; B = 8'h51; #100;
A = 8'h99; B = 8'h52; #100;
A = 8'h99; B = 8'h53; #100;
A = 8'h99; B = 8'h54; #100;
A = 8'h99; B = 8'h55; #100;
A = 8'h99; B = 8'h56; #100;
A = 8'h99; B = 8'h57; #100;
A = 8'h99; B = 8'h58; #100;
A = 8'h99; B = 8'h59; #100;
A = 8'h99; B = 8'h5A; #100;
A = 8'h99; B = 8'h5B; #100;
A = 8'h99; B = 8'h5C; #100;
A = 8'h99; B = 8'h5D; #100;
A = 8'h99; B = 8'h5E; #100;
A = 8'h99; B = 8'h5F; #100;
A = 8'h99; B = 8'h60; #100;
A = 8'h99; B = 8'h61; #100;
A = 8'h99; B = 8'h62; #100;
A = 8'h99; B = 8'h63; #100;
A = 8'h99; B = 8'h64; #100;
A = 8'h99; B = 8'h65; #100;
A = 8'h99; B = 8'h66; #100;
A = 8'h99; B = 8'h67; #100;
A = 8'h99; B = 8'h68; #100;
A = 8'h99; B = 8'h69; #100;
A = 8'h99; B = 8'h6A; #100;
A = 8'h99; B = 8'h6B; #100;
A = 8'h99; B = 8'h6C; #100;
A = 8'h99; B = 8'h6D; #100;
A = 8'h99; B = 8'h6E; #100;
A = 8'h99; B = 8'h6F; #100;
A = 8'h99; B = 8'h70; #100;
A = 8'h99; B = 8'h71; #100;
A = 8'h99; B = 8'h72; #100;
A = 8'h99; B = 8'h73; #100;
A = 8'h99; B = 8'h74; #100;
A = 8'h99; B = 8'h75; #100;
A = 8'h99; B = 8'h76; #100;
A = 8'h99; B = 8'h77; #100;
A = 8'h99; B = 8'h78; #100;
A = 8'h99; B = 8'h79; #100;
A = 8'h99; B = 8'h7A; #100;
A = 8'h99; B = 8'h7B; #100;
A = 8'h99; B = 8'h7C; #100;
A = 8'h99; B = 8'h7D; #100;
A = 8'h99; B = 8'h7E; #100;
A = 8'h99; B = 8'h7F; #100;
A = 8'h99; B = 8'h80; #100;
A = 8'h99; B = 8'h81; #100;
A = 8'h99; B = 8'h82; #100;
A = 8'h99; B = 8'h83; #100;
A = 8'h99; B = 8'h84; #100;
A = 8'h99; B = 8'h85; #100;
A = 8'h99; B = 8'h86; #100;
A = 8'h99; B = 8'h87; #100;
A = 8'h99; B = 8'h88; #100;
A = 8'h99; B = 8'h89; #100;
A = 8'h99; B = 8'h8A; #100;
A = 8'h99; B = 8'h8B; #100;
A = 8'h99; B = 8'h8C; #100;
A = 8'h99; B = 8'h8D; #100;
A = 8'h99; B = 8'h8E; #100;
A = 8'h99; B = 8'h8F; #100;
A = 8'h99; B = 8'h90; #100;
A = 8'h99; B = 8'h91; #100;
A = 8'h99; B = 8'h92; #100;
A = 8'h99; B = 8'h93; #100;
A = 8'h99; B = 8'h94; #100;
A = 8'h99; B = 8'h95; #100;
A = 8'h99; B = 8'h96; #100;
A = 8'h99; B = 8'h97; #100;
A = 8'h99; B = 8'h98; #100;
A = 8'h99; B = 8'h99; #100;
A = 8'h99; B = 8'h9A; #100;
A = 8'h99; B = 8'h9B; #100;
A = 8'h99; B = 8'h9C; #100;
A = 8'h99; B = 8'h9D; #100;
A = 8'h99; B = 8'h9E; #100;
A = 8'h99; B = 8'h9F; #100;
A = 8'h99; B = 8'hA0; #100;
A = 8'h99; B = 8'hA1; #100;
A = 8'h99; B = 8'hA2; #100;
A = 8'h99; B = 8'hA3; #100;
A = 8'h99; B = 8'hA4; #100;
A = 8'h99; B = 8'hA5; #100;
A = 8'h99; B = 8'hA6; #100;
A = 8'h99; B = 8'hA7; #100;
A = 8'h99; B = 8'hA8; #100;
A = 8'h99; B = 8'hA9; #100;
A = 8'h99; B = 8'hAA; #100;
A = 8'h99; B = 8'hAB; #100;
A = 8'h99; B = 8'hAC; #100;
A = 8'h99; B = 8'hAD; #100;
A = 8'h99; B = 8'hAE; #100;
A = 8'h99; B = 8'hAF; #100;
A = 8'h99; B = 8'hB0; #100;
A = 8'h99; B = 8'hB1; #100;
A = 8'h99; B = 8'hB2; #100;
A = 8'h99; B = 8'hB3; #100;
A = 8'h99; B = 8'hB4; #100;
A = 8'h99; B = 8'hB5; #100;
A = 8'h99; B = 8'hB6; #100;
A = 8'h99; B = 8'hB7; #100;
A = 8'h99; B = 8'hB8; #100;
A = 8'h99; B = 8'hB9; #100;
A = 8'h99; B = 8'hBA; #100;
A = 8'h99; B = 8'hBB; #100;
A = 8'h99; B = 8'hBC; #100;
A = 8'h99; B = 8'hBD; #100;
A = 8'h99; B = 8'hBE; #100;
A = 8'h99; B = 8'hBF; #100;
A = 8'h99; B = 8'hC0; #100;
A = 8'h99; B = 8'hC1; #100;
A = 8'h99; B = 8'hC2; #100;
A = 8'h99; B = 8'hC3; #100;
A = 8'h99; B = 8'hC4; #100;
A = 8'h99; B = 8'hC5; #100;
A = 8'h99; B = 8'hC6; #100;
A = 8'h99; B = 8'hC7; #100;
A = 8'h99; B = 8'hC8; #100;
A = 8'h99; B = 8'hC9; #100;
A = 8'h99; B = 8'hCA; #100;
A = 8'h99; B = 8'hCB; #100;
A = 8'h99; B = 8'hCC; #100;
A = 8'h99; B = 8'hCD; #100;
A = 8'h99; B = 8'hCE; #100;
A = 8'h99; B = 8'hCF; #100;
A = 8'h99; B = 8'hD0; #100;
A = 8'h99; B = 8'hD1; #100;
A = 8'h99; B = 8'hD2; #100;
A = 8'h99; B = 8'hD3; #100;
A = 8'h99; B = 8'hD4; #100;
A = 8'h99; B = 8'hD5; #100;
A = 8'h99; B = 8'hD6; #100;
A = 8'h99; B = 8'hD7; #100;
A = 8'h99; B = 8'hD8; #100;
A = 8'h99; B = 8'hD9; #100;
A = 8'h99; B = 8'hDA; #100;
A = 8'h99; B = 8'hDB; #100;
A = 8'h99; B = 8'hDC; #100;
A = 8'h99; B = 8'hDD; #100;
A = 8'h99; B = 8'hDE; #100;
A = 8'h99; B = 8'hDF; #100;
A = 8'h99; B = 8'hE0; #100;
A = 8'h99; B = 8'hE1; #100;
A = 8'h99; B = 8'hE2; #100;
A = 8'h99; B = 8'hE3; #100;
A = 8'h99; B = 8'hE4; #100;
A = 8'h99; B = 8'hE5; #100;
A = 8'h99; B = 8'hE6; #100;
A = 8'h99; B = 8'hE7; #100;
A = 8'h99; B = 8'hE8; #100;
A = 8'h99; B = 8'hE9; #100;
A = 8'h99; B = 8'hEA; #100;
A = 8'h99; B = 8'hEB; #100;
A = 8'h99; B = 8'hEC; #100;
A = 8'h99; B = 8'hED; #100;
A = 8'h99; B = 8'hEE; #100;
A = 8'h99; B = 8'hEF; #100;
A = 8'h99; B = 8'hF0; #100;
A = 8'h99; B = 8'hF1; #100;
A = 8'h99; B = 8'hF2; #100;
A = 8'h99; B = 8'hF3; #100;
A = 8'h99; B = 8'hF4; #100;
A = 8'h99; B = 8'hF5; #100;
A = 8'h99; B = 8'hF6; #100;
A = 8'h99; B = 8'hF7; #100;
A = 8'h99; B = 8'hF8; #100;
A = 8'h99; B = 8'hF9; #100;
A = 8'h99; B = 8'hFA; #100;
A = 8'h99; B = 8'hFB; #100;
A = 8'h99; B = 8'hFC; #100;
A = 8'h99; B = 8'hFD; #100;
A = 8'h99; B = 8'hFE; #100;
A = 8'h99; B = 8'hFF; #100;
A = 8'h9A; B = 8'h0; #100;
A = 8'h9A; B = 8'h1; #100;
A = 8'h9A; B = 8'h2; #100;
A = 8'h9A; B = 8'h3; #100;
A = 8'h9A; B = 8'h4; #100;
A = 8'h9A; B = 8'h5; #100;
A = 8'h9A; B = 8'h6; #100;
A = 8'h9A; B = 8'h7; #100;
A = 8'h9A; B = 8'h8; #100;
A = 8'h9A; B = 8'h9; #100;
A = 8'h9A; B = 8'hA; #100;
A = 8'h9A; B = 8'hB; #100;
A = 8'h9A; B = 8'hC; #100;
A = 8'h9A; B = 8'hD; #100;
A = 8'h9A; B = 8'hE; #100;
A = 8'h9A; B = 8'hF; #100;
A = 8'h9A; B = 8'h10; #100;
A = 8'h9A; B = 8'h11; #100;
A = 8'h9A; B = 8'h12; #100;
A = 8'h9A; B = 8'h13; #100;
A = 8'h9A; B = 8'h14; #100;
A = 8'h9A; B = 8'h15; #100;
A = 8'h9A; B = 8'h16; #100;
A = 8'h9A; B = 8'h17; #100;
A = 8'h9A; B = 8'h18; #100;
A = 8'h9A; B = 8'h19; #100;
A = 8'h9A; B = 8'h1A; #100;
A = 8'h9A; B = 8'h1B; #100;
A = 8'h9A; B = 8'h1C; #100;
A = 8'h9A; B = 8'h1D; #100;
A = 8'h9A; B = 8'h1E; #100;
A = 8'h9A; B = 8'h1F; #100;
A = 8'h9A; B = 8'h20; #100;
A = 8'h9A; B = 8'h21; #100;
A = 8'h9A; B = 8'h22; #100;
A = 8'h9A; B = 8'h23; #100;
A = 8'h9A; B = 8'h24; #100;
A = 8'h9A; B = 8'h25; #100;
A = 8'h9A; B = 8'h26; #100;
A = 8'h9A; B = 8'h27; #100;
A = 8'h9A; B = 8'h28; #100;
A = 8'h9A; B = 8'h29; #100;
A = 8'h9A; B = 8'h2A; #100;
A = 8'h9A; B = 8'h2B; #100;
A = 8'h9A; B = 8'h2C; #100;
A = 8'h9A; B = 8'h2D; #100;
A = 8'h9A; B = 8'h2E; #100;
A = 8'h9A; B = 8'h2F; #100;
A = 8'h9A; B = 8'h30; #100;
A = 8'h9A; B = 8'h31; #100;
A = 8'h9A; B = 8'h32; #100;
A = 8'h9A; B = 8'h33; #100;
A = 8'h9A; B = 8'h34; #100;
A = 8'h9A; B = 8'h35; #100;
A = 8'h9A; B = 8'h36; #100;
A = 8'h9A; B = 8'h37; #100;
A = 8'h9A; B = 8'h38; #100;
A = 8'h9A; B = 8'h39; #100;
A = 8'h9A; B = 8'h3A; #100;
A = 8'h9A; B = 8'h3B; #100;
A = 8'h9A; B = 8'h3C; #100;
A = 8'h9A; B = 8'h3D; #100;
A = 8'h9A; B = 8'h3E; #100;
A = 8'h9A; B = 8'h3F; #100;
A = 8'h9A; B = 8'h40; #100;
A = 8'h9A; B = 8'h41; #100;
A = 8'h9A; B = 8'h42; #100;
A = 8'h9A; B = 8'h43; #100;
A = 8'h9A; B = 8'h44; #100;
A = 8'h9A; B = 8'h45; #100;
A = 8'h9A; B = 8'h46; #100;
A = 8'h9A; B = 8'h47; #100;
A = 8'h9A; B = 8'h48; #100;
A = 8'h9A; B = 8'h49; #100;
A = 8'h9A; B = 8'h4A; #100;
A = 8'h9A; B = 8'h4B; #100;
A = 8'h9A; B = 8'h4C; #100;
A = 8'h9A; B = 8'h4D; #100;
A = 8'h9A; B = 8'h4E; #100;
A = 8'h9A; B = 8'h4F; #100;
A = 8'h9A; B = 8'h50; #100;
A = 8'h9A; B = 8'h51; #100;
A = 8'h9A; B = 8'h52; #100;
A = 8'h9A; B = 8'h53; #100;
A = 8'h9A; B = 8'h54; #100;
A = 8'h9A; B = 8'h55; #100;
A = 8'h9A; B = 8'h56; #100;
A = 8'h9A; B = 8'h57; #100;
A = 8'h9A; B = 8'h58; #100;
A = 8'h9A; B = 8'h59; #100;
A = 8'h9A; B = 8'h5A; #100;
A = 8'h9A; B = 8'h5B; #100;
A = 8'h9A; B = 8'h5C; #100;
A = 8'h9A; B = 8'h5D; #100;
A = 8'h9A; B = 8'h5E; #100;
A = 8'h9A; B = 8'h5F; #100;
A = 8'h9A; B = 8'h60; #100;
A = 8'h9A; B = 8'h61; #100;
A = 8'h9A; B = 8'h62; #100;
A = 8'h9A; B = 8'h63; #100;
A = 8'h9A; B = 8'h64; #100;
A = 8'h9A; B = 8'h65; #100;
A = 8'h9A; B = 8'h66; #100;
A = 8'h9A; B = 8'h67; #100;
A = 8'h9A; B = 8'h68; #100;
A = 8'h9A; B = 8'h69; #100;
A = 8'h9A; B = 8'h6A; #100;
A = 8'h9A; B = 8'h6B; #100;
A = 8'h9A; B = 8'h6C; #100;
A = 8'h9A; B = 8'h6D; #100;
A = 8'h9A; B = 8'h6E; #100;
A = 8'h9A; B = 8'h6F; #100;
A = 8'h9A; B = 8'h70; #100;
A = 8'h9A; B = 8'h71; #100;
A = 8'h9A; B = 8'h72; #100;
A = 8'h9A; B = 8'h73; #100;
A = 8'h9A; B = 8'h74; #100;
A = 8'h9A; B = 8'h75; #100;
A = 8'h9A; B = 8'h76; #100;
A = 8'h9A; B = 8'h77; #100;
A = 8'h9A; B = 8'h78; #100;
A = 8'h9A; B = 8'h79; #100;
A = 8'h9A; B = 8'h7A; #100;
A = 8'h9A; B = 8'h7B; #100;
A = 8'h9A; B = 8'h7C; #100;
A = 8'h9A; B = 8'h7D; #100;
A = 8'h9A; B = 8'h7E; #100;
A = 8'h9A; B = 8'h7F; #100;
A = 8'h9A; B = 8'h80; #100;
A = 8'h9A; B = 8'h81; #100;
A = 8'h9A; B = 8'h82; #100;
A = 8'h9A; B = 8'h83; #100;
A = 8'h9A; B = 8'h84; #100;
A = 8'h9A; B = 8'h85; #100;
A = 8'h9A; B = 8'h86; #100;
A = 8'h9A; B = 8'h87; #100;
A = 8'h9A; B = 8'h88; #100;
A = 8'h9A; B = 8'h89; #100;
A = 8'h9A; B = 8'h8A; #100;
A = 8'h9A; B = 8'h8B; #100;
A = 8'h9A; B = 8'h8C; #100;
A = 8'h9A; B = 8'h8D; #100;
A = 8'h9A; B = 8'h8E; #100;
A = 8'h9A; B = 8'h8F; #100;
A = 8'h9A; B = 8'h90; #100;
A = 8'h9A; B = 8'h91; #100;
A = 8'h9A; B = 8'h92; #100;
A = 8'h9A; B = 8'h93; #100;
A = 8'h9A; B = 8'h94; #100;
A = 8'h9A; B = 8'h95; #100;
A = 8'h9A; B = 8'h96; #100;
A = 8'h9A; B = 8'h97; #100;
A = 8'h9A; B = 8'h98; #100;
A = 8'h9A; B = 8'h99; #100;
A = 8'h9A; B = 8'h9A; #100;
A = 8'h9A; B = 8'h9B; #100;
A = 8'h9A; B = 8'h9C; #100;
A = 8'h9A; B = 8'h9D; #100;
A = 8'h9A; B = 8'h9E; #100;
A = 8'h9A; B = 8'h9F; #100;
A = 8'h9A; B = 8'hA0; #100;
A = 8'h9A; B = 8'hA1; #100;
A = 8'h9A; B = 8'hA2; #100;
A = 8'h9A; B = 8'hA3; #100;
A = 8'h9A; B = 8'hA4; #100;
A = 8'h9A; B = 8'hA5; #100;
A = 8'h9A; B = 8'hA6; #100;
A = 8'h9A; B = 8'hA7; #100;
A = 8'h9A; B = 8'hA8; #100;
A = 8'h9A; B = 8'hA9; #100;
A = 8'h9A; B = 8'hAA; #100;
A = 8'h9A; B = 8'hAB; #100;
A = 8'h9A; B = 8'hAC; #100;
A = 8'h9A; B = 8'hAD; #100;
A = 8'h9A; B = 8'hAE; #100;
A = 8'h9A; B = 8'hAF; #100;
A = 8'h9A; B = 8'hB0; #100;
A = 8'h9A; B = 8'hB1; #100;
A = 8'h9A; B = 8'hB2; #100;
A = 8'h9A; B = 8'hB3; #100;
A = 8'h9A; B = 8'hB4; #100;
A = 8'h9A; B = 8'hB5; #100;
A = 8'h9A; B = 8'hB6; #100;
A = 8'h9A; B = 8'hB7; #100;
A = 8'h9A; B = 8'hB8; #100;
A = 8'h9A; B = 8'hB9; #100;
A = 8'h9A; B = 8'hBA; #100;
A = 8'h9A; B = 8'hBB; #100;
A = 8'h9A; B = 8'hBC; #100;
A = 8'h9A; B = 8'hBD; #100;
A = 8'h9A; B = 8'hBE; #100;
A = 8'h9A; B = 8'hBF; #100;
A = 8'h9A; B = 8'hC0; #100;
A = 8'h9A; B = 8'hC1; #100;
A = 8'h9A; B = 8'hC2; #100;
A = 8'h9A; B = 8'hC3; #100;
A = 8'h9A; B = 8'hC4; #100;
A = 8'h9A; B = 8'hC5; #100;
A = 8'h9A; B = 8'hC6; #100;
A = 8'h9A; B = 8'hC7; #100;
A = 8'h9A; B = 8'hC8; #100;
A = 8'h9A; B = 8'hC9; #100;
A = 8'h9A; B = 8'hCA; #100;
A = 8'h9A; B = 8'hCB; #100;
A = 8'h9A; B = 8'hCC; #100;
A = 8'h9A; B = 8'hCD; #100;
A = 8'h9A; B = 8'hCE; #100;
A = 8'h9A; B = 8'hCF; #100;
A = 8'h9A; B = 8'hD0; #100;
A = 8'h9A; B = 8'hD1; #100;
A = 8'h9A; B = 8'hD2; #100;
A = 8'h9A; B = 8'hD3; #100;
A = 8'h9A; B = 8'hD4; #100;
A = 8'h9A; B = 8'hD5; #100;
A = 8'h9A; B = 8'hD6; #100;
A = 8'h9A; B = 8'hD7; #100;
A = 8'h9A; B = 8'hD8; #100;
A = 8'h9A; B = 8'hD9; #100;
A = 8'h9A; B = 8'hDA; #100;
A = 8'h9A; B = 8'hDB; #100;
A = 8'h9A; B = 8'hDC; #100;
A = 8'h9A; B = 8'hDD; #100;
A = 8'h9A; B = 8'hDE; #100;
A = 8'h9A; B = 8'hDF; #100;
A = 8'h9A; B = 8'hE0; #100;
A = 8'h9A; B = 8'hE1; #100;
A = 8'h9A; B = 8'hE2; #100;
A = 8'h9A; B = 8'hE3; #100;
A = 8'h9A; B = 8'hE4; #100;
A = 8'h9A; B = 8'hE5; #100;
A = 8'h9A; B = 8'hE6; #100;
A = 8'h9A; B = 8'hE7; #100;
A = 8'h9A; B = 8'hE8; #100;
A = 8'h9A; B = 8'hE9; #100;
A = 8'h9A; B = 8'hEA; #100;
A = 8'h9A; B = 8'hEB; #100;
A = 8'h9A; B = 8'hEC; #100;
A = 8'h9A; B = 8'hED; #100;
A = 8'h9A; B = 8'hEE; #100;
A = 8'h9A; B = 8'hEF; #100;
A = 8'h9A; B = 8'hF0; #100;
A = 8'h9A; B = 8'hF1; #100;
A = 8'h9A; B = 8'hF2; #100;
A = 8'h9A; B = 8'hF3; #100;
A = 8'h9A; B = 8'hF4; #100;
A = 8'h9A; B = 8'hF5; #100;
A = 8'h9A; B = 8'hF6; #100;
A = 8'h9A; B = 8'hF7; #100;
A = 8'h9A; B = 8'hF8; #100;
A = 8'h9A; B = 8'hF9; #100;
A = 8'h9A; B = 8'hFA; #100;
A = 8'h9A; B = 8'hFB; #100;
A = 8'h9A; B = 8'hFC; #100;
A = 8'h9A; B = 8'hFD; #100;
A = 8'h9A; B = 8'hFE; #100;
A = 8'h9A; B = 8'hFF; #100;
A = 8'h9B; B = 8'h0; #100;
A = 8'h9B; B = 8'h1; #100;
A = 8'h9B; B = 8'h2; #100;
A = 8'h9B; B = 8'h3; #100;
A = 8'h9B; B = 8'h4; #100;
A = 8'h9B; B = 8'h5; #100;
A = 8'h9B; B = 8'h6; #100;
A = 8'h9B; B = 8'h7; #100;
A = 8'h9B; B = 8'h8; #100;
A = 8'h9B; B = 8'h9; #100;
A = 8'h9B; B = 8'hA; #100;
A = 8'h9B; B = 8'hB; #100;
A = 8'h9B; B = 8'hC; #100;
A = 8'h9B; B = 8'hD; #100;
A = 8'h9B; B = 8'hE; #100;
A = 8'h9B; B = 8'hF; #100;
A = 8'h9B; B = 8'h10; #100;
A = 8'h9B; B = 8'h11; #100;
A = 8'h9B; B = 8'h12; #100;
A = 8'h9B; B = 8'h13; #100;
A = 8'h9B; B = 8'h14; #100;
A = 8'h9B; B = 8'h15; #100;
A = 8'h9B; B = 8'h16; #100;
A = 8'h9B; B = 8'h17; #100;
A = 8'h9B; B = 8'h18; #100;
A = 8'h9B; B = 8'h19; #100;
A = 8'h9B; B = 8'h1A; #100;
A = 8'h9B; B = 8'h1B; #100;
A = 8'h9B; B = 8'h1C; #100;
A = 8'h9B; B = 8'h1D; #100;
A = 8'h9B; B = 8'h1E; #100;
A = 8'h9B; B = 8'h1F; #100;
A = 8'h9B; B = 8'h20; #100;
A = 8'h9B; B = 8'h21; #100;
A = 8'h9B; B = 8'h22; #100;
A = 8'h9B; B = 8'h23; #100;
A = 8'h9B; B = 8'h24; #100;
A = 8'h9B; B = 8'h25; #100;
A = 8'h9B; B = 8'h26; #100;
A = 8'h9B; B = 8'h27; #100;
A = 8'h9B; B = 8'h28; #100;
A = 8'h9B; B = 8'h29; #100;
A = 8'h9B; B = 8'h2A; #100;
A = 8'h9B; B = 8'h2B; #100;
A = 8'h9B; B = 8'h2C; #100;
A = 8'h9B; B = 8'h2D; #100;
A = 8'h9B; B = 8'h2E; #100;
A = 8'h9B; B = 8'h2F; #100;
A = 8'h9B; B = 8'h30; #100;
A = 8'h9B; B = 8'h31; #100;
A = 8'h9B; B = 8'h32; #100;
A = 8'h9B; B = 8'h33; #100;
A = 8'h9B; B = 8'h34; #100;
A = 8'h9B; B = 8'h35; #100;
A = 8'h9B; B = 8'h36; #100;
A = 8'h9B; B = 8'h37; #100;
A = 8'h9B; B = 8'h38; #100;
A = 8'h9B; B = 8'h39; #100;
A = 8'h9B; B = 8'h3A; #100;
A = 8'h9B; B = 8'h3B; #100;
A = 8'h9B; B = 8'h3C; #100;
A = 8'h9B; B = 8'h3D; #100;
A = 8'h9B; B = 8'h3E; #100;
A = 8'h9B; B = 8'h3F; #100;
A = 8'h9B; B = 8'h40; #100;
A = 8'h9B; B = 8'h41; #100;
A = 8'h9B; B = 8'h42; #100;
A = 8'h9B; B = 8'h43; #100;
A = 8'h9B; B = 8'h44; #100;
A = 8'h9B; B = 8'h45; #100;
A = 8'h9B; B = 8'h46; #100;
A = 8'h9B; B = 8'h47; #100;
A = 8'h9B; B = 8'h48; #100;
A = 8'h9B; B = 8'h49; #100;
A = 8'h9B; B = 8'h4A; #100;
A = 8'h9B; B = 8'h4B; #100;
A = 8'h9B; B = 8'h4C; #100;
A = 8'h9B; B = 8'h4D; #100;
A = 8'h9B; B = 8'h4E; #100;
A = 8'h9B; B = 8'h4F; #100;
A = 8'h9B; B = 8'h50; #100;
A = 8'h9B; B = 8'h51; #100;
A = 8'h9B; B = 8'h52; #100;
A = 8'h9B; B = 8'h53; #100;
A = 8'h9B; B = 8'h54; #100;
A = 8'h9B; B = 8'h55; #100;
A = 8'h9B; B = 8'h56; #100;
A = 8'h9B; B = 8'h57; #100;
A = 8'h9B; B = 8'h58; #100;
A = 8'h9B; B = 8'h59; #100;
A = 8'h9B; B = 8'h5A; #100;
A = 8'h9B; B = 8'h5B; #100;
A = 8'h9B; B = 8'h5C; #100;
A = 8'h9B; B = 8'h5D; #100;
A = 8'h9B; B = 8'h5E; #100;
A = 8'h9B; B = 8'h5F; #100;
A = 8'h9B; B = 8'h60; #100;
A = 8'h9B; B = 8'h61; #100;
A = 8'h9B; B = 8'h62; #100;
A = 8'h9B; B = 8'h63; #100;
A = 8'h9B; B = 8'h64; #100;
A = 8'h9B; B = 8'h65; #100;
A = 8'h9B; B = 8'h66; #100;
A = 8'h9B; B = 8'h67; #100;
A = 8'h9B; B = 8'h68; #100;
A = 8'h9B; B = 8'h69; #100;
A = 8'h9B; B = 8'h6A; #100;
A = 8'h9B; B = 8'h6B; #100;
A = 8'h9B; B = 8'h6C; #100;
A = 8'h9B; B = 8'h6D; #100;
A = 8'h9B; B = 8'h6E; #100;
A = 8'h9B; B = 8'h6F; #100;
A = 8'h9B; B = 8'h70; #100;
A = 8'h9B; B = 8'h71; #100;
A = 8'h9B; B = 8'h72; #100;
A = 8'h9B; B = 8'h73; #100;
A = 8'h9B; B = 8'h74; #100;
A = 8'h9B; B = 8'h75; #100;
A = 8'h9B; B = 8'h76; #100;
A = 8'h9B; B = 8'h77; #100;
A = 8'h9B; B = 8'h78; #100;
A = 8'h9B; B = 8'h79; #100;
A = 8'h9B; B = 8'h7A; #100;
A = 8'h9B; B = 8'h7B; #100;
A = 8'h9B; B = 8'h7C; #100;
A = 8'h9B; B = 8'h7D; #100;
A = 8'h9B; B = 8'h7E; #100;
A = 8'h9B; B = 8'h7F; #100;
A = 8'h9B; B = 8'h80; #100;
A = 8'h9B; B = 8'h81; #100;
A = 8'h9B; B = 8'h82; #100;
A = 8'h9B; B = 8'h83; #100;
A = 8'h9B; B = 8'h84; #100;
A = 8'h9B; B = 8'h85; #100;
A = 8'h9B; B = 8'h86; #100;
A = 8'h9B; B = 8'h87; #100;
A = 8'h9B; B = 8'h88; #100;
A = 8'h9B; B = 8'h89; #100;
A = 8'h9B; B = 8'h8A; #100;
A = 8'h9B; B = 8'h8B; #100;
A = 8'h9B; B = 8'h8C; #100;
A = 8'h9B; B = 8'h8D; #100;
A = 8'h9B; B = 8'h8E; #100;
A = 8'h9B; B = 8'h8F; #100;
A = 8'h9B; B = 8'h90; #100;
A = 8'h9B; B = 8'h91; #100;
A = 8'h9B; B = 8'h92; #100;
A = 8'h9B; B = 8'h93; #100;
A = 8'h9B; B = 8'h94; #100;
A = 8'h9B; B = 8'h95; #100;
A = 8'h9B; B = 8'h96; #100;
A = 8'h9B; B = 8'h97; #100;
A = 8'h9B; B = 8'h98; #100;
A = 8'h9B; B = 8'h99; #100;
A = 8'h9B; B = 8'h9A; #100;
A = 8'h9B; B = 8'h9B; #100;
A = 8'h9B; B = 8'h9C; #100;
A = 8'h9B; B = 8'h9D; #100;
A = 8'h9B; B = 8'h9E; #100;
A = 8'h9B; B = 8'h9F; #100;
A = 8'h9B; B = 8'hA0; #100;
A = 8'h9B; B = 8'hA1; #100;
A = 8'h9B; B = 8'hA2; #100;
A = 8'h9B; B = 8'hA3; #100;
A = 8'h9B; B = 8'hA4; #100;
A = 8'h9B; B = 8'hA5; #100;
A = 8'h9B; B = 8'hA6; #100;
A = 8'h9B; B = 8'hA7; #100;
A = 8'h9B; B = 8'hA8; #100;
A = 8'h9B; B = 8'hA9; #100;
A = 8'h9B; B = 8'hAA; #100;
A = 8'h9B; B = 8'hAB; #100;
A = 8'h9B; B = 8'hAC; #100;
A = 8'h9B; B = 8'hAD; #100;
A = 8'h9B; B = 8'hAE; #100;
A = 8'h9B; B = 8'hAF; #100;
A = 8'h9B; B = 8'hB0; #100;
A = 8'h9B; B = 8'hB1; #100;
A = 8'h9B; B = 8'hB2; #100;
A = 8'h9B; B = 8'hB3; #100;
A = 8'h9B; B = 8'hB4; #100;
A = 8'h9B; B = 8'hB5; #100;
A = 8'h9B; B = 8'hB6; #100;
A = 8'h9B; B = 8'hB7; #100;
A = 8'h9B; B = 8'hB8; #100;
A = 8'h9B; B = 8'hB9; #100;
A = 8'h9B; B = 8'hBA; #100;
A = 8'h9B; B = 8'hBB; #100;
A = 8'h9B; B = 8'hBC; #100;
A = 8'h9B; B = 8'hBD; #100;
A = 8'h9B; B = 8'hBE; #100;
A = 8'h9B; B = 8'hBF; #100;
A = 8'h9B; B = 8'hC0; #100;
A = 8'h9B; B = 8'hC1; #100;
A = 8'h9B; B = 8'hC2; #100;
A = 8'h9B; B = 8'hC3; #100;
A = 8'h9B; B = 8'hC4; #100;
A = 8'h9B; B = 8'hC5; #100;
A = 8'h9B; B = 8'hC6; #100;
A = 8'h9B; B = 8'hC7; #100;
A = 8'h9B; B = 8'hC8; #100;
A = 8'h9B; B = 8'hC9; #100;
A = 8'h9B; B = 8'hCA; #100;
A = 8'h9B; B = 8'hCB; #100;
A = 8'h9B; B = 8'hCC; #100;
A = 8'h9B; B = 8'hCD; #100;
A = 8'h9B; B = 8'hCE; #100;
A = 8'h9B; B = 8'hCF; #100;
A = 8'h9B; B = 8'hD0; #100;
A = 8'h9B; B = 8'hD1; #100;
A = 8'h9B; B = 8'hD2; #100;
A = 8'h9B; B = 8'hD3; #100;
A = 8'h9B; B = 8'hD4; #100;
A = 8'h9B; B = 8'hD5; #100;
A = 8'h9B; B = 8'hD6; #100;
A = 8'h9B; B = 8'hD7; #100;
A = 8'h9B; B = 8'hD8; #100;
A = 8'h9B; B = 8'hD9; #100;
A = 8'h9B; B = 8'hDA; #100;
A = 8'h9B; B = 8'hDB; #100;
A = 8'h9B; B = 8'hDC; #100;
A = 8'h9B; B = 8'hDD; #100;
A = 8'h9B; B = 8'hDE; #100;
A = 8'h9B; B = 8'hDF; #100;
A = 8'h9B; B = 8'hE0; #100;
A = 8'h9B; B = 8'hE1; #100;
A = 8'h9B; B = 8'hE2; #100;
A = 8'h9B; B = 8'hE3; #100;
A = 8'h9B; B = 8'hE4; #100;
A = 8'h9B; B = 8'hE5; #100;
A = 8'h9B; B = 8'hE6; #100;
A = 8'h9B; B = 8'hE7; #100;
A = 8'h9B; B = 8'hE8; #100;
A = 8'h9B; B = 8'hE9; #100;
A = 8'h9B; B = 8'hEA; #100;
A = 8'h9B; B = 8'hEB; #100;
A = 8'h9B; B = 8'hEC; #100;
A = 8'h9B; B = 8'hED; #100;
A = 8'h9B; B = 8'hEE; #100;
A = 8'h9B; B = 8'hEF; #100;
A = 8'h9B; B = 8'hF0; #100;
A = 8'h9B; B = 8'hF1; #100;
A = 8'h9B; B = 8'hF2; #100;
A = 8'h9B; B = 8'hF3; #100;
A = 8'h9B; B = 8'hF4; #100;
A = 8'h9B; B = 8'hF5; #100;
A = 8'h9B; B = 8'hF6; #100;
A = 8'h9B; B = 8'hF7; #100;
A = 8'h9B; B = 8'hF8; #100;
A = 8'h9B; B = 8'hF9; #100;
A = 8'h9B; B = 8'hFA; #100;
A = 8'h9B; B = 8'hFB; #100;
A = 8'h9B; B = 8'hFC; #100;
A = 8'h9B; B = 8'hFD; #100;
A = 8'h9B; B = 8'hFE; #100;
A = 8'h9B; B = 8'hFF; #100;
A = 8'h9C; B = 8'h0; #100;
A = 8'h9C; B = 8'h1; #100;
A = 8'h9C; B = 8'h2; #100;
A = 8'h9C; B = 8'h3; #100;
A = 8'h9C; B = 8'h4; #100;
A = 8'h9C; B = 8'h5; #100;
A = 8'h9C; B = 8'h6; #100;
A = 8'h9C; B = 8'h7; #100;
A = 8'h9C; B = 8'h8; #100;
A = 8'h9C; B = 8'h9; #100;
A = 8'h9C; B = 8'hA; #100;
A = 8'h9C; B = 8'hB; #100;
A = 8'h9C; B = 8'hC; #100;
A = 8'h9C; B = 8'hD; #100;
A = 8'h9C; B = 8'hE; #100;
A = 8'h9C; B = 8'hF; #100;
A = 8'h9C; B = 8'h10; #100;
A = 8'h9C; B = 8'h11; #100;
A = 8'h9C; B = 8'h12; #100;
A = 8'h9C; B = 8'h13; #100;
A = 8'h9C; B = 8'h14; #100;
A = 8'h9C; B = 8'h15; #100;
A = 8'h9C; B = 8'h16; #100;
A = 8'h9C; B = 8'h17; #100;
A = 8'h9C; B = 8'h18; #100;
A = 8'h9C; B = 8'h19; #100;
A = 8'h9C; B = 8'h1A; #100;
A = 8'h9C; B = 8'h1B; #100;
A = 8'h9C; B = 8'h1C; #100;
A = 8'h9C; B = 8'h1D; #100;
A = 8'h9C; B = 8'h1E; #100;
A = 8'h9C; B = 8'h1F; #100;
A = 8'h9C; B = 8'h20; #100;
A = 8'h9C; B = 8'h21; #100;
A = 8'h9C; B = 8'h22; #100;
A = 8'h9C; B = 8'h23; #100;
A = 8'h9C; B = 8'h24; #100;
A = 8'h9C; B = 8'h25; #100;
A = 8'h9C; B = 8'h26; #100;
A = 8'h9C; B = 8'h27; #100;
A = 8'h9C; B = 8'h28; #100;
A = 8'h9C; B = 8'h29; #100;
A = 8'h9C; B = 8'h2A; #100;
A = 8'h9C; B = 8'h2B; #100;
A = 8'h9C; B = 8'h2C; #100;
A = 8'h9C; B = 8'h2D; #100;
A = 8'h9C; B = 8'h2E; #100;
A = 8'h9C; B = 8'h2F; #100;
A = 8'h9C; B = 8'h30; #100;
A = 8'h9C; B = 8'h31; #100;
A = 8'h9C; B = 8'h32; #100;
A = 8'h9C; B = 8'h33; #100;
A = 8'h9C; B = 8'h34; #100;
A = 8'h9C; B = 8'h35; #100;
A = 8'h9C; B = 8'h36; #100;
A = 8'h9C; B = 8'h37; #100;
A = 8'h9C; B = 8'h38; #100;
A = 8'h9C; B = 8'h39; #100;
A = 8'h9C; B = 8'h3A; #100;
A = 8'h9C; B = 8'h3B; #100;
A = 8'h9C; B = 8'h3C; #100;
A = 8'h9C; B = 8'h3D; #100;
A = 8'h9C; B = 8'h3E; #100;
A = 8'h9C; B = 8'h3F; #100;
A = 8'h9C; B = 8'h40; #100;
A = 8'h9C; B = 8'h41; #100;
A = 8'h9C; B = 8'h42; #100;
A = 8'h9C; B = 8'h43; #100;
A = 8'h9C; B = 8'h44; #100;
A = 8'h9C; B = 8'h45; #100;
A = 8'h9C; B = 8'h46; #100;
A = 8'h9C; B = 8'h47; #100;
A = 8'h9C; B = 8'h48; #100;
A = 8'h9C; B = 8'h49; #100;
A = 8'h9C; B = 8'h4A; #100;
A = 8'h9C; B = 8'h4B; #100;
A = 8'h9C; B = 8'h4C; #100;
A = 8'h9C; B = 8'h4D; #100;
A = 8'h9C; B = 8'h4E; #100;
A = 8'h9C; B = 8'h4F; #100;
A = 8'h9C; B = 8'h50; #100;
A = 8'h9C; B = 8'h51; #100;
A = 8'h9C; B = 8'h52; #100;
A = 8'h9C; B = 8'h53; #100;
A = 8'h9C; B = 8'h54; #100;
A = 8'h9C; B = 8'h55; #100;
A = 8'h9C; B = 8'h56; #100;
A = 8'h9C; B = 8'h57; #100;
A = 8'h9C; B = 8'h58; #100;
A = 8'h9C; B = 8'h59; #100;
A = 8'h9C; B = 8'h5A; #100;
A = 8'h9C; B = 8'h5B; #100;
A = 8'h9C; B = 8'h5C; #100;
A = 8'h9C; B = 8'h5D; #100;
A = 8'h9C; B = 8'h5E; #100;
A = 8'h9C; B = 8'h5F; #100;
A = 8'h9C; B = 8'h60; #100;
A = 8'h9C; B = 8'h61; #100;
A = 8'h9C; B = 8'h62; #100;
A = 8'h9C; B = 8'h63; #100;
A = 8'h9C; B = 8'h64; #100;
A = 8'h9C; B = 8'h65; #100;
A = 8'h9C; B = 8'h66; #100;
A = 8'h9C; B = 8'h67; #100;
A = 8'h9C; B = 8'h68; #100;
A = 8'h9C; B = 8'h69; #100;
A = 8'h9C; B = 8'h6A; #100;
A = 8'h9C; B = 8'h6B; #100;
A = 8'h9C; B = 8'h6C; #100;
A = 8'h9C; B = 8'h6D; #100;
A = 8'h9C; B = 8'h6E; #100;
A = 8'h9C; B = 8'h6F; #100;
A = 8'h9C; B = 8'h70; #100;
A = 8'h9C; B = 8'h71; #100;
A = 8'h9C; B = 8'h72; #100;
A = 8'h9C; B = 8'h73; #100;
A = 8'h9C; B = 8'h74; #100;
A = 8'h9C; B = 8'h75; #100;
A = 8'h9C; B = 8'h76; #100;
A = 8'h9C; B = 8'h77; #100;
A = 8'h9C; B = 8'h78; #100;
A = 8'h9C; B = 8'h79; #100;
A = 8'h9C; B = 8'h7A; #100;
A = 8'h9C; B = 8'h7B; #100;
A = 8'h9C; B = 8'h7C; #100;
A = 8'h9C; B = 8'h7D; #100;
A = 8'h9C; B = 8'h7E; #100;
A = 8'h9C; B = 8'h7F; #100;
A = 8'h9C; B = 8'h80; #100;
A = 8'h9C; B = 8'h81; #100;
A = 8'h9C; B = 8'h82; #100;
A = 8'h9C; B = 8'h83; #100;
A = 8'h9C; B = 8'h84; #100;
A = 8'h9C; B = 8'h85; #100;
A = 8'h9C; B = 8'h86; #100;
A = 8'h9C; B = 8'h87; #100;
A = 8'h9C; B = 8'h88; #100;
A = 8'h9C; B = 8'h89; #100;
A = 8'h9C; B = 8'h8A; #100;
A = 8'h9C; B = 8'h8B; #100;
A = 8'h9C; B = 8'h8C; #100;
A = 8'h9C; B = 8'h8D; #100;
A = 8'h9C; B = 8'h8E; #100;
A = 8'h9C; B = 8'h8F; #100;
A = 8'h9C; B = 8'h90; #100;
A = 8'h9C; B = 8'h91; #100;
A = 8'h9C; B = 8'h92; #100;
A = 8'h9C; B = 8'h93; #100;
A = 8'h9C; B = 8'h94; #100;
A = 8'h9C; B = 8'h95; #100;
A = 8'h9C; B = 8'h96; #100;
A = 8'h9C; B = 8'h97; #100;
A = 8'h9C; B = 8'h98; #100;
A = 8'h9C; B = 8'h99; #100;
A = 8'h9C; B = 8'h9A; #100;
A = 8'h9C; B = 8'h9B; #100;
A = 8'h9C; B = 8'h9C; #100;
A = 8'h9C; B = 8'h9D; #100;
A = 8'h9C; B = 8'h9E; #100;
A = 8'h9C; B = 8'h9F; #100;
A = 8'h9C; B = 8'hA0; #100;
A = 8'h9C; B = 8'hA1; #100;
A = 8'h9C; B = 8'hA2; #100;
A = 8'h9C; B = 8'hA3; #100;
A = 8'h9C; B = 8'hA4; #100;
A = 8'h9C; B = 8'hA5; #100;
A = 8'h9C; B = 8'hA6; #100;
A = 8'h9C; B = 8'hA7; #100;
A = 8'h9C; B = 8'hA8; #100;
A = 8'h9C; B = 8'hA9; #100;
A = 8'h9C; B = 8'hAA; #100;
A = 8'h9C; B = 8'hAB; #100;
A = 8'h9C; B = 8'hAC; #100;
A = 8'h9C; B = 8'hAD; #100;
A = 8'h9C; B = 8'hAE; #100;
A = 8'h9C; B = 8'hAF; #100;
A = 8'h9C; B = 8'hB0; #100;
A = 8'h9C; B = 8'hB1; #100;
A = 8'h9C; B = 8'hB2; #100;
A = 8'h9C; B = 8'hB3; #100;
A = 8'h9C; B = 8'hB4; #100;
A = 8'h9C; B = 8'hB5; #100;
A = 8'h9C; B = 8'hB6; #100;
A = 8'h9C; B = 8'hB7; #100;
A = 8'h9C; B = 8'hB8; #100;
A = 8'h9C; B = 8'hB9; #100;
A = 8'h9C; B = 8'hBA; #100;
A = 8'h9C; B = 8'hBB; #100;
A = 8'h9C; B = 8'hBC; #100;
A = 8'h9C; B = 8'hBD; #100;
A = 8'h9C; B = 8'hBE; #100;
A = 8'h9C; B = 8'hBF; #100;
A = 8'h9C; B = 8'hC0; #100;
A = 8'h9C; B = 8'hC1; #100;
A = 8'h9C; B = 8'hC2; #100;
A = 8'h9C; B = 8'hC3; #100;
A = 8'h9C; B = 8'hC4; #100;
A = 8'h9C; B = 8'hC5; #100;
A = 8'h9C; B = 8'hC6; #100;
A = 8'h9C; B = 8'hC7; #100;
A = 8'h9C; B = 8'hC8; #100;
A = 8'h9C; B = 8'hC9; #100;
A = 8'h9C; B = 8'hCA; #100;
A = 8'h9C; B = 8'hCB; #100;
A = 8'h9C; B = 8'hCC; #100;
A = 8'h9C; B = 8'hCD; #100;
A = 8'h9C; B = 8'hCE; #100;
A = 8'h9C; B = 8'hCF; #100;
A = 8'h9C; B = 8'hD0; #100;
A = 8'h9C; B = 8'hD1; #100;
A = 8'h9C; B = 8'hD2; #100;
A = 8'h9C; B = 8'hD3; #100;
A = 8'h9C; B = 8'hD4; #100;
A = 8'h9C; B = 8'hD5; #100;
A = 8'h9C; B = 8'hD6; #100;
A = 8'h9C; B = 8'hD7; #100;
A = 8'h9C; B = 8'hD8; #100;
A = 8'h9C; B = 8'hD9; #100;
A = 8'h9C; B = 8'hDA; #100;
A = 8'h9C; B = 8'hDB; #100;
A = 8'h9C; B = 8'hDC; #100;
A = 8'h9C; B = 8'hDD; #100;
A = 8'h9C; B = 8'hDE; #100;
A = 8'h9C; B = 8'hDF; #100;
A = 8'h9C; B = 8'hE0; #100;
A = 8'h9C; B = 8'hE1; #100;
A = 8'h9C; B = 8'hE2; #100;
A = 8'h9C; B = 8'hE3; #100;
A = 8'h9C; B = 8'hE4; #100;
A = 8'h9C; B = 8'hE5; #100;
A = 8'h9C; B = 8'hE6; #100;
A = 8'h9C; B = 8'hE7; #100;
A = 8'h9C; B = 8'hE8; #100;
A = 8'h9C; B = 8'hE9; #100;
A = 8'h9C; B = 8'hEA; #100;
A = 8'h9C; B = 8'hEB; #100;
A = 8'h9C; B = 8'hEC; #100;
A = 8'h9C; B = 8'hED; #100;
A = 8'h9C; B = 8'hEE; #100;
A = 8'h9C; B = 8'hEF; #100;
A = 8'h9C; B = 8'hF0; #100;
A = 8'h9C; B = 8'hF1; #100;
A = 8'h9C; B = 8'hF2; #100;
A = 8'h9C; B = 8'hF3; #100;
A = 8'h9C; B = 8'hF4; #100;
A = 8'h9C; B = 8'hF5; #100;
A = 8'h9C; B = 8'hF6; #100;
A = 8'h9C; B = 8'hF7; #100;
A = 8'h9C; B = 8'hF8; #100;
A = 8'h9C; B = 8'hF9; #100;
A = 8'h9C; B = 8'hFA; #100;
A = 8'h9C; B = 8'hFB; #100;
A = 8'h9C; B = 8'hFC; #100;
A = 8'h9C; B = 8'hFD; #100;
A = 8'h9C; B = 8'hFE; #100;
A = 8'h9C; B = 8'hFF; #100;
A = 8'h9D; B = 8'h0; #100;
A = 8'h9D; B = 8'h1; #100;
A = 8'h9D; B = 8'h2; #100;
A = 8'h9D; B = 8'h3; #100;
A = 8'h9D; B = 8'h4; #100;
A = 8'h9D; B = 8'h5; #100;
A = 8'h9D; B = 8'h6; #100;
A = 8'h9D; B = 8'h7; #100;
A = 8'h9D; B = 8'h8; #100;
A = 8'h9D; B = 8'h9; #100;
A = 8'h9D; B = 8'hA; #100;
A = 8'h9D; B = 8'hB; #100;
A = 8'h9D; B = 8'hC; #100;
A = 8'h9D; B = 8'hD; #100;
A = 8'h9D; B = 8'hE; #100;
A = 8'h9D; B = 8'hF; #100;
A = 8'h9D; B = 8'h10; #100;
A = 8'h9D; B = 8'h11; #100;
A = 8'h9D; B = 8'h12; #100;
A = 8'h9D; B = 8'h13; #100;
A = 8'h9D; B = 8'h14; #100;
A = 8'h9D; B = 8'h15; #100;
A = 8'h9D; B = 8'h16; #100;
A = 8'h9D; B = 8'h17; #100;
A = 8'h9D; B = 8'h18; #100;
A = 8'h9D; B = 8'h19; #100;
A = 8'h9D; B = 8'h1A; #100;
A = 8'h9D; B = 8'h1B; #100;
A = 8'h9D; B = 8'h1C; #100;
A = 8'h9D; B = 8'h1D; #100;
A = 8'h9D; B = 8'h1E; #100;
A = 8'h9D; B = 8'h1F; #100;
A = 8'h9D; B = 8'h20; #100;
A = 8'h9D; B = 8'h21; #100;
A = 8'h9D; B = 8'h22; #100;
A = 8'h9D; B = 8'h23; #100;
A = 8'h9D; B = 8'h24; #100;
A = 8'h9D; B = 8'h25; #100;
A = 8'h9D; B = 8'h26; #100;
A = 8'h9D; B = 8'h27; #100;
A = 8'h9D; B = 8'h28; #100;
A = 8'h9D; B = 8'h29; #100;
A = 8'h9D; B = 8'h2A; #100;
A = 8'h9D; B = 8'h2B; #100;
A = 8'h9D; B = 8'h2C; #100;
A = 8'h9D; B = 8'h2D; #100;
A = 8'h9D; B = 8'h2E; #100;
A = 8'h9D; B = 8'h2F; #100;
A = 8'h9D; B = 8'h30; #100;
A = 8'h9D; B = 8'h31; #100;
A = 8'h9D; B = 8'h32; #100;
A = 8'h9D; B = 8'h33; #100;
A = 8'h9D; B = 8'h34; #100;
A = 8'h9D; B = 8'h35; #100;
A = 8'h9D; B = 8'h36; #100;
A = 8'h9D; B = 8'h37; #100;
A = 8'h9D; B = 8'h38; #100;
A = 8'h9D; B = 8'h39; #100;
A = 8'h9D; B = 8'h3A; #100;
A = 8'h9D; B = 8'h3B; #100;
A = 8'h9D; B = 8'h3C; #100;
A = 8'h9D; B = 8'h3D; #100;
A = 8'h9D; B = 8'h3E; #100;
A = 8'h9D; B = 8'h3F; #100;
A = 8'h9D; B = 8'h40; #100;
A = 8'h9D; B = 8'h41; #100;
A = 8'h9D; B = 8'h42; #100;
A = 8'h9D; B = 8'h43; #100;
A = 8'h9D; B = 8'h44; #100;
A = 8'h9D; B = 8'h45; #100;
A = 8'h9D; B = 8'h46; #100;
A = 8'h9D; B = 8'h47; #100;
A = 8'h9D; B = 8'h48; #100;
A = 8'h9D; B = 8'h49; #100;
A = 8'h9D; B = 8'h4A; #100;
A = 8'h9D; B = 8'h4B; #100;
A = 8'h9D; B = 8'h4C; #100;
A = 8'h9D; B = 8'h4D; #100;
A = 8'h9D; B = 8'h4E; #100;
A = 8'h9D; B = 8'h4F; #100;
A = 8'h9D; B = 8'h50; #100;
A = 8'h9D; B = 8'h51; #100;
A = 8'h9D; B = 8'h52; #100;
A = 8'h9D; B = 8'h53; #100;
A = 8'h9D; B = 8'h54; #100;
A = 8'h9D; B = 8'h55; #100;
A = 8'h9D; B = 8'h56; #100;
A = 8'h9D; B = 8'h57; #100;
A = 8'h9D; B = 8'h58; #100;
A = 8'h9D; B = 8'h59; #100;
A = 8'h9D; B = 8'h5A; #100;
A = 8'h9D; B = 8'h5B; #100;
A = 8'h9D; B = 8'h5C; #100;
A = 8'h9D; B = 8'h5D; #100;
A = 8'h9D; B = 8'h5E; #100;
A = 8'h9D; B = 8'h5F; #100;
A = 8'h9D; B = 8'h60; #100;
A = 8'h9D; B = 8'h61; #100;
A = 8'h9D; B = 8'h62; #100;
A = 8'h9D; B = 8'h63; #100;
A = 8'h9D; B = 8'h64; #100;
A = 8'h9D; B = 8'h65; #100;
A = 8'h9D; B = 8'h66; #100;
A = 8'h9D; B = 8'h67; #100;
A = 8'h9D; B = 8'h68; #100;
A = 8'h9D; B = 8'h69; #100;
A = 8'h9D; B = 8'h6A; #100;
A = 8'h9D; B = 8'h6B; #100;
A = 8'h9D; B = 8'h6C; #100;
A = 8'h9D; B = 8'h6D; #100;
A = 8'h9D; B = 8'h6E; #100;
A = 8'h9D; B = 8'h6F; #100;
A = 8'h9D; B = 8'h70; #100;
A = 8'h9D; B = 8'h71; #100;
A = 8'h9D; B = 8'h72; #100;
A = 8'h9D; B = 8'h73; #100;
A = 8'h9D; B = 8'h74; #100;
A = 8'h9D; B = 8'h75; #100;
A = 8'h9D; B = 8'h76; #100;
A = 8'h9D; B = 8'h77; #100;
A = 8'h9D; B = 8'h78; #100;
A = 8'h9D; B = 8'h79; #100;
A = 8'h9D; B = 8'h7A; #100;
A = 8'h9D; B = 8'h7B; #100;
A = 8'h9D; B = 8'h7C; #100;
A = 8'h9D; B = 8'h7D; #100;
A = 8'h9D; B = 8'h7E; #100;
A = 8'h9D; B = 8'h7F; #100;
A = 8'h9D; B = 8'h80; #100;
A = 8'h9D; B = 8'h81; #100;
A = 8'h9D; B = 8'h82; #100;
A = 8'h9D; B = 8'h83; #100;
A = 8'h9D; B = 8'h84; #100;
A = 8'h9D; B = 8'h85; #100;
A = 8'h9D; B = 8'h86; #100;
A = 8'h9D; B = 8'h87; #100;
A = 8'h9D; B = 8'h88; #100;
A = 8'h9D; B = 8'h89; #100;
A = 8'h9D; B = 8'h8A; #100;
A = 8'h9D; B = 8'h8B; #100;
A = 8'h9D; B = 8'h8C; #100;
A = 8'h9D; B = 8'h8D; #100;
A = 8'h9D; B = 8'h8E; #100;
A = 8'h9D; B = 8'h8F; #100;
A = 8'h9D; B = 8'h90; #100;
A = 8'h9D; B = 8'h91; #100;
A = 8'h9D; B = 8'h92; #100;
A = 8'h9D; B = 8'h93; #100;
A = 8'h9D; B = 8'h94; #100;
A = 8'h9D; B = 8'h95; #100;
A = 8'h9D; B = 8'h96; #100;
A = 8'h9D; B = 8'h97; #100;
A = 8'h9D; B = 8'h98; #100;
A = 8'h9D; B = 8'h99; #100;
A = 8'h9D; B = 8'h9A; #100;
A = 8'h9D; B = 8'h9B; #100;
A = 8'h9D; B = 8'h9C; #100;
A = 8'h9D; B = 8'h9D; #100;
A = 8'h9D; B = 8'h9E; #100;
A = 8'h9D; B = 8'h9F; #100;
A = 8'h9D; B = 8'hA0; #100;
A = 8'h9D; B = 8'hA1; #100;
A = 8'h9D; B = 8'hA2; #100;
A = 8'h9D; B = 8'hA3; #100;
A = 8'h9D; B = 8'hA4; #100;
A = 8'h9D; B = 8'hA5; #100;
A = 8'h9D; B = 8'hA6; #100;
A = 8'h9D; B = 8'hA7; #100;
A = 8'h9D; B = 8'hA8; #100;
A = 8'h9D; B = 8'hA9; #100;
A = 8'h9D; B = 8'hAA; #100;
A = 8'h9D; B = 8'hAB; #100;
A = 8'h9D; B = 8'hAC; #100;
A = 8'h9D; B = 8'hAD; #100;
A = 8'h9D; B = 8'hAE; #100;
A = 8'h9D; B = 8'hAF; #100;
A = 8'h9D; B = 8'hB0; #100;
A = 8'h9D; B = 8'hB1; #100;
A = 8'h9D; B = 8'hB2; #100;
A = 8'h9D; B = 8'hB3; #100;
A = 8'h9D; B = 8'hB4; #100;
A = 8'h9D; B = 8'hB5; #100;
A = 8'h9D; B = 8'hB6; #100;
A = 8'h9D; B = 8'hB7; #100;
A = 8'h9D; B = 8'hB8; #100;
A = 8'h9D; B = 8'hB9; #100;
A = 8'h9D; B = 8'hBA; #100;
A = 8'h9D; B = 8'hBB; #100;
A = 8'h9D; B = 8'hBC; #100;
A = 8'h9D; B = 8'hBD; #100;
A = 8'h9D; B = 8'hBE; #100;
A = 8'h9D; B = 8'hBF; #100;
A = 8'h9D; B = 8'hC0; #100;
A = 8'h9D; B = 8'hC1; #100;
A = 8'h9D; B = 8'hC2; #100;
A = 8'h9D; B = 8'hC3; #100;
A = 8'h9D; B = 8'hC4; #100;
A = 8'h9D; B = 8'hC5; #100;
A = 8'h9D; B = 8'hC6; #100;
A = 8'h9D; B = 8'hC7; #100;
A = 8'h9D; B = 8'hC8; #100;
A = 8'h9D; B = 8'hC9; #100;
A = 8'h9D; B = 8'hCA; #100;
A = 8'h9D; B = 8'hCB; #100;
A = 8'h9D; B = 8'hCC; #100;
A = 8'h9D; B = 8'hCD; #100;
A = 8'h9D; B = 8'hCE; #100;
A = 8'h9D; B = 8'hCF; #100;
A = 8'h9D; B = 8'hD0; #100;
A = 8'h9D; B = 8'hD1; #100;
A = 8'h9D; B = 8'hD2; #100;
A = 8'h9D; B = 8'hD3; #100;
A = 8'h9D; B = 8'hD4; #100;
A = 8'h9D; B = 8'hD5; #100;
A = 8'h9D; B = 8'hD6; #100;
A = 8'h9D; B = 8'hD7; #100;
A = 8'h9D; B = 8'hD8; #100;
A = 8'h9D; B = 8'hD9; #100;
A = 8'h9D; B = 8'hDA; #100;
A = 8'h9D; B = 8'hDB; #100;
A = 8'h9D; B = 8'hDC; #100;
A = 8'h9D; B = 8'hDD; #100;
A = 8'h9D; B = 8'hDE; #100;
A = 8'h9D; B = 8'hDF; #100;
A = 8'h9D; B = 8'hE0; #100;
A = 8'h9D; B = 8'hE1; #100;
A = 8'h9D; B = 8'hE2; #100;
A = 8'h9D; B = 8'hE3; #100;
A = 8'h9D; B = 8'hE4; #100;
A = 8'h9D; B = 8'hE5; #100;
A = 8'h9D; B = 8'hE6; #100;
A = 8'h9D; B = 8'hE7; #100;
A = 8'h9D; B = 8'hE8; #100;
A = 8'h9D; B = 8'hE9; #100;
A = 8'h9D; B = 8'hEA; #100;
A = 8'h9D; B = 8'hEB; #100;
A = 8'h9D; B = 8'hEC; #100;
A = 8'h9D; B = 8'hED; #100;
A = 8'h9D; B = 8'hEE; #100;
A = 8'h9D; B = 8'hEF; #100;
A = 8'h9D; B = 8'hF0; #100;
A = 8'h9D; B = 8'hF1; #100;
A = 8'h9D; B = 8'hF2; #100;
A = 8'h9D; B = 8'hF3; #100;
A = 8'h9D; B = 8'hF4; #100;
A = 8'h9D; B = 8'hF5; #100;
A = 8'h9D; B = 8'hF6; #100;
A = 8'h9D; B = 8'hF7; #100;
A = 8'h9D; B = 8'hF8; #100;
A = 8'h9D; B = 8'hF9; #100;
A = 8'h9D; B = 8'hFA; #100;
A = 8'h9D; B = 8'hFB; #100;
A = 8'h9D; B = 8'hFC; #100;
A = 8'h9D; B = 8'hFD; #100;
A = 8'h9D; B = 8'hFE; #100;
A = 8'h9D; B = 8'hFF; #100;
A = 8'h9E; B = 8'h0; #100;
A = 8'h9E; B = 8'h1; #100;
A = 8'h9E; B = 8'h2; #100;
A = 8'h9E; B = 8'h3; #100;
A = 8'h9E; B = 8'h4; #100;
A = 8'h9E; B = 8'h5; #100;
A = 8'h9E; B = 8'h6; #100;
A = 8'h9E; B = 8'h7; #100;
A = 8'h9E; B = 8'h8; #100;
A = 8'h9E; B = 8'h9; #100;
A = 8'h9E; B = 8'hA; #100;
A = 8'h9E; B = 8'hB; #100;
A = 8'h9E; B = 8'hC; #100;
A = 8'h9E; B = 8'hD; #100;
A = 8'h9E; B = 8'hE; #100;
A = 8'h9E; B = 8'hF; #100;
A = 8'h9E; B = 8'h10; #100;
A = 8'h9E; B = 8'h11; #100;
A = 8'h9E; B = 8'h12; #100;
A = 8'h9E; B = 8'h13; #100;
A = 8'h9E; B = 8'h14; #100;
A = 8'h9E; B = 8'h15; #100;
A = 8'h9E; B = 8'h16; #100;
A = 8'h9E; B = 8'h17; #100;
A = 8'h9E; B = 8'h18; #100;
A = 8'h9E; B = 8'h19; #100;
A = 8'h9E; B = 8'h1A; #100;
A = 8'h9E; B = 8'h1B; #100;
A = 8'h9E; B = 8'h1C; #100;
A = 8'h9E; B = 8'h1D; #100;
A = 8'h9E; B = 8'h1E; #100;
A = 8'h9E; B = 8'h1F; #100;
A = 8'h9E; B = 8'h20; #100;
A = 8'h9E; B = 8'h21; #100;
A = 8'h9E; B = 8'h22; #100;
A = 8'h9E; B = 8'h23; #100;
A = 8'h9E; B = 8'h24; #100;
A = 8'h9E; B = 8'h25; #100;
A = 8'h9E; B = 8'h26; #100;
A = 8'h9E; B = 8'h27; #100;
A = 8'h9E; B = 8'h28; #100;
A = 8'h9E; B = 8'h29; #100;
A = 8'h9E; B = 8'h2A; #100;
A = 8'h9E; B = 8'h2B; #100;
A = 8'h9E; B = 8'h2C; #100;
A = 8'h9E; B = 8'h2D; #100;
A = 8'h9E; B = 8'h2E; #100;
A = 8'h9E; B = 8'h2F; #100;
A = 8'h9E; B = 8'h30; #100;
A = 8'h9E; B = 8'h31; #100;
A = 8'h9E; B = 8'h32; #100;
A = 8'h9E; B = 8'h33; #100;
A = 8'h9E; B = 8'h34; #100;
A = 8'h9E; B = 8'h35; #100;
A = 8'h9E; B = 8'h36; #100;
A = 8'h9E; B = 8'h37; #100;
A = 8'h9E; B = 8'h38; #100;
A = 8'h9E; B = 8'h39; #100;
A = 8'h9E; B = 8'h3A; #100;
A = 8'h9E; B = 8'h3B; #100;
A = 8'h9E; B = 8'h3C; #100;
A = 8'h9E; B = 8'h3D; #100;
A = 8'h9E; B = 8'h3E; #100;
A = 8'h9E; B = 8'h3F; #100;
A = 8'h9E; B = 8'h40; #100;
A = 8'h9E; B = 8'h41; #100;
A = 8'h9E; B = 8'h42; #100;
A = 8'h9E; B = 8'h43; #100;
A = 8'h9E; B = 8'h44; #100;
A = 8'h9E; B = 8'h45; #100;
A = 8'h9E; B = 8'h46; #100;
A = 8'h9E; B = 8'h47; #100;
A = 8'h9E; B = 8'h48; #100;
A = 8'h9E; B = 8'h49; #100;
A = 8'h9E; B = 8'h4A; #100;
A = 8'h9E; B = 8'h4B; #100;
A = 8'h9E; B = 8'h4C; #100;
A = 8'h9E; B = 8'h4D; #100;
A = 8'h9E; B = 8'h4E; #100;
A = 8'h9E; B = 8'h4F; #100;
A = 8'h9E; B = 8'h50; #100;
A = 8'h9E; B = 8'h51; #100;
A = 8'h9E; B = 8'h52; #100;
A = 8'h9E; B = 8'h53; #100;
A = 8'h9E; B = 8'h54; #100;
A = 8'h9E; B = 8'h55; #100;
A = 8'h9E; B = 8'h56; #100;
A = 8'h9E; B = 8'h57; #100;
A = 8'h9E; B = 8'h58; #100;
A = 8'h9E; B = 8'h59; #100;
A = 8'h9E; B = 8'h5A; #100;
A = 8'h9E; B = 8'h5B; #100;
A = 8'h9E; B = 8'h5C; #100;
A = 8'h9E; B = 8'h5D; #100;
A = 8'h9E; B = 8'h5E; #100;
A = 8'h9E; B = 8'h5F; #100;
A = 8'h9E; B = 8'h60; #100;
A = 8'h9E; B = 8'h61; #100;
A = 8'h9E; B = 8'h62; #100;
A = 8'h9E; B = 8'h63; #100;
A = 8'h9E; B = 8'h64; #100;
A = 8'h9E; B = 8'h65; #100;
A = 8'h9E; B = 8'h66; #100;
A = 8'h9E; B = 8'h67; #100;
A = 8'h9E; B = 8'h68; #100;
A = 8'h9E; B = 8'h69; #100;
A = 8'h9E; B = 8'h6A; #100;
A = 8'h9E; B = 8'h6B; #100;
A = 8'h9E; B = 8'h6C; #100;
A = 8'h9E; B = 8'h6D; #100;
A = 8'h9E; B = 8'h6E; #100;
A = 8'h9E; B = 8'h6F; #100;
A = 8'h9E; B = 8'h70; #100;
A = 8'h9E; B = 8'h71; #100;
A = 8'h9E; B = 8'h72; #100;
A = 8'h9E; B = 8'h73; #100;
A = 8'h9E; B = 8'h74; #100;
A = 8'h9E; B = 8'h75; #100;
A = 8'h9E; B = 8'h76; #100;
A = 8'h9E; B = 8'h77; #100;
A = 8'h9E; B = 8'h78; #100;
A = 8'h9E; B = 8'h79; #100;
A = 8'h9E; B = 8'h7A; #100;
A = 8'h9E; B = 8'h7B; #100;
A = 8'h9E; B = 8'h7C; #100;
A = 8'h9E; B = 8'h7D; #100;
A = 8'h9E; B = 8'h7E; #100;
A = 8'h9E; B = 8'h7F; #100;
A = 8'h9E; B = 8'h80; #100;
A = 8'h9E; B = 8'h81; #100;
A = 8'h9E; B = 8'h82; #100;
A = 8'h9E; B = 8'h83; #100;
A = 8'h9E; B = 8'h84; #100;
A = 8'h9E; B = 8'h85; #100;
A = 8'h9E; B = 8'h86; #100;
A = 8'h9E; B = 8'h87; #100;
A = 8'h9E; B = 8'h88; #100;
A = 8'h9E; B = 8'h89; #100;
A = 8'h9E; B = 8'h8A; #100;
A = 8'h9E; B = 8'h8B; #100;
A = 8'h9E; B = 8'h8C; #100;
A = 8'h9E; B = 8'h8D; #100;
A = 8'h9E; B = 8'h8E; #100;
A = 8'h9E; B = 8'h8F; #100;
A = 8'h9E; B = 8'h90; #100;
A = 8'h9E; B = 8'h91; #100;
A = 8'h9E; B = 8'h92; #100;
A = 8'h9E; B = 8'h93; #100;
A = 8'h9E; B = 8'h94; #100;
A = 8'h9E; B = 8'h95; #100;
A = 8'h9E; B = 8'h96; #100;
A = 8'h9E; B = 8'h97; #100;
A = 8'h9E; B = 8'h98; #100;
A = 8'h9E; B = 8'h99; #100;
A = 8'h9E; B = 8'h9A; #100;
A = 8'h9E; B = 8'h9B; #100;
A = 8'h9E; B = 8'h9C; #100;
A = 8'h9E; B = 8'h9D; #100;
A = 8'h9E; B = 8'h9E; #100;
A = 8'h9E; B = 8'h9F; #100;
A = 8'h9E; B = 8'hA0; #100;
A = 8'h9E; B = 8'hA1; #100;
A = 8'h9E; B = 8'hA2; #100;
A = 8'h9E; B = 8'hA3; #100;
A = 8'h9E; B = 8'hA4; #100;
A = 8'h9E; B = 8'hA5; #100;
A = 8'h9E; B = 8'hA6; #100;
A = 8'h9E; B = 8'hA7; #100;
A = 8'h9E; B = 8'hA8; #100;
A = 8'h9E; B = 8'hA9; #100;
A = 8'h9E; B = 8'hAA; #100;
A = 8'h9E; B = 8'hAB; #100;
A = 8'h9E; B = 8'hAC; #100;
A = 8'h9E; B = 8'hAD; #100;
A = 8'h9E; B = 8'hAE; #100;
A = 8'h9E; B = 8'hAF; #100;
A = 8'h9E; B = 8'hB0; #100;
A = 8'h9E; B = 8'hB1; #100;
A = 8'h9E; B = 8'hB2; #100;
A = 8'h9E; B = 8'hB3; #100;
A = 8'h9E; B = 8'hB4; #100;
A = 8'h9E; B = 8'hB5; #100;
A = 8'h9E; B = 8'hB6; #100;
A = 8'h9E; B = 8'hB7; #100;
A = 8'h9E; B = 8'hB8; #100;
A = 8'h9E; B = 8'hB9; #100;
A = 8'h9E; B = 8'hBA; #100;
A = 8'h9E; B = 8'hBB; #100;
A = 8'h9E; B = 8'hBC; #100;
A = 8'h9E; B = 8'hBD; #100;
A = 8'h9E; B = 8'hBE; #100;
A = 8'h9E; B = 8'hBF; #100;
A = 8'h9E; B = 8'hC0; #100;
A = 8'h9E; B = 8'hC1; #100;
A = 8'h9E; B = 8'hC2; #100;
A = 8'h9E; B = 8'hC3; #100;
A = 8'h9E; B = 8'hC4; #100;
A = 8'h9E; B = 8'hC5; #100;
A = 8'h9E; B = 8'hC6; #100;
A = 8'h9E; B = 8'hC7; #100;
A = 8'h9E; B = 8'hC8; #100;
A = 8'h9E; B = 8'hC9; #100;
A = 8'h9E; B = 8'hCA; #100;
A = 8'h9E; B = 8'hCB; #100;
A = 8'h9E; B = 8'hCC; #100;
A = 8'h9E; B = 8'hCD; #100;
A = 8'h9E; B = 8'hCE; #100;
A = 8'h9E; B = 8'hCF; #100;
A = 8'h9E; B = 8'hD0; #100;
A = 8'h9E; B = 8'hD1; #100;
A = 8'h9E; B = 8'hD2; #100;
A = 8'h9E; B = 8'hD3; #100;
A = 8'h9E; B = 8'hD4; #100;
A = 8'h9E; B = 8'hD5; #100;
A = 8'h9E; B = 8'hD6; #100;
A = 8'h9E; B = 8'hD7; #100;
A = 8'h9E; B = 8'hD8; #100;
A = 8'h9E; B = 8'hD9; #100;
A = 8'h9E; B = 8'hDA; #100;
A = 8'h9E; B = 8'hDB; #100;
A = 8'h9E; B = 8'hDC; #100;
A = 8'h9E; B = 8'hDD; #100;
A = 8'h9E; B = 8'hDE; #100;
A = 8'h9E; B = 8'hDF; #100;
A = 8'h9E; B = 8'hE0; #100;
A = 8'h9E; B = 8'hE1; #100;
A = 8'h9E; B = 8'hE2; #100;
A = 8'h9E; B = 8'hE3; #100;
A = 8'h9E; B = 8'hE4; #100;
A = 8'h9E; B = 8'hE5; #100;
A = 8'h9E; B = 8'hE6; #100;
A = 8'h9E; B = 8'hE7; #100;
A = 8'h9E; B = 8'hE8; #100;
A = 8'h9E; B = 8'hE9; #100;
A = 8'h9E; B = 8'hEA; #100;
A = 8'h9E; B = 8'hEB; #100;
A = 8'h9E; B = 8'hEC; #100;
A = 8'h9E; B = 8'hED; #100;
A = 8'h9E; B = 8'hEE; #100;
A = 8'h9E; B = 8'hEF; #100;
A = 8'h9E; B = 8'hF0; #100;
A = 8'h9E; B = 8'hF1; #100;
A = 8'h9E; B = 8'hF2; #100;
A = 8'h9E; B = 8'hF3; #100;
A = 8'h9E; B = 8'hF4; #100;
A = 8'h9E; B = 8'hF5; #100;
A = 8'h9E; B = 8'hF6; #100;
A = 8'h9E; B = 8'hF7; #100;
A = 8'h9E; B = 8'hF8; #100;
A = 8'h9E; B = 8'hF9; #100;
A = 8'h9E; B = 8'hFA; #100;
A = 8'h9E; B = 8'hFB; #100;
A = 8'h9E; B = 8'hFC; #100;
A = 8'h9E; B = 8'hFD; #100;
A = 8'h9E; B = 8'hFE; #100;
A = 8'h9E; B = 8'hFF; #100;
A = 8'h9F; B = 8'h0; #100;
A = 8'h9F; B = 8'h1; #100;
A = 8'h9F; B = 8'h2; #100;
A = 8'h9F; B = 8'h3; #100;
A = 8'h9F; B = 8'h4; #100;
A = 8'h9F; B = 8'h5; #100;
A = 8'h9F; B = 8'h6; #100;
A = 8'h9F; B = 8'h7; #100;
A = 8'h9F; B = 8'h8; #100;
A = 8'h9F; B = 8'h9; #100;
A = 8'h9F; B = 8'hA; #100;
A = 8'h9F; B = 8'hB; #100;
A = 8'h9F; B = 8'hC; #100;
A = 8'h9F; B = 8'hD; #100;
A = 8'h9F; B = 8'hE; #100;
A = 8'h9F; B = 8'hF; #100;
A = 8'h9F; B = 8'h10; #100;
A = 8'h9F; B = 8'h11; #100;
A = 8'h9F; B = 8'h12; #100;
A = 8'h9F; B = 8'h13; #100;
A = 8'h9F; B = 8'h14; #100;
A = 8'h9F; B = 8'h15; #100;
A = 8'h9F; B = 8'h16; #100;
A = 8'h9F; B = 8'h17; #100;
A = 8'h9F; B = 8'h18; #100;
A = 8'h9F; B = 8'h19; #100;
A = 8'h9F; B = 8'h1A; #100;
A = 8'h9F; B = 8'h1B; #100;
A = 8'h9F; B = 8'h1C; #100;
A = 8'h9F; B = 8'h1D; #100;
A = 8'h9F; B = 8'h1E; #100;
A = 8'h9F; B = 8'h1F; #100;
A = 8'h9F; B = 8'h20; #100;
A = 8'h9F; B = 8'h21; #100;
A = 8'h9F; B = 8'h22; #100;
A = 8'h9F; B = 8'h23; #100;
A = 8'h9F; B = 8'h24; #100;
A = 8'h9F; B = 8'h25; #100;
A = 8'h9F; B = 8'h26; #100;
A = 8'h9F; B = 8'h27; #100;
A = 8'h9F; B = 8'h28; #100;
A = 8'h9F; B = 8'h29; #100;
A = 8'h9F; B = 8'h2A; #100;
A = 8'h9F; B = 8'h2B; #100;
A = 8'h9F; B = 8'h2C; #100;
A = 8'h9F; B = 8'h2D; #100;
A = 8'h9F; B = 8'h2E; #100;
A = 8'h9F; B = 8'h2F; #100;
A = 8'h9F; B = 8'h30; #100;
A = 8'h9F; B = 8'h31; #100;
A = 8'h9F; B = 8'h32; #100;
A = 8'h9F; B = 8'h33; #100;
A = 8'h9F; B = 8'h34; #100;
A = 8'h9F; B = 8'h35; #100;
A = 8'h9F; B = 8'h36; #100;
A = 8'h9F; B = 8'h37; #100;
A = 8'h9F; B = 8'h38; #100;
A = 8'h9F; B = 8'h39; #100;
A = 8'h9F; B = 8'h3A; #100;
A = 8'h9F; B = 8'h3B; #100;
A = 8'h9F; B = 8'h3C; #100;
A = 8'h9F; B = 8'h3D; #100;
A = 8'h9F; B = 8'h3E; #100;
A = 8'h9F; B = 8'h3F; #100;
A = 8'h9F; B = 8'h40; #100;
A = 8'h9F; B = 8'h41; #100;
A = 8'h9F; B = 8'h42; #100;
A = 8'h9F; B = 8'h43; #100;
A = 8'h9F; B = 8'h44; #100;
A = 8'h9F; B = 8'h45; #100;
A = 8'h9F; B = 8'h46; #100;
A = 8'h9F; B = 8'h47; #100;
A = 8'h9F; B = 8'h48; #100;
A = 8'h9F; B = 8'h49; #100;
A = 8'h9F; B = 8'h4A; #100;
A = 8'h9F; B = 8'h4B; #100;
A = 8'h9F; B = 8'h4C; #100;
A = 8'h9F; B = 8'h4D; #100;
A = 8'h9F; B = 8'h4E; #100;
A = 8'h9F; B = 8'h4F; #100;
A = 8'h9F; B = 8'h50; #100;
A = 8'h9F; B = 8'h51; #100;
A = 8'h9F; B = 8'h52; #100;
A = 8'h9F; B = 8'h53; #100;
A = 8'h9F; B = 8'h54; #100;
A = 8'h9F; B = 8'h55; #100;
A = 8'h9F; B = 8'h56; #100;
A = 8'h9F; B = 8'h57; #100;
A = 8'h9F; B = 8'h58; #100;
A = 8'h9F; B = 8'h59; #100;
A = 8'h9F; B = 8'h5A; #100;
A = 8'h9F; B = 8'h5B; #100;
A = 8'h9F; B = 8'h5C; #100;
A = 8'h9F; B = 8'h5D; #100;
A = 8'h9F; B = 8'h5E; #100;
A = 8'h9F; B = 8'h5F; #100;
A = 8'h9F; B = 8'h60; #100;
A = 8'h9F; B = 8'h61; #100;
A = 8'h9F; B = 8'h62; #100;
A = 8'h9F; B = 8'h63; #100;
A = 8'h9F; B = 8'h64; #100;
A = 8'h9F; B = 8'h65; #100;
A = 8'h9F; B = 8'h66; #100;
A = 8'h9F; B = 8'h67; #100;
A = 8'h9F; B = 8'h68; #100;
A = 8'h9F; B = 8'h69; #100;
A = 8'h9F; B = 8'h6A; #100;
A = 8'h9F; B = 8'h6B; #100;
A = 8'h9F; B = 8'h6C; #100;
A = 8'h9F; B = 8'h6D; #100;
A = 8'h9F; B = 8'h6E; #100;
A = 8'h9F; B = 8'h6F; #100;
A = 8'h9F; B = 8'h70; #100;
A = 8'h9F; B = 8'h71; #100;
A = 8'h9F; B = 8'h72; #100;
A = 8'h9F; B = 8'h73; #100;
A = 8'h9F; B = 8'h74; #100;
A = 8'h9F; B = 8'h75; #100;
A = 8'h9F; B = 8'h76; #100;
A = 8'h9F; B = 8'h77; #100;
A = 8'h9F; B = 8'h78; #100;
A = 8'h9F; B = 8'h79; #100;
A = 8'h9F; B = 8'h7A; #100;
A = 8'h9F; B = 8'h7B; #100;
A = 8'h9F; B = 8'h7C; #100;
A = 8'h9F; B = 8'h7D; #100;
A = 8'h9F; B = 8'h7E; #100;
A = 8'h9F; B = 8'h7F; #100;
A = 8'h9F; B = 8'h80; #100;
A = 8'h9F; B = 8'h81; #100;
A = 8'h9F; B = 8'h82; #100;
A = 8'h9F; B = 8'h83; #100;
A = 8'h9F; B = 8'h84; #100;
A = 8'h9F; B = 8'h85; #100;
A = 8'h9F; B = 8'h86; #100;
A = 8'h9F; B = 8'h87; #100;
A = 8'h9F; B = 8'h88; #100;
A = 8'h9F; B = 8'h89; #100;
A = 8'h9F; B = 8'h8A; #100;
A = 8'h9F; B = 8'h8B; #100;
A = 8'h9F; B = 8'h8C; #100;
A = 8'h9F; B = 8'h8D; #100;
A = 8'h9F; B = 8'h8E; #100;
A = 8'h9F; B = 8'h8F; #100;
A = 8'h9F; B = 8'h90; #100;
A = 8'h9F; B = 8'h91; #100;
A = 8'h9F; B = 8'h92; #100;
A = 8'h9F; B = 8'h93; #100;
A = 8'h9F; B = 8'h94; #100;
A = 8'h9F; B = 8'h95; #100;
A = 8'h9F; B = 8'h96; #100;
A = 8'h9F; B = 8'h97; #100;
A = 8'h9F; B = 8'h98; #100;
A = 8'h9F; B = 8'h99; #100;
A = 8'h9F; B = 8'h9A; #100;
A = 8'h9F; B = 8'h9B; #100;
A = 8'h9F; B = 8'h9C; #100;
A = 8'h9F; B = 8'h9D; #100;
A = 8'h9F; B = 8'h9E; #100;
A = 8'h9F; B = 8'h9F; #100;
A = 8'h9F; B = 8'hA0; #100;
A = 8'h9F; B = 8'hA1; #100;
A = 8'h9F; B = 8'hA2; #100;
A = 8'h9F; B = 8'hA3; #100;
A = 8'h9F; B = 8'hA4; #100;
A = 8'h9F; B = 8'hA5; #100;
A = 8'h9F; B = 8'hA6; #100;
A = 8'h9F; B = 8'hA7; #100;
A = 8'h9F; B = 8'hA8; #100;
A = 8'h9F; B = 8'hA9; #100;
A = 8'h9F; B = 8'hAA; #100;
A = 8'h9F; B = 8'hAB; #100;
A = 8'h9F; B = 8'hAC; #100;
A = 8'h9F; B = 8'hAD; #100;
A = 8'h9F; B = 8'hAE; #100;
A = 8'h9F; B = 8'hAF; #100;
A = 8'h9F; B = 8'hB0; #100;
A = 8'h9F; B = 8'hB1; #100;
A = 8'h9F; B = 8'hB2; #100;
A = 8'h9F; B = 8'hB3; #100;
A = 8'h9F; B = 8'hB4; #100;
A = 8'h9F; B = 8'hB5; #100;
A = 8'h9F; B = 8'hB6; #100;
A = 8'h9F; B = 8'hB7; #100;
A = 8'h9F; B = 8'hB8; #100;
A = 8'h9F; B = 8'hB9; #100;
A = 8'h9F; B = 8'hBA; #100;
A = 8'h9F; B = 8'hBB; #100;
A = 8'h9F; B = 8'hBC; #100;
A = 8'h9F; B = 8'hBD; #100;
A = 8'h9F; B = 8'hBE; #100;
A = 8'h9F; B = 8'hBF; #100;
A = 8'h9F; B = 8'hC0; #100;
A = 8'h9F; B = 8'hC1; #100;
A = 8'h9F; B = 8'hC2; #100;
A = 8'h9F; B = 8'hC3; #100;
A = 8'h9F; B = 8'hC4; #100;
A = 8'h9F; B = 8'hC5; #100;
A = 8'h9F; B = 8'hC6; #100;
A = 8'h9F; B = 8'hC7; #100;
A = 8'h9F; B = 8'hC8; #100;
A = 8'h9F; B = 8'hC9; #100;
A = 8'h9F; B = 8'hCA; #100;
A = 8'h9F; B = 8'hCB; #100;
A = 8'h9F; B = 8'hCC; #100;
A = 8'h9F; B = 8'hCD; #100;
A = 8'h9F; B = 8'hCE; #100;
A = 8'h9F; B = 8'hCF; #100;
A = 8'h9F; B = 8'hD0; #100;
A = 8'h9F; B = 8'hD1; #100;
A = 8'h9F; B = 8'hD2; #100;
A = 8'h9F; B = 8'hD3; #100;
A = 8'h9F; B = 8'hD4; #100;
A = 8'h9F; B = 8'hD5; #100;
A = 8'h9F; B = 8'hD6; #100;
A = 8'h9F; B = 8'hD7; #100;
A = 8'h9F; B = 8'hD8; #100;
A = 8'h9F; B = 8'hD9; #100;
A = 8'h9F; B = 8'hDA; #100;
A = 8'h9F; B = 8'hDB; #100;
A = 8'h9F; B = 8'hDC; #100;
A = 8'h9F; B = 8'hDD; #100;
A = 8'h9F; B = 8'hDE; #100;
A = 8'h9F; B = 8'hDF; #100;
A = 8'h9F; B = 8'hE0; #100;
A = 8'h9F; B = 8'hE1; #100;
A = 8'h9F; B = 8'hE2; #100;
A = 8'h9F; B = 8'hE3; #100;
A = 8'h9F; B = 8'hE4; #100;
A = 8'h9F; B = 8'hE5; #100;
A = 8'h9F; B = 8'hE6; #100;
A = 8'h9F; B = 8'hE7; #100;
A = 8'h9F; B = 8'hE8; #100;
A = 8'h9F; B = 8'hE9; #100;
A = 8'h9F; B = 8'hEA; #100;
A = 8'h9F; B = 8'hEB; #100;
A = 8'h9F; B = 8'hEC; #100;
A = 8'h9F; B = 8'hED; #100;
A = 8'h9F; B = 8'hEE; #100;
A = 8'h9F; B = 8'hEF; #100;
A = 8'h9F; B = 8'hF0; #100;
A = 8'h9F; B = 8'hF1; #100;
A = 8'h9F; B = 8'hF2; #100;
A = 8'h9F; B = 8'hF3; #100;
A = 8'h9F; B = 8'hF4; #100;
A = 8'h9F; B = 8'hF5; #100;
A = 8'h9F; B = 8'hF6; #100;
A = 8'h9F; B = 8'hF7; #100;
A = 8'h9F; B = 8'hF8; #100;
A = 8'h9F; B = 8'hF9; #100;
A = 8'h9F; B = 8'hFA; #100;
A = 8'h9F; B = 8'hFB; #100;
A = 8'h9F; B = 8'hFC; #100;
A = 8'h9F; B = 8'hFD; #100;
A = 8'h9F; B = 8'hFE; #100;
A = 8'h9F; B = 8'hFF; #100;
A = 8'hA0; B = 8'h0; #100;
A = 8'hA0; B = 8'h1; #100;
A = 8'hA0; B = 8'h2; #100;
A = 8'hA0; B = 8'h3; #100;
A = 8'hA0; B = 8'h4; #100;
A = 8'hA0; B = 8'h5; #100;
A = 8'hA0; B = 8'h6; #100;
A = 8'hA0; B = 8'h7; #100;
A = 8'hA0; B = 8'h8; #100;
A = 8'hA0; B = 8'h9; #100;
A = 8'hA0; B = 8'hA; #100;
A = 8'hA0; B = 8'hB; #100;
A = 8'hA0; B = 8'hC; #100;
A = 8'hA0; B = 8'hD; #100;
A = 8'hA0; B = 8'hE; #100;
A = 8'hA0; B = 8'hF; #100;
A = 8'hA0; B = 8'h10; #100;
A = 8'hA0; B = 8'h11; #100;
A = 8'hA0; B = 8'h12; #100;
A = 8'hA0; B = 8'h13; #100;
A = 8'hA0; B = 8'h14; #100;
A = 8'hA0; B = 8'h15; #100;
A = 8'hA0; B = 8'h16; #100;
A = 8'hA0; B = 8'h17; #100;
A = 8'hA0; B = 8'h18; #100;
A = 8'hA0; B = 8'h19; #100;
A = 8'hA0; B = 8'h1A; #100;
A = 8'hA0; B = 8'h1B; #100;
A = 8'hA0; B = 8'h1C; #100;
A = 8'hA0; B = 8'h1D; #100;
A = 8'hA0; B = 8'h1E; #100;
A = 8'hA0; B = 8'h1F; #100;
A = 8'hA0; B = 8'h20; #100;
A = 8'hA0; B = 8'h21; #100;
A = 8'hA0; B = 8'h22; #100;
A = 8'hA0; B = 8'h23; #100;
A = 8'hA0; B = 8'h24; #100;
A = 8'hA0; B = 8'h25; #100;
A = 8'hA0; B = 8'h26; #100;
A = 8'hA0; B = 8'h27; #100;
A = 8'hA0; B = 8'h28; #100;
A = 8'hA0; B = 8'h29; #100;
A = 8'hA0; B = 8'h2A; #100;
A = 8'hA0; B = 8'h2B; #100;
A = 8'hA0; B = 8'h2C; #100;
A = 8'hA0; B = 8'h2D; #100;
A = 8'hA0; B = 8'h2E; #100;
A = 8'hA0; B = 8'h2F; #100;
A = 8'hA0; B = 8'h30; #100;
A = 8'hA0; B = 8'h31; #100;
A = 8'hA0; B = 8'h32; #100;
A = 8'hA0; B = 8'h33; #100;
A = 8'hA0; B = 8'h34; #100;
A = 8'hA0; B = 8'h35; #100;
A = 8'hA0; B = 8'h36; #100;
A = 8'hA0; B = 8'h37; #100;
A = 8'hA0; B = 8'h38; #100;
A = 8'hA0; B = 8'h39; #100;
A = 8'hA0; B = 8'h3A; #100;
A = 8'hA0; B = 8'h3B; #100;
A = 8'hA0; B = 8'h3C; #100;
A = 8'hA0; B = 8'h3D; #100;
A = 8'hA0; B = 8'h3E; #100;
A = 8'hA0; B = 8'h3F; #100;
A = 8'hA0; B = 8'h40; #100;
A = 8'hA0; B = 8'h41; #100;
A = 8'hA0; B = 8'h42; #100;
A = 8'hA0; B = 8'h43; #100;
A = 8'hA0; B = 8'h44; #100;
A = 8'hA0; B = 8'h45; #100;
A = 8'hA0; B = 8'h46; #100;
A = 8'hA0; B = 8'h47; #100;
A = 8'hA0; B = 8'h48; #100;
A = 8'hA0; B = 8'h49; #100;
A = 8'hA0; B = 8'h4A; #100;
A = 8'hA0; B = 8'h4B; #100;
A = 8'hA0; B = 8'h4C; #100;
A = 8'hA0; B = 8'h4D; #100;
A = 8'hA0; B = 8'h4E; #100;
A = 8'hA0; B = 8'h4F; #100;
A = 8'hA0; B = 8'h50; #100;
A = 8'hA0; B = 8'h51; #100;
A = 8'hA0; B = 8'h52; #100;
A = 8'hA0; B = 8'h53; #100;
A = 8'hA0; B = 8'h54; #100;
A = 8'hA0; B = 8'h55; #100;
A = 8'hA0; B = 8'h56; #100;
A = 8'hA0; B = 8'h57; #100;
A = 8'hA0; B = 8'h58; #100;
A = 8'hA0; B = 8'h59; #100;
A = 8'hA0; B = 8'h5A; #100;
A = 8'hA0; B = 8'h5B; #100;
A = 8'hA0; B = 8'h5C; #100;
A = 8'hA0; B = 8'h5D; #100;
A = 8'hA0; B = 8'h5E; #100;
A = 8'hA0; B = 8'h5F; #100;
A = 8'hA0; B = 8'h60; #100;
A = 8'hA0; B = 8'h61; #100;
A = 8'hA0; B = 8'h62; #100;
A = 8'hA0; B = 8'h63; #100;
A = 8'hA0; B = 8'h64; #100;
A = 8'hA0; B = 8'h65; #100;
A = 8'hA0; B = 8'h66; #100;
A = 8'hA0; B = 8'h67; #100;
A = 8'hA0; B = 8'h68; #100;
A = 8'hA0; B = 8'h69; #100;
A = 8'hA0; B = 8'h6A; #100;
A = 8'hA0; B = 8'h6B; #100;
A = 8'hA0; B = 8'h6C; #100;
A = 8'hA0; B = 8'h6D; #100;
A = 8'hA0; B = 8'h6E; #100;
A = 8'hA0; B = 8'h6F; #100;
A = 8'hA0; B = 8'h70; #100;
A = 8'hA0; B = 8'h71; #100;
A = 8'hA0; B = 8'h72; #100;
A = 8'hA0; B = 8'h73; #100;
A = 8'hA0; B = 8'h74; #100;
A = 8'hA0; B = 8'h75; #100;
A = 8'hA0; B = 8'h76; #100;
A = 8'hA0; B = 8'h77; #100;
A = 8'hA0; B = 8'h78; #100;
A = 8'hA0; B = 8'h79; #100;
A = 8'hA0; B = 8'h7A; #100;
A = 8'hA0; B = 8'h7B; #100;
A = 8'hA0; B = 8'h7C; #100;
A = 8'hA0; B = 8'h7D; #100;
A = 8'hA0; B = 8'h7E; #100;
A = 8'hA0; B = 8'h7F; #100;
A = 8'hA0; B = 8'h80; #100;
A = 8'hA0; B = 8'h81; #100;
A = 8'hA0; B = 8'h82; #100;
A = 8'hA0; B = 8'h83; #100;
A = 8'hA0; B = 8'h84; #100;
A = 8'hA0; B = 8'h85; #100;
A = 8'hA0; B = 8'h86; #100;
A = 8'hA0; B = 8'h87; #100;
A = 8'hA0; B = 8'h88; #100;
A = 8'hA0; B = 8'h89; #100;
A = 8'hA0; B = 8'h8A; #100;
A = 8'hA0; B = 8'h8B; #100;
A = 8'hA0; B = 8'h8C; #100;
A = 8'hA0; B = 8'h8D; #100;
A = 8'hA0; B = 8'h8E; #100;
A = 8'hA0; B = 8'h8F; #100;
A = 8'hA0; B = 8'h90; #100;
A = 8'hA0; B = 8'h91; #100;
A = 8'hA0; B = 8'h92; #100;
A = 8'hA0; B = 8'h93; #100;
A = 8'hA0; B = 8'h94; #100;
A = 8'hA0; B = 8'h95; #100;
A = 8'hA0; B = 8'h96; #100;
A = 8'hA0; B = 8'h97; #100;
A = 8'hA0; B = 8'h98; #100;
A = 8'hA0; B = 8'h99; #100;
A = 8'hA0; B = 8'h9A; #100;
A = 8'hA0; B = 8'h9B; #100;
A = 8'hA0; B = 8'h9C; #100;
A = 8'hA0; B = 8'h9D; #100;
A = 8'hA0; B = 8'h9E; #100;
A = 8'hA0; B = 8'h9F; #100;
A = 8'hA0; B = 8'hA0; #100;
A = 8'hA0; B = 8'hA1; #100;
A = 8'hA0; B = 8'hA2; #100;
A = 8'hA0; B = 8'hA3; #100;
A = 8'hA0; B = 8'hA4; #100;
A = 8'hA0; B = 8'hA5; #100;
A = 8'hA0; B = 8'hA6; #100;
A = 8'hA0; B = 8'hA7; #100;
A = 8'hA0; B = 8'hA8; #100;
A = 8'hA0; B = 8'hA9; #100;
A = 8'hA0; B = 8'hAA; #100;
A = 8'hA0; B = 8'hAB; #100;
A = 8'hA0; B = 8'hAC; #100;
A = 8'hA0; B = 8'hAD; #100;
A = 8'hA0; B = 8'hAE; #100;
A = 8'hA0; B = 8'hAF; #100;
A = 8'hA0; B = 8'hB0; #100;
A = 8'hA0; B = 8'hB1; #100;
A = 8'hA0; B = 8'hB2; #100;
A = 8'hA0; B = 8'hB3; #100;
A = 8'hA0; B = 8'hB4; #100;
A = 8'hA0; B = 8'hB5; #100;
A = 8'hA0; B = 8'hB6; #100;
A = 8'hA0; B = 8'hB7; #100;
A = 8'hA0; B = 8'hB8; #100;
A = 8'hA0; B = 8'hB9; #100;
A = 8'hA0; B = 8'hBA; #100;
A = 8'hA0; B = 8'hBB; #100;
A = 8'hA0; B = 8'hBC; #100;
A = 8'hA0; B = 8'hBD; #100;
A = 8'hA0; B = 8'hBE; #100;
A = 8'hA0; B = 8'hBF; #100;
A = 8'hA0; B = 8'hC0; #100;
A = 8'hA0; B = 8'hC1; #100;
A = 8'hA0; B = 8'hC2; #100;
A = 8'hA0; B = 8'hC3; #100;
A = 8'hA0; B = 8'hC4; #100;
A = 8'hA0; B = 8'hC5; #100;
A = 8'hA0; B = 8'hC6; #100;
A = 8'hA0; B = 8'hC7; #100;
A = 8'hA0; B = 8'hC8; #100;
A = 8'hA0; B = 8'hC9; #100;
A = 8'hA0; B = 8'hCA; #100;
A = 8'hA0; B = 8'hCB; #100;
A = 8'hA0; B = 8'hCC; #100;
A = 8'hA0; B = 8'hCD; #100;
A = 8'hA0; B = 8'hCE; #100;
A = 8'hA0; B = 8'hCF; #100;
A = 8'hA0; B = 8'hD0; #100;
A = 8'hA0; B = 8'hD1; #100;
A = 8'hA0; B = 8'hD2; #100;
A = 8'hA0; B = 8'hD3; #100;
A = 8'hA0; B = 8'hD4; #100;
A = 8'hA0; B = 8'hD5; #100;
A = 8'hA0; B = 8'hD6; #100;
A = 8'hA0; B = 8'hD7; #100;
A = 8'hA0; B = 8'hD8; #100;
A = 8'hA0; B = 8'hD9; #100;
A = 8'hA0; B = 8'hDA; #100;
A = 8'hA0; B = 8'hDB; #100;
A = 8'hA0; B = 8'hDC; #100;
A = 8'hA0; B = 8'hDD; #100;
A = 8'hA0; B = 8'hDE; #100;
A = 8'hA0; B = 8'hDF; #100;
A = 8'hA0; B = 8'hE0; #100;
A = 8'hA0; B = 8'hE1; #100;
A = 8'hA0; B = 8'hE2; #100;
A = 8'hA0; B = 8'hE3; #100;
A = 8'hA0; B = 8'hE4; #100;
A = 8'hA0; B = 8'hE5; #100;
A = 8'hA0; B = 8'hE6; #100;
A = 8'hA0; B = 8'hE7; #100;
A = 8'hA0; B = 8'hE8; #100;
A = 8'hA0; B = 8'hE9; #100;
A = 8'hA0; B = 8'hEA; #100;
A = 8'hA0; B = 8'hEB; #100;
A = 8'hA0; B = 8'hEC; #100;
A = 8'hA0; B = 8'hED; #100;
A = 8'hA0; B = 8'hEE; #100;
A = 8'hA0; B = 8'hEF; #100;
A = 8'hA0; B = 8'hF0; #100;
A = 8'hA0; B = 8'hF1; #100;
A = 8'hA0; B = 8'hF2; #100;
A = 8'hA0; B = 8'hF3; #100;
A = 8'hA0; B = 8'hF4; #100;
A = 8'hA0; B = 8'hF5; #100;
A = 8'hA0; B = 8'hF6; #100;
A = 8'hA0; B = 8'hF7; #100;
A = 8'hA0; B = 8'hF8; #100;
A = 8'hA0; B = 8'hF9; #100;
A = 8'hA0; B = 8'hFA; #100;
A = 8'hA0; B = 8'hFB; #100;
A = 8'hA0; B = 8'hFC; #100;
A = 8'hA0; B = 8'hFD; #100;
A = 8'hA0; B = 8'hFE; #100;
A = 8'hA0; B = 8'hFF; #100;
A = 8'hA1; B = 8'h0; #100;
A = 8'hA1; B = 8'h1; #100;
A = 8'hA1; B = 8'h2; #100;
A = 8'hA1; B = 8'h3; #100;
A = 8'hA1; B = 8'h4; #100;
A = 8'hA1; B = 8'h5; #100;
A = 8'hA1; B = 8'h6; #100;
A = 8'hA1; B = 8'h7; #100;
A = 8'hA1; B = 8'h8; #100;
A = 8'hA1; B = 8'h9; #100;
A = 8'hA1; B = 8'hA; #100;
A = 8'hA1; B = 8'hB; #100;
A = 8'hA1; B = 8'hC; #100;
A = 8'hA1; B = 8'hD; #100;
A = 8'hA1; B = 8'hE; #100;
A = 8'hA1; B = 8'hF; #100;
A = 8'hA1; B = 8'h10; #100;
A = 8'hA1; B = 8'h11; #100;
A = 8'hA1; B = 8'h12; #100;
A = 8'hA1; B = 8'h13; #100;
A = 8'hA1; B = 8'h14; #100;
A = 8'hA1; B = 8'h15; #100;
A = 8'hA1; B = 8'h16; #100;
A = 8'hA1; B = 8'h17; #100;
A = 8'hA1; B = 8'h18; #100;
A = 8'hA1; B = 8'h19; #100;
A = 8'hA1; B = 8'h1A; #100;
A = 8'hA1; B = 8'h1B; #100;
A = 8'hA1; B = 8'h1C; #100;
A = 8'hA1; B = 8'h1D; #100;
A = 8'hA1; B = 8'h1E; #100;
A = 8'hA1; B = 8'h1F; #100;
A = 8'hA1; B = 8'h20; #100;
A = 8'hA1; B = 8'h21; #100;
A = 8'hA1; B = 8'h22; #100;
A = 8'hA1; B = 8'h23; #100;
A = 8'hA1; B = 8'h24; #100;
A = 8'hA1; B = 8'h25; #100;
A = 8'hA1; B = 8'h26; #100;
A = 8'hA1; B = 8'h27; #100;
A = 8'hA1; B = 8'h28; #100;
A = 8'hA1; B = 8'h29; #100;
A = 8'hA1; B = 8'h2A; #100;
A = 8'hA1; B = 8'h2B; #100;
A = 8'hA1; B = 8'h2C; #100;
A = 8'hA1; B = 8'h2D; #100;
A = 8'hA1; B = 8'h2E; #100;
A = 8'hA1; B = 8'h2F; #100;
A = 8'hA1; B = 8'h30; #100;
A = 8'hA1; B = 8'h31; #100;
A = 8'hA1; B = 8'h32; #100;
A = 8'hA1; B = 8'h33; #100;
A = 8'hA1; B = 8'h34; #100;
A = 8'hA1; B = 8'h35; #100;
A = 8'hA1; B = 8'h36; #100;
A = 8'hA1; B = 8'h37; #100;
A = 8'hA1; B = 8'h38; #100;
A = 8'hA1; B = 8'h39; #100;
A = 8'hA1; B = 8'h3A; #100;
A = 8'hA1; B = 8'h3B; #100;
A = 8'hA1; B = 8'h3C; #100;
A = 8'hA1; B = 8'h3D; #100;
A = 8'hA1; B = 8'h3E; #100;
A = 8'hA1; B = 8'h3F; #100;
A = 8'hA1; B = 8'h40; #100;
A = 8'hA1; B = 8'h41; #100;
A = 8'hA1; B = 8'h42; #100;
A = 8'hA1; B = 8'h43; #100;
A = 8'hA1; B = 8'h44; #100;
A = 8'hA1; B = 8'h45; #100;
A = 8'hA1; B = 8'h46; #100;
A = 8'hA1; B = 8'h47; #100;
A = 8'hA1; B = 8'h48; #100;
A = 8'hA1; B = 8'h49; #100;
A = 8'hA1; B = 8'h4A; #100;
A = 8'hA1; B = 8'h4B; #100;
A = 8'hA1; B = 8'h4C; #100;
A = 8'hA1; B = 8'h4D; #100;
A = 8'hA1; B = 8'h4E; #100;
A = 8'hA1; B = 8'h4F; #100;
A = 8'hA1; B = 8'h50; #100;
A = 8'hA1; B = 8'h51; #100;
A = 8'hA1; B = 8'h52; #100;
A = 8'hA1; B = 8'h53; #100;
A = 8'hA1; B = 8'h54; #100;
A = 8'hA1; B = 8'h55; #100;
A = 8'hA1; B = 8'h56; #100;
A = 8'hA1; B = 8'h57; #100;
A = 8'hA1; B = 8'h58; #100;
A = 8'hA1; B = 8'h59; #100;
A = 8'hA1; B = 8'h5A; #100;
A = 8'hA1; B = 8'h5B; #100;
A = 8'hA1; B = 8'h5C; #100;
A = 8'hA1; B = 8'h5D; #100;
A = 8'hA1; B = 8'h5E; #100;
A = 8'hA1; B = 8'h5F; #100;
A = 8'hA1; B = 8'h60; #100;
A = 8'hA1; B = 8'h61; #100;
A = 8'hA1; B = 8'h62; #100;
A = 8'hA1; B = 8'h63; #100;
A = 8'hA1; B = 8'h64; #100;
A = 8'hA1; B = 8'h65; #100;
A = 8'hA1; B = 8'h66; #100;
A = 8'hA1; B = 8'h67; #100;
A = 8'hA1; B = 8'h68; #100;
A = 8'hA1; B = 8'h69; #100;
A = 8'hA1; B = 8'h6A; #100;
A = 8'hA1; B = 8'h6B; #100;
A = 8'hA1; B = 8'h6C; #100;
A = 8'hA1; B = 8'h6D; #100;
A = 8'hA1; B = 8'h6E; #100;
A = 8'hA1; B = 8'h6F; #100;
A = 8'hA1; B = 8'h70; #100;
A = 8'hA1; B = 8'h71; #100;
A = 8'hA1; B = 8'h72; #100;
A = 8'hA1; B = 8'h73; #100;
A = 8'hA1; B = 8'h74; #100;
A = 8'hA1; B = 8'h75; #100;
A = 8'hA1; B = 8'h76; #100;
A = 8'hA1; B = 8'h77; #100;
A = 8'hA1; B = 8'h78; #100;
A = 8'hA1; B = 8'h79; #100;
A = 8'hA1; B = 8'h7A; #100;
A = 8'hA1; B = 8'h7B; #100;
A = 8'hA1; B = 8'h7C; #100;
A = 8'hA1; B = 8'h7D; #100;
A = 8'hA1; B = 8'h7E; #100;
A = 8'hA1; B = 8'h7F; #100;
A = 8'hA1; B = 8'h80; #100;
A = 8'hA1; B = 8'h81; #100;
A = 8'hA1; B = 8'h82; #100;
A = 8'hA1; B = 8'h83; #100;
A = 8'hA1; B = 8'h84; #100;
A = 8'hA1; B = 8'h85; #100;
A = 8'hA1; B = 8'h86; #100;
A = 8'hA1; B = 8'h87; #100;
A = 8'hA1; B = 8'h88; #100;
A = 8'hA1; B = 8'h89; #100;
A = 8'hA1; B = 8'h8A; #100;
A = 8'hA1; B = 8'h8B; #100;
A = 8'hA1; B = 8'h8C; #100;
A = 8'hA1; B = 8'h8D; #100;
A = 8'hA1; B = 8'h8E; #100;
A = 8'hA1; B = 8'h8F; #100;
A = 8'hA1; B = 8'h90; #100;
A = 8'hA1; B = 8'h91; #100;
A = 8'hA1; B = 8'h92; #100;
A = 8'hA1; B = 8'h93; #100;
A = 8'hA1; B = 8'h94; #100;
A = 8'hA1; B = 8'h95; #100;
A = 8'hA1; B = 8'h96; #100;
A = 8'hA1; B = 8'h97; #100;
A = 8'hA1; B = 8'h98; #100;
A = 8'hA1; B = 8'h99; #100;
A = 8'hA1; B = 8'h9A; #100;
A = 8'hA1; B = 8'h9B; #100;
A = 8'hA1; B = 8'h9C; #100;
A = 8'hA1; B = 8'h9D; #100;
A = 8'hA1; B = 8'h9E; #100;
A = 8'hA1; B = 8'h9F; #100;
A = 8'hA1; B = 8'hA0; #100;
A = 8'hA1; B = 8'hA1; #100;
A = 8'hA1; B = 8'hA2; #100;
A = 8'hA1; B = 8'hA3; #100;
A = 8'hA1; B = 8'hA4; #100;
A = 8'hA1; B = 8'hA5; #100;
A = 8'hA1; B = 8'hA6; #100;
A = 8'hA1; B = 8'hA7; #100;
A = 8'hA1; B = 8'hA8; #100;
A = 8'hA1; B = 8'hA9; #100;
A = 8'hA1; B = 8'hAA; #100;
A = 8'hA1; B = 8'hAB; #100;
A = 8'hA1; B = 8'hAC; #100;
A = 8'hA1; B = 8'hAD; #100;
A = 8'hA1; B = 8'hAE; #100;
A = 8'hA1; B = 8'hAF; #100;
A = 8'hA1; B = 8'hB0; #100;
A = 8'hA1; B = 8'hB1; #100;
A = 8'hA1; B = 8'hB2; #100;
A = 8'hA1; B = 8'hB3; #100;
A = 8'hA1; B = 8'hB4; #100;
A = 8'hA1; B = 8'hB5; #100;
A = 8'hA1; B = 8'hB6; #100;
A = 8'hA1; B = 8'hB7; #100;
A = 8'hA1; B = 8'hB8; #100;
A = 8'hA1; B = 8'hB9; #100;
A = 8'hA1; B = 8'hBA; #100;
A = 8'hA1; B = 8'hBB; #100;
A = 8'hA1; B = 8'hBC; #100;
A = 8'hA1; B = 8'hBD; #100;
A = 8'hA1; B = 8'hBE; #100;
A = 8'hA1; B = 8'hBF; #100;
A = 8'hA1; B = 8'hC0; #100;
A = 8'hA1; B = 8'hC1; #100;
A = 8'hA1; B = 8'hC2; #100;
A = 8'hA1; B = 8'hC3; #100;
A = 8'hA1; B = 8'hC4; #100;
A = 8'hA1; B = 8'hC5; #100;
A = 8'hA1; B = 8'hC6; #100;
A = 8'hA1; B = 8'hC7; #100;
A = 8'hA1; B = 8'hC8; #100;
A = 8'hA1; B = 8'hC9; #100;
A = 8'hA1; B = 8'hCA; #100;
A = 8'hA1; B = 8'hCB; #100;
A = 8'hA1; B = 8'hCC; #100;
A = 8'hA1; B = 8'hCD; #100;
A = 8'hA1; B = 8'hCE; #100;
A = 8'hA1; B = 8'hCF; #100;
A = 8'hA1; B = 8'hD0; #100;
A = 8'hA1; B = 8'hD1; #100;
A = 8'hA1; B = 8'hD2; #100;
A = 8'hA1; B = 8'hD3; #100;
A = 8'hA1; B = 8'hD4; #100;
A = 8'hA1; B = 8'hD5; #100;
A = 8'hA1; B = 8'hD6; #100;
A = 8'hA1; B = 8'hD7; #100;
A = 8'hA1; B = 8'hD8; #100;
A = 8'hA1; B = 8'hD9; #100;
A = 8'hA1; B = 8'hDA; #100;
A = 8'hA1; B = 8'hDB; #100;
A = 8'hA1; B = 8'hDC; #100;
A = 8'hA1; B = 8'hDD; #100;
A = 8'hA1; B = 8'hDE; #100;
A = 8'hA1; B = 8'hDF; #100;
A = 8'hA1; B = 8'hE0; #100;
A = 8'hA1; B = 8'hE1; #100;
A = 8'hA1; B = 8'hE2; #100;
A = 8'hA1; B = 8'hE3; #100;
A = 8'hA1; B = 8'hE4; #100;
A = 8'hA1; B = 8'hE5; #100;
A = 8'hA1; B = 8'hE6; #100;
A = 8'hA1; B = 8'hE7; #100;
A = 8'hA1; B = 8'hE8; #100;
A = 8'hA1; B = 8'hE9; #100;
A = 8'hA1; B = 8'hEA; #100;
A = 8'hA1; B = 8'hEB; #100;
A = 8'hA1; B = 8'hEC; #100;
A = 8'hA1; B = 8'hED; #100;
A = 8'hA1; B = 8'hEE; #100;
A = 8'hA1; B = 8'hEF; #100;
A = 8'hA1; B = 8'hF0; #100;
A = 8'hA1; B = 8'hF1; #100;
A = 8'hA1; B = 8'hF2; #100;
A = 8'hA1; B = 8'hF3; #100;
A = 8'hA1; B = 8'hF4; #100;
A = 8'hA1; B = 8'hF5; #100;
A = 8'hA1; B = 8'hF6; #100;
A = 8'hA1; B = 8'hF7; #100;
A = 8'hA1; B = 8'hF8; #100;
A = 8'hA1; B = 8'hF9; #100;
A = 8'hA1; B = 8'hFA; #100;
A = 8'hA1; B = 8'hFB; #100;
A = 8'hA1; B = 8'hFC; #100;
A = 8'hA1; B = 8'hFD; #100;
A = 8'hA1; B = 8'hFE; #100;
A = 8'hA1; B = 8'hFF; #100;
A = 8'hA2; B = 8'h0; #100;
A = 8'hA2; B = 8'h1; #100;
A = 8'hA2; B = 8'h2; #100;
A = 8'hA2; B = 8'h3; #100;
A = 8'hA2; B = 8'h4; #100;
A = 8'hA2; B = 8'h5; #100;
A = 8'hA2; B = 8'h6; #100;
A = 8'hA2; B = 8'h7; #100;
A = 8'hA2; B = 8'h8; #100;
A = 8'hA2; B = 8'h9; #100;
A = 8'hA2; B = 8'hA; #100;
A = 8'hA2; B = 8'hB; #100;
A = 8'hA2; B = 8'hC; #100;
A = 8'hA2; B = 8'hD; #100;
A = 8'hA2; B = 8'hE; #100;
A = 8'hA2; B = 8'hF; #100;
A = 8'hA2; B = 8'h10; #100;
A = 8'hA2; B = 8'h11; #100;
A = 8'hA2; B = 8'h12; #100;
A = 8'hA2; B = 8'h13; #100;
A = 8'hA2; B = 8'h14; #100;
A = 8'hA2; B = 8'h15; #100;
A = 8'hA2; B = 8'h16; #100;
A = 8'hA2; B = 8'h17; #100;
A = 8'hA2; B = 8'h18; #100;
A = 8'hA2; B = 8'h19; #100;
A = 8'hA2; B = 8'h1A; #100;
A = 8'hA2; B = 8'h1B; #100;
A = 8'hA2; B = 8'h1C; #100;
A = 8'hA2; B = 8'h1D; #100;
A = 8'hA2; B = 8'h1E; #100;
A = 8'hA2; B = 8'h1F; #100;
A = 8'hA2; B = 8'h20; #100;
A = 8'hA2; B = 8'h21; #100;
A = 8'hA2; B = 8'h22; #100;
A = 8'hA2; B = 8'h23; #100;
A = 8'hA2; B = 8'h24; #100;
A = 8'hA2; B = 8'h25; #100;
A = 8'hA2; B = 8'h26; #100;
A = 8'hA2; B = 8'h27; #100;
A = 8'hA2; B = 8'h28; #100;
A = 8'hA2; B = 8'h29; #100;
A = 8'hA2; B = 8'h2A; #100;
A = 8'hA2; B = 8'h2B; #100;
A = 8'hA2; B = 8'h2C; #100;
A = 8'hA2; B = 8'h2D; #100;
A = 8'hA2; B = 8'h2E; #100;
A = 8'hA2; B = 8'h2F; #100;
A = 8'hA2; B = 8'h30; #100;
A = 8'hA2; B = 8'h31; #100;
A = 8'hA2; B = 8'h32; #100;
A = 8'hA2; B = 8'h33; #100;
A = 8'hA2; B = 8'h34; #100;
A = 8'hA2; B = 8'h35; #100;
A = 8'hA2; B = 8'h36; #100;
A = 8'hA2; B = 8'h37; #100;
A = 8'hA2; B = 8'h38; #100;
A = 8'hA2; B = 8'h39; #100;
A = 8'hA2; B = 8'h3A; #100;
A = 8'hA2; B = 8'h3B; #100;
A = 8'hA2; B = 8'h3C; #100;
A = 8'hA2; B = 8'h3D; #100;
A = 8'hA2; B = 8'h3E; #100;
A = 8'hA2; B = 8'h3F; #100;
A = 8'hA2; B = 8'h40; #100;
A = 8'hA2; B = 8'h41; #100;
A = 8'hA2; B = 8'h42; #100;
A = 8'hA2; B = 8'h43; #100;
A = 8'hA2; B = 8'h44; #100;
A = 8'hA2; B = 8'h45; #100;
A = 8'hA2; B = 8'h46; #100;
A = 8'hA2; B = 8'h47; #100;
A = 8'hA2; B = 8'h48; #100;
A = 8'hA2; B = 8'h49; #100;
A = 8'hA2; B = 8'h4A; #100;
A = 8'hA2; B = 8'h4B; #100;
A = 8'hA2; B = 8'h4C; #100;
A = 8'hA2; B = 8'h4D; #100;
A = 8'hA2; B = 8'h4E; #100;
A = 8'hA2; B = 8'h4F; #100;
A = 8'hA2; B = 8'h50; #100;
A = 8'hA2; B = 8'h51; #100;
A = 8'hA2; B = 8'h52; #100;
A = 8'hA2; B = 8'h53; #100;
A = 8'hA2; B = 8'h54; #100;
A = 8'hA2; B = 8'h55; #100;
A = 8'hA2; B = 8'h56; #100;
A = 8'hA2; B = 8'h57; #100;
A = 8'hA2; B = 8'h58; #100;
A = 8'hA2; B = 8'h59; #100;
A = 8'hA2; B = 8'h5A; #100;
A = 8'hA2; B = 8'h5B; #100;
A = 8'hA2; B = 8'h5C; #100;
A = 8'hA2; B = 8'h5D; #100;
A = 8'hA2; B = 8'h5E; #100;
A = 8'hA2; B = 8'h5F; #100;
A = 8'hA2; B = 8'h60; #100;
A = 8'hA2; B = 8'h61; #100;
A = 8'hA2; B = 8'h62; #100;
A = 8'hA2; B = 8'h63; #100;
A = 8'hA2; B = 8'h64; #100;
A = 8'hA2; B = 8'h65; #100;
A = 8'hA2; B = 8'h66; #100;
A = 8'hA2; B = 8'h67; #100;
A = 8'hA2; B = 8'h68; #100;
A = 8'hA2; B = 8'h69; #100;
A = 8'hA2; B = 8'h6A; #100;
A = 8'hA2; B = 8'h6B; #100;
A = 8'hA2; B = 8'h6C; #100;
A = 8'hA2; B = 8'h6D; #100;
A = 8'hA2; B = 8'h6E; #100;
A = 8'hA2; B = 8'h6F; #100;
A = 8'hA2; B = 8'h70; #100;
A = 8'hA2; B = 8'h71; #100;
A = 8'hA2; B = 8'h72; #100;
A = 8'hA2; B = 8'h73; #100;
A = 8'hA2; B = 8'h74; #100;
A = 8'hA2; B = 8'h75; #100;
A = 8'hA2; B = 8'h76; #100;
A = 8'hA2; B = 8'h77; #100;
A = 8'hA2; B = 8'h78; #100;
A = 8'hA2; B = 8'h79; #100;
A = 8'hA2; B = 8'h7A; #100;
A = 8'hA2; B = 8'h7B; #100;
A = 8'hA2; B = 8'h7C; #100;
A = 8'hA2; B = 8'h7D; #100;
A = 8'hA2; B = 8'h7E; #100;
A = 8'hA2; B = 8'h7F; #100;
A = 8'hA2; B = 8'h80; #100;
A = 8'hA2; B = 8'h81; #100;
A = 8'hA2; B = 8'h82; #100;
A = 8'hA2; B = 8'h83; #100;
A = 8'hA2; B = 8'h84; #100;
A = 8'hA2; B = 8'h85; #100;
A = 8'hA2; B = 8'h86; #100;
A = 8'hA2; B = 8'h87; #100;
A = 8'hA2; B = 8'h88; #100;
A = 8'hA2; B = 8'h89; #100;
A = 8'hA2; B = 8'h8A; #100;
A = 8'hA2; B = 8'h8B; #100;
A = 8'hA2; B = 8'h8C; #100;
A = 8'hA2; B = 8'h8D; #100;
A = 8'hA2; B = 8'h8E; #100;
A = 8'hA2; B = 8'h8F; #100;
A = 8'hA2; B = 8'h90; #100;
A = 8'hA2; B = 8'h91; #100;
A = 8'hA2; B = 8'h92; #100;
A = 8'hA2; B = 8'h93; #100;
A = 8'hA2; B = 8'h94; #100;
A = 8'hA2; B = 8'h95; #100;
A = 8'hA2; B = 8'h96; #100;
A = 8'hA2; B = 8'h97; #100;
A = 8'hA2; B = 8'h98; #100;
A = 8'hA2; B = 8'h99; #100;
A = 8'hA2; B = 8'h9A; #100;
A = 8'hA2; B = 8'h9B; #100;
A = 8'hA2; B = 8'h9C; #100;
A = 8'hA2; B = 8'h9D; #100;
A = 8'hA2; B = 8'h9E; #100;
A = 8'hA2; B = 8'h9F; #100;
A = 8'hA2; B = 8'hA0; #100;
A = 8'hA2; B = 8'hA1; #100;
A = 8'hA2; B = 8'hA2; #100;
A = 8'hA2; B = 8'hA3; #100;
A = 8'hA2; B = 8'hA4; #100;
A = 8'hA2; B = 8'hA5; #100;
A = 8'hA2; B = 8'hA6; #100;
A = 8'hA2; B = 8'hA7; #100;
A = 8'hA2; B = 8'hA8; #100;
A = 8'hA2; B = 8'hA9; #100;
A = 8'hA2; B = 8'hAA; #100;
A = 8'hA2; B = 8'hAB; #100;
A = 8'hA2; B = 8'hAC; #100;
A = 8'hA2; B = 8'hAD; #100;
A = 8'hA2; B = 8'hAE; #100;
A = 8'hA2; B = 8'hAF; #100;
A = 8'hA2; B = 8'hB0; #100;
A = 8'hA2; B = 8'hB1; #100;
A = 8'hA2; B = 8'hB2; #100;
A = 8'hA2; B = 8'hB3; #100;
A = 8'hA2; B = 8'hB4; #100;
A = 8'hA2; B = 8'hB5; #100;
A = 8'hA2; B = 8'hB6; #100;
A = 8'hA2; B = 8'hB7; #100;
A = 8'hA2; B = 8'hB8; #100;
A = 8'hA2; B = 8'hB9; #100;
A = 8'hA2; B = 8'hBA; #100;
A = 8'hA2; B = 8'hBB; #100;
A = 8'hA2; B = 8'hBC; #100;
A = 8'hA2; B = 8'hBD; #100;
A = 8'hA2; B = 8'hBE; #100;
A = 8'hA2; B = 8'hBF; #100;
A = 8'hA2; B = 8'hC0; #100;
A = 8'hA2; B = 8'hC1; #100;
A = 8'hA2; B = 8'hC2; #100;
A = 8'hA2; B = 8'hC3; #100;
A = 8'hA2; B = 8'hC4; #100;
A = 8'hA2; B = 8'hC5; #100;
A = 8'hA2; B = 8'hC6; #100;
A = 8'hA2; B = 8'hC7; #100;
A = 8'hA2; B = 8'hC8; #100;
A = 8'hA2; B = 8'hC9; #100;
A = 8'hA2; B = 8'hCA; #100;
A = 8'hA2; B = 8'hCB; #100;
A = 8'hA2; B = 8'hCC; #100;
A = 8'hA2; B = 8'hCD; #100;
A = 8'hA2; B = 8'hCE; #100;
A = 8'hA2; B = 8'hCF; #100;
A = 8'hA2; B = 8'hD0; #100;
A = 8'hA2; B = 8'hD1; #100;
A = 8'hA2; B = 8'hD2; #100;
A = 8'hA2; B = 8'hD3; #100;
A = 8'hA2; B = 8'hD4; #100;
A = 8'hA2; B = 8'hD5; #100;
A = 8'hA2; B = 8'hD6; #100;
A = 8'hA2; B = 8'hD7; #100;
A = 8'hA2; B = 8'hD8; #100;
A = 8'hA2; B = 8'hD9; #100;
A = 8'hA2; B = 8'hDA; #100;
A = 8'hA2; B = 8'hDB; #100;
A = 8'hA2; B = 8'hDC; #100;
A = 8'hA2; B = 8'hDD; #100;
A = 8'hA2; B = 8'hDE; #100;
A = 8'hA2; B = 8'hDF; #100;
A = 8'hA2; B = 8'hE0; #100;
A = 8'hA2; B = 8'hE1; #100;
A = 8'hA2; B = 8'hE2; #100;
A = 8'hA2; B = 8'hE3; #100;
A = 8'hA2; B = 8'hE4; #100;
A = 8'hA2; B = 8'hE5; #100;
A = 8'hA2; B = 8'hE6; #100;
A = 8'hA2; B = 8'hE7; #100;
A = 8'hA2; B = 8'hE8; #100;
A = 8'hA2; B = 8'hE9; #100;
A = 8'hA2; B = 8'hEA; #100;
A = 8'hA2; B = 8'hEB; #100;
A = 8'hA2; B = 8'hEC; #100;
A = 8'hA2; B = 8'hED; #100;
A = 8'hA2; B = 8'hEE; #100;
A = 8'hA2; B = 8'hEF; #100;
A = 8'hA2; B = 8'hF0; #100;
A = 8'hA2; B = 8'hF1; #100;
A = 8'hA2; B = 8'hF2; #100;
A = 8'hA2; B = 8'hF3; #100;
A = 8'hA2; B = 8'hF4; #100;
A = 8'hA2; B = 8'hF5; #100;
A = 8'hA2; B = 8'hF6; #100;
A = 8'hA2; B = 8'hF7; #100;
A = 8'hA2; B = 8'hF8; #100;
A = 8'hA2; B = 8'hF9; #100;
A = 8'hA2; B = 8'hFA; #100;
A = 8'hA2; B = 8'hFB; #100;
A = 8'hA2; B = 8'hFC; #100;
A = 8'hA2; B = 8'hFD; #100;
A = 8'hA2; B = 8'hFE; #100;
A = 8'hA2; B = 8'hFF; #100;
A = 8'hA3; B = 8'h0; #100;
A = 8'hA3; B = 8'h1; #100;
A = 8'hA3; B = 8'h2; #100;
A = 8'hA3; B = 8'h3; #100;
A = 8'hA3; B = 8'h4; #100;
A = 8'hA3; B = 8'h5; #100;
A = 8'hA3; B = 8'h6; #100;
A = 8'hA3; B = 8'h7; #100;
A = 8'hA3; B = 8'h8; #100;
A = 8'hA3; B = 8'h9; #100;
A = 8'hA3; B = 8'hA; #100;
A = 8'hA3; B = 8'hB; #100;
A = 8'hA3; B = 8'hC; #100;
A = 8'hA3; B = 8'hD; #100;
A = 8'hA3; B = 8'hE; #100;
A = 8'hA3; B = 8'hF; #100;
A = 8'hA3; B = 8'h10; #100;
A = 8'hA3; B = 8'h11; #100;
A = 8'hA3; B = 8'h12; #100;
A = 8'hA3; B = 8'h13; #100;
A = 8'hA3; B = 8'h14; #100;
A = 8'hA3; B = 8'h15; #100;
A = 8'hA3; B = 8'h16; #100;
A = 8'hA3; B = 8'h17; #100;
A = 8'hA3; B = 8'h18; #100;
A = 8'hA3; B = 8'h19; #100;
A = 8'hA3; B = 8'h1A; #100;
A = 8'hA3; B = 8'h1B; #100;
A = 8'hA3; B = 8'h1C; #100;
A = 8'hA3; B = 8'h1D; #100;
A = 8'hA3; B = 8'h1E; #100;
A = 8'hA3; B = 8'h1F; #100;
A = 8'hA3; B = 8'h20; #100;
A = 8'hA3; B = 8'h21; #100;
A = 8'hA3; B = 8'h22; #100;
A = 8'hA3; B = 8'h23; #100;
A = 8'hA3; B = 8'h24; #100;
A = 8'hA3; B = 8'h25; #100;
A = 8'hA3; B = 8'h26; #100;
A = 8'hA3; B = 8'h27; #100;
A = 8'hA3; B = 8'h28; #100;
A = 8'hA3; B = 8'h29; #100;
A = 8'hA3; B = 8'h2A; #100;
A = 8'hA3; B = 8'h2B; #100;
A = 8'hA3; B = 8'h2C; #100;
A = 8'hA3; B = 8'h2D; #100;
A = 8'hA3; B = 8'h2E; #100;
A = 8'hA3; B = 8'h2F; #100;
A = 8'hA3; B = 8'h30; #100;
A = 8'hA3; B = 8'h31; #100;
A = 8'hA3; B = 8'h32; #100;
A = 8'hA3; B = 8'h33; #100;
A = 8'hA3; B = 8'h34; #100;
A = 8'hA3; B = 8'h35; #100;
A = 8'hA3; B = 8'h36; #100;
A = 8'hA3; B = 8'h37; #100;
A = 8'hA3; B = 8'h38; #100;
A = 8'hA3; B = 8'h39; #100;
A = 8'hA3; B = 8'h3A; #100;
A = 8'hA3; B = 8'h3B; #100;
A = 8'hA3; B = 8'h3C; #100;
A = 8'hA3; B = 8'h3D; #100;
A = 8'hA3; B = 8'h3E; #100;
A = 8'hA3; B = 8'h3F; #100;
A = 8'hA3; B = 8'h40; #100;
A = 8'hA3; B = 8'h41; #100;
A = 8'hA3; B = 8'h42; #100;
A = 8'hA3; B = 8'h43; #100;
A = 8'hA3; B = 8'h44; #100;
A = 8'hA3; B = 8'h45; #100;
A = 8'hA3; B = 8'h46; #100;
A = 8'hA3; B = 8'h47; #100;
A = 8'hA3; B = 8'h48; #100;
A = 8'hA3; B = 8'h49; #100;
A = 8'hA3; B = 8'h4A; #100;
A = 8'hA3; B = 8'h4B; #100;
A = 8'hA3; B = 8'h4C; #100;
A = 8'hA3; B = 8'h4D; #100;
A = 8'hA3; B = 8'h4E; #100;
A = 8'hA3; B = 8'h4F; #100;
A = 8'hA3; B = 8'h50; #100;
A = 8'hA3; B = 8'h51; #100;
A = 8'hA3; B = 8'h52; #100;
A = 8'hA3; B = 8'h53; #100;
A = 8'hA3; B = 8'h54; #100;
A = 8'hA3; B = 8'h55; #100;
A = 8'hA3; B = 8'h56; #100;
A = 8'hA3; B = 8'h57; #100;
A = 8'hA3; B = 8'h58; #100;
A = 8'hA3; B = 8'h59; #100;
A = 8'hA3; B = 8'h5A; #100;
A = 8'hA3; B = 8'h5B; #100;
A = 8'hA3; B = 8'h5C; #100;
A = 8'hA3; B = 8'h5D; #100;
A = 8'hA3; B = 8'h5E; #100;
A = 8'hA3; B = 8'h5F; #100;
A = 8'hA3; B = 8'h60; #100;
A = 8'hA3; B = 8'h61; #100;
A = 8'hA3; B = 8'h62; #100;
A = 8'hA3; B = 8'h63; #100;
A = 8'hA3; B = 8'h64; #100;
A = 8'hA3; B = 8'h65; #100;
A = 8'hA3; B = 8'h66; #100;
A = 8'hA3; B = 8'h67; #100;
A = 8'hA3; B = 8'h68; #100;
A = 8'hA3; B = 8'h69; #100;
A = 8'hA3; B = 8'h6A; #100;
A = 8'hA3; B = 8'h6B; #100;
A = 8'hA3; B = 8'h6C; #100;
A = 8'hA3; B = 8'h6D; #100;
A = 8'hA3; B = 8'h6E; #100;
A = 8'hA3; B = 8'h6F; #100;
A = 8'hA3; B = 8'h70; #100;
A = 8'hA3; B = 8'h71; #100;
A = 8'hA3; B = 8'h72; #100;
A = 8'hA3; B = 8'h73; #100;
A = 8'hA3; B = 8'h74; #100;
A = 8'hA3; B = 8'h75; #100;
A = 8'hA3; B = 8'h76; #100;
A = 8'hA3; B = 8'h77; #100;
A = 8'hA3; B = 8'h78; #100;
A = 8'hA3; B = 8'h79; #100;
A = 8'hA3; B = 8'h7A; #100;
A = 8'hA3; B = 8'h7B; #100;
A = 8'hA3; B = 8'h7C; #100;
A = 8'hA3; B = 8'h7D; #100;
A = 8'hA3; B = 8'h7E; #100;
A = 8'hA3; B = 8'h7F; #100;
A = 8'hA3; B = 8'h80; #100;
A = 8'hA3; B = 8'h81; #100;
A = 8'hA3; B = 8'h82; #100;
A = 8'hA3; B = 8'h83; #100;
A = 8'hA3; B = 8'h84; #100;
A = 8'hA3; B = 8'h85; #100;
A = 8'hA3; B = 8'h86; #100;
A = 8'hA3; B = 8'h87; #100;
A = 8'hA3; B = 8'h88; #100;
A = 8'hA3; B = 8'h89; #100;
A = 8'hA3; B = 8'h8A; #100;
A = 8'hA3; B = 8'h8B; #100;
A = 8'hA3; B = 8'h8C; #100;
A = 8'hA3; B = 8'h8D; #100;
A = 8'hA3; B = 8'h8E; #100;
A = 8'hA3; B = 8'h8F; #100;
A = 8'hA3; B = 8'h90; #100;
A = 8'hA3; B = 8'h91; #100;
A = 8'hA3; B = 8'h92; #100;
A = 8'hA3; B = 8'h93; #100;
A = 8'hA3; B = 8'h94; #100;
A = 8'hA3; B = 8'h95; #100;
A = 8'hA3; B = 8'h96; #100;
A = 8'hA3; B = 8'h97; #100;
A = 8'hA3; B = 8'h98; #100;
A = 8'hA3; B = 8'h99; #100;
A = 8'hA3; B = 8'h9A; #100;
A = 8'hA3; B = 8'h9B; #100;
A = 8'hA3; B = 8'h9C; #100;
A = 8'hA3; B = 8'h9D; #100;
A = 8'hA3; B = 8'h9E; #100;
A = 8'hA3; B = 8'h9F; #100;
A = 8'hA3; B = 8'hA0; #100;
A = 8'hA3; B = 8'hA1; #100;
A = 8'hA3; B = 8'hA2; #100;
A = 8'hA3; B = 8'hA3; #100;
A = 8'hA3; B = 8'hA4; #100;
A = 8'hA3; B = 8'hA5; #100;
A = 8'hA3; B = 8'hA6; #100;
A = 8'hA3; B = 8'hA7; #100;
A = 8'hA3; B = 8'hA8; #100;
A = 8'hA3; B = 8'hA9; #100;
A = 8'hA3; B = 8'hAA; #100;
A = 8'hA3; B = 8'hAB; #100;
A = 8'hA3; B = 8'hAC; #100;
A = 8'hA3; B = 8'hAD; #100;
A = 8'hA3; B = 8'hAE; #100;
A = 8'hA3; B = 8'hAF; #100;
A = 8'hA3; B = 8'hB0; #100;
A = 8'hA3; B = 8'hB1; #100;
A = 8'hA3; B = 8'hB2; #100;
A = 8'hA3; B = 8'hB3; #100;
A = 8'hA3; B = 8'hB4; #100;
A = 8'hA3; B = 8'hB5; #100;
A = 8'hA3; B = 8'hB6; #100;
A = 8'hA3; B = 8'hB7; #100;
A = 8'hA3; B = 8'hB8; #100;
A = 8'hA3; B = 8'hB9; #100;
A = 8'hA3; B = 8'hBA; #100;
A = 8'hA3; B = 8'hBB; #100;
A = 8'hA3; B = 8'hBC; #100;
A = 8'hA3; B = 8'hBD; #100;
A = 8'hA3; B = 8'hBE; #100;
A = 8'hA3; B = 8'hBF; #100;
A = 8'hA3; B = 8'hC0; #100;
A = 8'hA3; B = 8'hC1; #100;
A = 8'hA3; B = 8'hC2; #100;
A = 8'hA3; B = 8'hC3; #100;
A = 8'hA3; B = 8'hC4; #100;
A = 8'hA3; B = 8'hC5; #100;
A = 8'hA3; B = 8'hC6; #100;
A = 8'hA3; B = 8'hC7; #100;
A = 8'hA3; B = 8'hC8; #100;
A = 8'hA3; B = 8'hC9; #100;
A = 8'hA3; B = 8'hCA; #100;
A = 8'hA3; B = 8'hCB; #100;
A = 8'hA3; B = 8'hCC; #100;
A = 8'hA3; B = 8'hCD; #100;
A = 8'hA3; B = 8'hCE; #100;
A = 8'hA3; B = 8'hCF; #100;
A = 8'hA3; B = 8'hD0; #100;
A = 8'hA3; B = 8'hD1; #100;
A = 8'hA3; B = 8'hD2; #100;
A = 8'hA3; B = 8'hD3; #100;
A = 8'hA3; B = 8'hD4; #100;
A = 8'hA3; B = 8'hD5; #100;
A = 8'hA3; B = 8'hD6; #100;
A = 8'hA3; B = 8'hD7; #100;
A = 8'hA3; B = 8'hD8; #100;
A = 8'hA3; B = 8'hD9; #100;
A = 8'hA3; B = 8'hDA; #100;
A = 8'hA3; B = 8'hDB; #100;
A = 8'hA3; B = 8'hDC; #100;
A = 8'hA3; B = 8'hDD; #100;
A = 8'hA3; B = 8'hDE; #100;
A = 8'hA3; B = 8'hDF; #100;
A = 8'hA3; B = 8'hE0; #100;
A = 8'hA3; B = 8'hE1; #100;
A = 8'hA3; B = 8'hE2; #100;
A = 8'hA3; B = 8'hE3; #100;
A = 8'hA3; B = 8'hE4; #100;
A = 8'hA3; B = 8'hE5; #100;
A = 8'hA3; B = 8'hE6; #100;
A = 8'hA3; B = 8'hE7; #100;
A = 8'hA3; B = 8'hE8; #100;
A = 8'hA3; B = 8'hE9; #100;
A = 8'hA3; B = 8'hEA; #100;
A = 8'hA3; B = 8'hEB; #100;
A = 8'hA3; B = 8'hEC; #100;
A = 8'hA3; B = 8'hED; #100;
A = 8'hA3; B = 8'hEE; #100;
A = 8'hA3; B = 8'hEF; #100;
A = 8'hA3; B = 8'hF0; #100;
A = 8'hA3; B = 8'hF1; #100;
A = 8'hA3; B = 8'hF2; #100;
A = 8'hA3; B = 8'hF3; #100;
A = 8'hA3; B = 8'hF4; #100;
A = 8'hA3; B = 8'hF5; #100;
A = 8'hA3; B = 8'hF6; #100;
A = 8'hA3; B = 8'hF7; #100;
A = 8'hA3; B = 8'hF8; #100;
A = 8'hA3; B = 8'hF9; #100;
A = 8'hA3; B = 8'hFA; #100;
A = 8'hA3; B = 8'hFB; #100;
A = 8'hA3; B = 8'hFC; #100;
A = 8'hA3; B = 8'hFD; #100;
A = 8'hA3; B = 8'hFE; #100;
A = 8'hA3; B = 8'hFF; #100;
A = 8'hA4; B = 8'h0; #100;
A = 8'hA4; B = 8'h1; #100;
A = 8'hA4; B = 8'h2; #100;
A = 8'hA4; B = 8'h3; #100;
A = 8'hA4; B = 8'h4; #100;
A = 8'hA4; B = 8'h5; #100;
A = 8'hA4; B = 8'h6; #100;
A = 8'hA4; B = 8'h7; #100;
A = 8'hA4; B = 8'h8; #100;
A = 8'hA4; B = 8'h9; #100;
A = 8'hA4; B = 8'hA; #100;
A = 8'hA4; B = 8'hB; #100;
A = 8'hA4; B = 8'hC; #100;
A = 8'hA4; B = 8'hD; #100;
A = 8'hA4; B = 8'hE; #100;
A = 8'hA4; B = 8'hF; #100;
A = 8'hA4; B = 8'h10; #100;
A = 8'hA4; B = 8'h11; #100;
A = 8'hA4; B = 8'h12; #100;
A = 8'hA4; B = 8'h13; #100;
A = 8'hA4; B = 8'h14; #100;
A = 8'hA4; B = 8'h15; #100;
A = 8'hA4; B = 8'h16; #100;
A = 8'hA4; B = 8'h17; #100;
A = 8'hA4; B = 8'h18; #100;
A = 8'hA4; B = 8'h19; #100;
A = 8'hA4; B = 8'h1A; #100;
A = 8'hA4; B = 8'h1B; #100;
A = 8'hA4; B = 8'h1C; #100;
A = 8'hA4; B = 8'h1D; #100;
A = 8'hA4; B = 8'h1E; #100;
A = 8'hA4; B = 8'h1F; #100;
A = 8'hA4; B = 8'h20; #100;
A = 8'hA4; B = 8'h21; #100;
A = 8'hA4; B = 8'h22; #100;
A = 8'hA4; B = 8'h23; #100;
A = 8'hA4; B = 8'h24; #100;
A = 8'hA4; B = 8'h25; #100;
A = 8'hA4; B = 8'h26; #100;
A = 8'hA4; B = 8'h27; #100;
A = 8'hA4; B = 8'h28; #100;
A = 8'hA4; B = 8'h29; #100;
A = 8'hA4; B = 8'h2A; #100;
A = 8'hA4; B = 8'h2B; #100;
A = 8'hA4; B = 8'h2C; #100;
A = 8'hA4; B = 8'h2D; #100;
A = 8'hA4; B = 8'h2E; #100;
A = 8'hA4; B = 8'h2F; #100;
A = 8'hA4; B = 8'h30; #100;
A = 8'hA4; B = 8'h31; #100;
A = 8'hA4; B = 8'h32; #100;
A = 8'hA4; B = 8'h33; #100;
A = 8'hA4; B = 8'h34; #100;
A = 8'hA4; B = 8'h35; #100;
A = 8'hA4; B = 8'h36; #100;
A = 8'hA4; B = 8'h37; #100;
A = 8'hA4; B = 8'h38; #100;
A = 8'hA4; B = 8'h39; #100;
A = 8'hA4; B = 8'h3A; #100;
A = 8'hA4; B = 8'h3B; #100;
A = 8'hA4; B = 8'h3C; #100;
A = 8'hA4; B = 8'h3D; #100;
A = 8'hA4; B = 8'h3E; #100;
A = 8'hA4; B = 8'h3F; #100;
A = 8'hA4; B = 8'h40; #100;
A = 8'hA4; B = 8'h41; #100;
A = 8'hA4; B = 8'h42; #100;
A = 8'hA4; B = 8'h43; #100;
A = 8'hA4; B = 8'h44; #100;
A = 8'hA4; B = 8'h45; #100;
A = 8'hA4; B = 8'h46; #100;
A = 8'hA4; B = 8'h47; #100;
A = 8'hA4; B = 8'h48; #100;
A = 8'hA4; B = 8'h49; #100;
A = 8'hA4; B = 8'h4A; #100;
A = 8'hA4; B = 8'h4B; #100;
A = 8'hA4; B = 8'h4C; #100;
A = 8'hA4; B = 8'h4D; #100;
A = 8'hA4; B = 8'h4E; #100;
A = 8'hA4; B = 8'h4F; #100;
A = 8'hA4; B = 8'h50; #100;
A = 8'hA4; B = 8'h51; #100;
A = 8'hA4; B = 8'h52; #100;
A = 8'hA4; B = 8'h53; #100;
A = 8'hA4; B = 8'h54; #100;
A = 8'hA4; B = 8'h55; #100;
A = 8'hA4; B = 8'h56; #100;
A = 8'hA4; B = 8'h57; #100;
A = 8'hA4; B = 8'h58; #100;
A = 8'hA4; B = 8'h59; #100;
A = 8'hA4; B = 8'h5A; #100;
A = 8'hA4; B = 8'h5B; #100;
A = 8'hA4; B = 8'h5C; #100;
A = 8'hA4; B = 8'h5D; #100;
A = 8'hA4; B = 8'h5E; #100;
A = 8'hA4; B = 8'h5F; #100;
A = 8'hA4; B = 8'h60; #100;
A = 8'hA4; B = 8'h61; #100;
A = 8'hA4; B = 8'h62; #100;
A = 8'hA4; B = 8'h63; #100;
A = 8'hA4; B = 8'h64; #100;
A = 8'hA4; B = 8'h65; #100;
A = 8'hA4; B = 8'h66; #100;
A = 8'hA4; B = 8'h67; #100;
A = 8'hA4; B = 8'h68; #100;
A = 8'hA4; B = 8'h69; #100;
A = 8'hA4; B = 8'h6A; #100;
A = 8'hA4; B = 8'h6B; #100;
A = 8'hA4; B = 8'h6C; #100;
A = 8'hA4; B = 8'h6D; #100;
A = 8'hA4; B = 8'h6E; #100;
A = 8'hA4; B = 8'h6F; #100;
A = 8'hA4; B = 8'h70; #100;
A = 8'hA4; B = 8'h71; #100;
A = 8'hA4; B = 8'h72; #100;
A = 8'hA4; B = 8'h73; #100;
A = 8'hA4; B = 8'h74; #100;
A = 8'hA4; B = 8'h75; #100;
A = 8'hA4; B = 8'h76; #100;
A = 8'hA4; B = 8'h77; #100;
A = 8'hA4; B = 8'h78; #100;
A = 8'hA4; B = 8'h79; #100;
A = 8'hA4; B = 8'h7A; #100;
A = 8'hA4; B = 8'h7B; #100;
A = 8'hA4; B = 8'h7C; #100;
A = 8'hA4; B = 8'h7D; #100;
A = 8'hA4; B = 8'h7E; #100;
A = 8'hA4; B = 8'h7F; #100;
A = 8'hA4; B = 8'h80; #100;
A = 8'hA4; B = 8'h81; #100;
A = 8'hA4; B = 8'h82; #100;
A = 8'hA4; B = 8'h83; #100;
A = 8'hA4; B = 8'h84; #100;
A = 8'hA4; B = 8'h85; #100;
A = 8'hA4; B = 8'h86; #100;
A = 8'hA4; B = 8'h87; #100;
A = 8'hA4; B = 8'h88; #100;
A = 8'hA4; B = 8'h89; #100;
A = 8'hA4; B = 8'h8A; #100;
A = 8'hA4; B = 8'h8B; #100;
A = 8'hA4; B = 8'h8C; #100;
A = 8'hA4; B = 8'h8D; #100;
A = 8'hA4; B = 8'h8E; #100;
A = 8'hA4; B = 8'h8F; #100;
A = 8'hA4; B = 8'h90; #100;
A = 8'hA4; B = 8'h91; #100;
A = 8'hA4; B = 8'h92; #100;
A = 8'hA4; B = 8'h93; #100;
A = 8'hA4; B = 8'h94; #100;
A = 8'hA4; B = 8'h95; #100;
A = 8'hA4; B = 8'h96; #100;
A = 8'hA4; B = 8'h97; #100;
A = 8'hA4; B = 8'h98; #100;
A = 8'hA4; B = 8'h99; #100;
A = 8'hA4; B = 8'h9A; #100;
A = 8'hA4; B = 8'h9B; #100;
A = 8'hA4; B = 8'h9C; #100;
A = 8'hA4; B = 8'h9D; #100;
A = 8'hA4; B = 8'h9E; #100;
A = 8'hA4; B = 8'h9F; #100;
A = 8'hA4; B = 8'hA0; #100;
A = 8'hA4; B = 8'hA1; #100;
A = 8'hA4; B = 8'hA2; #100;
A = 8'hA4; B = 8'hA3; #100;
A = 8'hA4; B = 8'hA4; #100;
A = 8'hA4; B = 8'hA5; #100;
A = 8'hA4; B = 8'hA6; #100;
A = 8'hA4; B = 8'hA7; #100;
A = 8'hA4; B = 8'hA8; #100;
A = 8'hA4; B = 8'hA9; #100;
A = 8'hA4; B = 8'hAA; #100;
A = 8'hA4; B = 8'hAB; #100;
A = 8'hA4; B = 8'hAC; #100;
A = 8'hA4; B = 8'hAD; #100;
A = 8'hA4; B = 8'hAE; #100;
A = 8'hA4; B = 8'hAF; #100;
A = 8'hA4; B = 8'hB0; #100;
A = 8'hA4; B = 8'hB1; #100;
A = 8'hA4; B = 8'hB2; #100;
A = 8'hA4; B = 8'hB3; #100;
A = 8'hA4; B = 8'hB4; #100;
A = 8'hA4; B = 8'hB5; #100;
A = 8'hA4; B = 8'hB6; #100;
A = 8'hA4; B = 8'hB7; #100;
A = 8'hA4; B = 8'hB8; #100;
A = 8'hA4; B = 8'hB9; #100;
A = 8'hA4; B = 8'hBA; #100;
A = 8'hA4; B = 8'hBB; #100;
A = 8'hA4; B = 8'hBC; #100;
A = 8'hA4; B = 8'hBD; #100;
A = 8'hA4; B = 8'hBE; #100;
A = 8'hA4; B = 8'hBF; #100;
A = 8'hA4; B = 8'hC0; #100;
A = 8'hA4; B = 8'hC1; #100;
A = 8'hA4; B = 8'hC2; #100;
A = 8'hA4; B = 8'hC3; #100;
A = 8'hA4; B = 8'hC4; #100;
A = 8'hA4; B = 8'hC5; #100;
A = 8'hA4; B = 8'hC6; #100;
A = 8'hA4; B = 8'hC7; #100;
A = 8'hA4; B = 8'hC8; #100;
A = 8'hA4; B = 8'hC9; #100;
A = 8'hA4; B = 8'hCA; #100;
A = 8'hA4; B = 8'hCB; #100;
A = 8'hA4; B = 8'hCC; #100;
A = 8'hA4; B = 8'hCD; #100;
A = 8'hA4; B = 8'hCE; #100;
A = 8'hA4; B = 8'hCF; #100;
A = 8'hA4; B = 8'hD0; #100;
A = 8'hA4; B = 8'hD1; #100;
A = 8'hA4; B = 8'hD2; #100;
A = 8'hA4; B = 8'hD3; #100;
A = 8'hA4; B = 8'hD4; #100;
A = 8'hA4; B = 8'hD5; #100;
A = 8'hA4; B = 8'hD6; #100;
A = 8'hA4; B = 8'hD7; #100;
A = 8'hA4; B = 8'hD8; #100;
A = 8'hA4; B = 8'hD9; #100;
A = 8'hA4; B = 8'hDA; #100;
A = 8'hA4; B = 8'hDB; #100;
A = 8'hA4; B = 8'hDC; #100;
A = 8'hA4; B = 8'hDD; #100;
A = 8'hA4; B = 8'hDE; #100;
A = 8'hA4; B = 8'hDF; #100;
A = 8'hA4; B = 8'hE0; #100;
A = 8'hA4; B = 8'hE1; #100;
A = 8'hA4; B = 8'hE2; #100;
A = 8'hA4; B = 8'hE3; #100;
A = 8'hA4; B = 8'hE4; #100;
A = 8'hA4; B = 8'hE5; #100;
A = 8'hA4; B = 8'hE6; #100;
A = 8'hA4; B = 8'hE7; #100;
A = 8'hA4; B = 8'hE8; #100;
A = 8'hA4; B = 8'hE9; #100;
A = 8'hA4; B = 8'hEA; #100;
A = 8'hA4; B = 8'hEB; #100;
A = 8'hA4; B = 8'hEC; #100;
A = 8'hA4; B = 8'hED; #100;
A = 8'hA4; B = 8'hEE; #100;
A = 8'hA4; B = 8'hEF; #100;
A = 8'hA4; B = 8'hF0; #100;
A = 8'hA4; B = 8'hF1; #100;
A = 8'hA4; B = 8'hF2; #100;
A = 8'hA4; B = 8'hF3; #100;
A = 8'hA4; B = 8'hF4; #100;
A = 8'hA4; B = 8'hF5; #100;
A = 8'hA4; B = 8'hF6; #100;
A = 8'hA4; B = 8'hF7; #100;
A = 8'hA4; B = 8'hF8; #100;
A = 8'hA4; B = 8'hF9; #100;
A = 8'hA4; B = 8'hFA; #100;
A = 8'hA4; B = 8'hFB; #100;
A = 8'hA4; B = 8'hFC; #100;
A = 8'hA4; B = 8'hFD; #100;
A = 8'hA4; B = 8'hFE; #100;
A = 8'hA4; B = 8'hFF; #100;
A = 8'hA5; B = 8'h0; #100;
A = 8'hA5; B = 8'h1; #100;
A = 8'hA5; B = 8'h2; #100;
A = 8'hA5; B = 8'h3; #100;
A = 8'hA5; B = 8'h4; #100;
A = 8'hA5; B = 8'h5; #100;
A = 8'hA5; B = 8'h6; #100;
A = 8'hA5; B = 8'h7; #100;
A = 8'hA5; B = 8'h8; #100;
A = 8'hA5; B = 8'h9; #100;
A = 8'hA5; B = 8'hA; #100;
A = 8'hA5; B = 8'hB; #100;
A = 8'hA5; B = 8'hC; #100;
A = 8'hA5; B = 8'hD; #100;
A = 8'hA5; B = 8'hE; #100;
A = 8'hA5; B = 8'hF; #100;
A = 8'hA5; B = 8'h10; #100;
A = 8'hA5; B = 8'h11; #100;
A = 8'hA5; B = 8'h12; #100;
A = 8'hA5; B = 8'h13; #100;
A = 8'hA5; B = 8'h14; #100;
A = 8'hA5; B = 8'h15; #100;
A = 8'hA5; B = 8'h16; #100;
A = 8'hA5; B = 8'h17; #100;
A = 8'hA5; B = 8'h18; #100;
A = 8'hA5; B = 8'h19; #100;
A = 8'hA5; B = 8'h1A; #100;
A = 8'hA5; B = 8'h1B; #100;
A = 8'hA5; B = 8'h1C; #100;
A = 8'hA5; B = 8'h1D; #100;
A = 8'hA5; B = 8'h1E; #100;
A = 8'hA5; B = 8'h1F; #100;
A = 8'hA5; B = 8'h20; #100;
A = 8'hA5; B = 8'h21; #100;
A = 8'hA5; B = 8'h22; #100;
A = 8'hA5; B = 8'h23; #100;
A = 8'hA5; B = 8'h24; #100;
A = 8'hA5; B = 8'h25; #100;
A = 8'hA5; B = 8'h26; #100;
A = 8'hA5; B = 8'h27; #100;
A = 8'hA5; B = 8'h28; #100;
A = 8'hA5; B = 8'h29; #100;
A = 8'hA5; B = 8'h2A; #100;
A = 8'hA5; B = 8'h2B; #100;
A = 8'hA5; B = 8'h2C; #100;
A = 8'hA5; B = 8'h2D; #100;
A = 8'hA5; B = 8'h2E; #100;
A = 8'hA5; B = 8'h2F; #100;
A = 8'hA5; B = 8'h30; #100;
A = 8'hA5; B = 8'h31; #100;
A = 8'hA5; B = 8'h32; #100;
A = 8'hA5; B = 8'h33; #100;
A = 8'hA5; B = 8'h34; #100;
A = 8'hA5; B = 8'h35; #100;
A = 8'hA5; B = 8'h36; #100;
A = 8'hA5; B = 8'h37; #100;
A = 8'hA5; B = 8'h38; #100;
A = 8'hA5; B = 8'h39; #100;
A = 8'hA5; B = 8'h3A; #100;
A = 8'hA5; B = 8'h3B; #100;
A = 8'hA5; B = 8'h3C; #100;
A = 8'hA5; B = 8'h3D; #100;
A = 8'hA5; B = 8'h3E; #100;
A = 8'hA5; B = 8'h3F; #100;
A = 8'hA5; B = 8'h40; #100;
A = 8'hA5; B = 8'h41; #100;
A = 8'hA5; B = 8'h42; #100;
A = 8'hA5; B = 8'h43; #100;
A = 8'hA5; B = 8'h44; #100;
A = 8'hA5; B = 8'h45; #100;
A = 8'hA5; B = 8'h46; #100;
A = 8'hA5; B = 8'h47; #100;
A = 8'hA5; B = 8'h48; #100;
A = 8'hA5; B = 8'h49; #100;
A = 8'hA5; B = 8'h4A; #100;
A = 8'hA5; B = 8'h4B; #100;
A = 8'hA5; B = 8'h4C; #100;
A = 8'hA5; B = 8'h4D; #100;
A = 8'hA5; B = 8'h4E; #100;
A = 8'hA5; B = 8'h4F; #100;
A = 8'hA5; B = 8'h50; #100;
A = 8'hA5; B = 8'h51; #100;
A = 8'hA5; B = 8'h52; #100;
A = 8'hA5; B = 8'h53; #100;
A = 8'hA5; B = 8'h54; #100;
A = 8'hA5; B = 8'h55; #100;
A = 8'hA5; B = 8'h56; #100;
A = 8'hA5; B = 8'h57; #100;
A = 8'hA5; B = 8'h58; #100;
A = 8'hA5; B = 8'h59; #100;
A = 8'hA5; B = 8'h5A; #100;
A = 8'hA5; B = 8'h5B; #100;
A = 8'hA5; B = 8'h5C; #100;
A = 8'hA5; B = 8'h5D; #100;
A = 8'hA5; B = 8'h5E; #100;
A = 8'hA5; B = 8'h5F; #100;
A = 8'hA5; B = 8'h60; #100;
A = 8'hA5; B = 8'h61; #100;
A = 8'hA5; B = 8'h62; #100;
A = 8'hA5; B = 8'h63; #100;
A = 8'hA5; B = 8'h64; #100;
A = 8'hA5; B = 8'h65; #100;
A = 8'hA5; B = 8'h66; #100;
A = 8'hA5; B = 8'h67; #100;
A = 8'hA5; B = 8'h68; #100;
A = 8'hA5; B = 8'h69; #100;
A = 8'hA5; B = 8'h6A; #100;
A = 8'hA5; B = 8'h6B; #100;
A = 8'hA5; B = 8'h6C; #100;
A = 8'hA5; B = 8'h6D; #100;
A = 8'hA5; B = 8'h6E; #100;
A = 8'hA5; B = 8'h6F; #100;
A = 8'hA5; B = 8'h70; #100;
A = 8'hA5; B = 8'h71; #100;
A = 8'hA5; B = 8'h72; #100;
A = 8'hA5; B = 8'h73; #100;
A = 8'hA5; B = 8'h74; #100;
A = 8'hA5; B = 8'h75; #100;
A = 8'hA5; B = 8'h76; #100;
A = 8'hA5; B = 8'h77; #100;
A = 8'hA5; B = 8'h78; #100;
A = 8'hA5; B = 8'h79; #100;
A = 8'hA5; B = 8'h7A; #100;
A = 8'hA5; B = 8'h7B; #100;
A = 8'hA5; B = 8'h7C; #100;
A = 8'hA5; B = 8'h7D; #100;
A = 8'hA5; B = 8'h7E; #100;
A = 8'hA5; B = 8'h7F; #100;
A = 8'hA5; B = 8'h80; #100;
A = 8'hA5; B = 8'h81; #100;
A = 8'hA5; B = 8'h82; #100;
A = 8'hA5; B = 8'h83; #100;
A = 8'hA5; B = 8'h84; #100;
A = 8'hA5; B = 8'h85; #100;
A = 8'hA5; B = 8'h86; #100;
A = 8'hA5; B = 8'h87; #100;
A = 8'hA5; B = 8'h88; #100;
A = 8'hA5; B = 8'h89; #100;
A = 8'hA5; B = 8'h8A; #100;
A = 8'hA5; B = 8'h8B; #100;
A = 8'hA5; B = 8'h8C; #100;
A = 8'hA5; B = 8'h8D; #100;
A = 8'hA5; B = 8'h8E; #100;
A = 8'hA5; B = 8'h8F; #100;
A = 8'hA5; B = 8'h90; #100;
A = 8'hA5; B = 8'h91; #100;
A = 8'hA5; B = 8'h92; #100;
A = 8'hA5; B = 8'h93; #100;
A = 8'hA5; B = 8'h94; #100;
A = 8'hA5; B = 8'h95; #100;
A = 8'hA5; B = 8'h96; #100;
A = 8'hA5; B = 8'h97; #100;
A = 8'hA5; B = 8'h98; #100;
A = 8'hA5; B = 8'h99; #100;
A = 8'hA5; B = 8'h9A; #100;
A = 8'hA5; B = 8'h9B; #100;
A = 8'hA5; B = 8'h9C; #100;
A = 8'hA5; B = 8'h9D; #100;
A = 8'hA5; B = 8'h9E; #100;
A = 8'hA5; B = 8'h9F; #100;
A = 8'hA5; B = 8'hA0; #100;
A = 8'hA5; B = 8'hA1; #100;
A = 8'hA5; B = 8'hA2; #100;
A = 8'hA5; B = 8'hA3; #100;
A = 8'hA5; B = 8'hA4; #100;
A = 8'hA5; B = 8'hA5; #100;
A = 8'hA5; B = 8'hA6; #100;
A = 8'hA5; B = 8'hA7; #100;
A = 8'hA5; B = 8'hA8; #100;
A = 8'hA5; B = 8'hA9; #100;
A = 8'hA5; B = 8'hAA; #100;
A = 8'hA5; B = 8'hAB; #100;
A = 8'hA5; B = 8'hAC; #100;
A = 8'hA5; B = 8'hAD; #100;
A = 8'hA5; B = 8'hAE; #100;
A = 8'hA5; B = 8'hAF; #100;
A = 8'hA5; B = 8'hB0; #100;
A = 8'hA5; B = 8'hB1; #100;
A = 8'hA5; B = 8'hB2; #100;
A = 8'hA5; B = 8'hB3; #100;
A = 8'hA5; B = 8'hB4; #100;
A = 8'hA5; B = 8'hB5; #100;
A = 8'hA5; B = 8'hB6; #100;
A = 8'hA5; B = 8'hB7; #100;
A = 8'hA5; B = 8'hB8; #100;
A = 8'hA5; B = 8'hB9; #100;
A = 8'hA5; B = 8'hBA; #100;
A = 8'hA5; B = 8'hBB; #100;
A = 8'hA5; B = 8'hBC; #100;
A = 8'hA5; B = 8'hBD; #100;
A = 8'hA5; B = 8'hBE; #100;
A = 8'hA5; B = 8'hBF; #100;
A = 8'hA5; B = 8'hC0; #100;
A = 8'hA5; B = 8'hC1; #100;
A = 8'hA5; B = 8'hC2; #100;
A = 8'hA5; B = 8'hC3; #100;
A = 8'hA5; B = 8'hC4; #100;
A = 8'hA5; B = 8'hC5; #100;
A = 8'hA5; B = 8'hC6; #100;
A = 8'hA5; B = 8'hC7; #100;
A = 8'hA5; B = 8'hC8; #100;
A = 8'hA5; B = 8'hC9; #100;
A = 8'hA5; B = 8'hCA; #100;
A = 8'hA5; B = 8'hCB; #100;
A = 8'hA5; B = 8'hCC; #100;
A = 8'hA5; B = 8'hCD; #100;
A = 8'hA5; B = 8'hCE; #100;
A = 8'hA5; B = 8'hCF; #100;
A = 8'hA5; B = 8'hD0; #100;
A = 8'hA5; B = 8'hD1; #100;
A = 8'hA5; B = 8'hD2; #100;
A = 8'hA5; B = 8'hD3; #100;
A = 8'hA5; B = 8'hD4; #100;
A = 8'hA5; B = 8'hD5; #100;
A = 8'hA5; B = 8'hD6; #100;
A = 8'hA5; B = 8'hD7; #100;
A = 8'hA5; B = 8'hD8; #100;
A = 8'hA5; B = 8'hD9; #100;
A = 8'hA5; B = 8'hDA; #100;
A = 8'hA5; B = 8'hDB; #100;
A = 8'hA5; B = 8'hDC; #100;
A = 8'hA5; B = 8'hDD; #100;
A = 8'hA5; B = 8'hDE; #100;
A = 8'hA5; B = 8'hDF; #100;
A = 8'hA5; B = 8'hE0; #100;
A = 8'hA5; B = 8'hE1; #100;
A = 8'hA5; B = 8'hE2; #100;
A = 8'hA5; B = 8'hE3; #100;
A = 8'hA5; B = 8'hE4; #100;
A = 8'hA5; B = 8'hE5; #100;
A = 8'hA5; B = 8'hE6; #100;
A = 8'hA5; B = 8'hE7; #100;
A = 8'hA5; B = 8'hE8; #100;
A = 8'hA5; B = 8'hE9; #100;
A = 8'hA5; B = 8'hEA; #100;
A = 8'hA5; B = 8'hEB; #100;
A = 8'hA5; B = 8'hEC; #100;
A = 8'hA5; B = 8'hED; #100;
A = 8'hA5; B = 8'hEE; #100;
A = 8'hA5; B = 8'hEF; #100;
A = 8'hA5; B = 8'hF0; #100;
A = 8'hA5; B = 8'hF1; #100;
A = 8'hA5; B = 8'hF2; #100;
A = 8'hA5; B = 8'hF3; #100;
A = 8'hA5; B = 8'hF4; #100;
A = 8'hA5; B = 8'hF5; #100;
A = 8'hA5; B = 8'hF6; #100;
A = 8'hA5; B = 8'hF7; #100;
A = 8'hA5; B = 8'hF8; #100;
A = 8'hA5; B = 8'hF9; #100;
A = 8'hA5; B = 8'hFA; #100;
A = 8'hA5; B = 8'hFB; #100;
A = 8'hA5; B = 8'hFC; #100;
A = 8'hA5; B = 8'hFD; #100;
A = 8'hA5; B = 8'hFE; #100;
A = 8'hA5; B = 8'hFF; #100;
A = 8'hA6; B = 8'h0; #100;
A = 8'hA6; B = 8'h1; #100;
A = 8'hA6; B = 8'h2; #100;
A = 8'hA6; B = 8'h3; #100;
A = 8'hA6; B = 8'h4; #100;
A = 8'hA6; B = 8'h5; #100;
A = 8'hA6; B = 8'h6; #100;
A = 8'hA6; B = 8'h7; #100;
A = 8'hA6; B = 8'h8; #100;
A = 8'hA6; B = 8'h9; #100;
A = 8'hA6; B = 8'hA; #100;
A = 8'hA6; B = 8'hB; #100;
A = 8'hA6; B = 8'hC; #100;
A = 8'hA6; B = 8'hD; #100;
A = 8'hA6; B = 8'hE; #100;
A = 8'hA6; B = 8'hF; #100;
A = 8'hA6; B = 8'h10; #100;
A = 8'hA6; B = 8'h11; #100;
A = 8'hA6; B = 8'h12; #100;
A = 8'hA6; B = 8'h13; #100;
A = 8'hA6; B = 8'h14; #100;
A = 8'hA6; B = 8'h15; #100;
A = 8'hA6; B = 8'h16; #100;
A = 8'hA6; B = 8'h17; #100;
A = 8'hA6; B = 8'h18; #100;
A = 8'hA6; B = 8'h19; #100;
A = 8'hA6; B = 8'h1A; #100;
A = 8'hA6; B = 8'h1B; #100;
A = 8'hA6; B = 8'h1C; #100;
A = 8'hA6; B = 8'h1D; #100;
A = 8'hA6; B = 8'h1E; #100;
A = 8'hA6; B = 8'h1F; #100;
A = 8'hA6; B = 8'h20; #100;
A = 8'hA6; B = 8'h21; #100;
A = 8'hA6; B = 8'h22; #100;
A = 8'hA6; B = 8'h23; #100;
A = 8'hA6; B = 8'h24; #100;
A = 8'hA6; B = 8'h25; #100;
A = 8'hA6; B = 8'h26; #100;
A = 8'hA6; B = 8'h27; #100;
A = 8'hA6; B = 8'h28; #100;
A = 8'hA6; B = 8'h29; #100;
A = 8'hA6; B = 8'h2A; #100;
A = 8'hA6; B = 8'h2B; #100;
A = 8'hA6; B = 8'h2C; #100;
A = 8'hA6; B = 8'h2D; #100;
A = 8'hA6; B = 8'h2E; #100;
A = 8'hA6; B = 8'h2F; #100;
A = 8'hA6; B = 8'h30; #100;
A = 8'hA6; B = 8'h31; #100;
A = 8'hA6; B = 8'h32; #100;
A = 8'hA6; B = 8'h33; #100;
A = 8'hA6; B = 8'h34; #100;
A = 8'hA6; B = 8'h35; #100;
A = 8'hA6; B = 8'h36; #100;
A = 8'hA6; B = 8'h37; #100;
A = 8'hA6; B = 8'h38; #100;
A = 8'hA6; B = 8'h39; #100;
A = 8'hA6; B = 8'h3A; #100;
A = 8'hA6; B = 8'h3B; #100;
A = 8'hA6; B = 8'h3C; #100;
A = 8'hA6; B = 8'h3D; #100;
A = 8'hA6; B = 8'h3E; #100;
A = 8'hA6; B = 8'h3F; #100;
A = 8'hA6; B = 8'h40; #100;
A = 8'hA6; B = 8'h41; #100;
A = 8'hA6; B = 8'h42; #100;
A = 8'hA6; B = 8'h43; #100;
A = 8'hA6; B = 8'h44; #100;
A = 8'hA6; B = 8'h45; #100;
A = 8'hA6; B = 8'h46; #100;
A = 8'hA6; B = 8'h47; #100;
A = 8'hA6; B = 8'h48; #100;
A = 8'hA6; B = 8'h49; #100;
A = 8'hA6; B = 8'h4A; #100;
A = 8'hA6; B = 8'h4B; #100;
A = 8'hA6; B = 8'h4C; #100;
A = 8'hA6; B = 8'h4D; #100;
A = 8'hA6; B = 8'h4E; #100;
A = 8'hA6; B = 8'h4F; #100;
A = 8'hA6; B = 8'h50; #100;
A = 8'hA6; B = 8'h51; #100;
A = 8'hA6; B = 8'h52; #100;
A = 8'hA6; B = 8'h53; #100;
A = 8'hA6; B = 8'h54; #100;
A = 8'hA6; B = 8'h55; #100;
A = 8'hA6; B = 8'h56; #100;
A = 8'hA6; B = 8'h57; #100;
A = 8'hA6; B = 8'h58; #100;
A = 8'hA6; B = 8'h59; #100;
A = 8'hA6; B = 8'h5A; #100;
A = 8'hA6; B = 8'h5B; #100;
A = 8'hA6; B = 8'h5C; #100;
A = 8'hA6; B = 8'h5D; #100;
A = 8'hA6; B = 8'h5E; #100;
A = 8'hA6; B = 8'h5F; #100;
A = 8'hA6; B = 8'h60; #100;
A = 8'hA6; B = 8'h61; #100;
A = 8'hA6; B = 8'h62; #100;
A = 8'hA6; B = 8'h63; #100;
A = 8'hA6; B = 8'h64; #100;
A = 8'hA6; B = 8'h65; #100;
A = 8'hA6; B = 8'h66; #100;
A = 8'hA6; B = 8'h67; #100;
A = 8'hA6; B = 8'h68; #100;
A = 8'hA6; B = 8'h69; #100;
A = 8'hA6; B = 8'h6A; #100;
A = 8'hA6; B = 8'h6B; #100;
A = 8'hA6; B = 8'h6C; #100;
A = 8'hA6; B = 8'h6D; #100;
A = 8'hA6; B = 8'h6E; #100;
A = 8'hA6; B = 8'h6F; #100;
A = 8'hA6; B = 8'h70; #100;
A = 8'hA6; B = 8'h71; #100;
A = 8'hA6; B = 8'h72; #100;
A = 8'hA6; B = 8'h73; #100;
A = 8'hA6; B = 8'h74; #100;
A = 8'hA6; B = 8'h75; #100;
A = 8'hA6; B = 8'h76; #100;
A = 8'hA6; B = 8'h77; #100;
A = 8'hA6; B = 8'h78; #100;
A = 8'hA6; B = 8'h79; #100;
A = 8'hA6; B = 8'h7A; #100;
A = 8'hA6; B = 8'h7B; #100;
A = 8'hA6; B = 8'h7C; #100;
A = 8'hA6; B = 8'h7D; #100;
A = 8'hA6; B = 8'h7E; #100;
A = 8'hA6; B = 8'h7F; #100;
A = 8'hA6; B = 8'h80; #100;
A = 8'hA6; B = 8'h81; #100;
A = 8'hA6; B = 8'h82; #100;
A = 8'hA6; B = 8'h83; #100;
A = 8'hA6; B = 8'h84; #100;
A = 8'hA6; B = 8'h85; #100;
A = 8'hA6; B = 8'h86; #100;
A = 8'hA6; B = 8'h87; #100;
A = 8'hA6; B = 8'h88; #100;
A = 8'hA6; B = 8'h89; #100;
A = 8'hA6; B = 8'h8A; #100;
A = 8'hA6; B = 8'h8B; #100;
A = 8'hA6; B = 8'h8C; #100;
A = 8'hA6; B = 8'h8D; #100;
A = 8'hA6; B = 8'h8E; #100;
A = 8'hA6; B = 8'h8F; #100;
A = 8'hA6; B = 8'h90; #100;
A = 8'hA6; B = 8'h91; #100;
A = 8'hA6; B = 8'h92; #100;
A = 8'hA6; B = 8'h93; #100;
A = 8'hA6; B = 8'h94; #100;
A = 8'hA6; B = 8'h95; #100;
A = 8'hA6; B = 8'h96; #100;
A = 8'hA6; B = 8'h97; #100;
A = 8'hA6; B = 8'h98; #100;
A = 8'hA6; B = 8'h99; #100;
A = 8'hA6; B = 8'h9A; #100;
A = 8'hA6; B = 8'h9B; #100;
A = 8'hA6; B = 8'h9C; #100;
A = 8'hA6; B = 8'h9D; #100;
A = 8'hA6; B = 8'h9E; #100;
A = 8'hA6; B = 8'h9F; #100;
A = 8'hA6; B = 8'hA0; #100;
A = 8'hA6; B = 8'hA1; #100;
A = 8'hA6; B = 8'hA2; #100;
A = 8'hA6; B = 8'hA3; #100;
A = 8'hA6; B = 8'hA4; #100;
A = 8'hA6; B = 8'hA5; #100;
A = 8'hA6; B = 8'hA6; #100;
A = 8'hA6; B = 8'hA7; #100;
A = 8'hA6; B = 8'hA8; #100;
A = 8'hA6; B = 8'hA9; #100;
A = 8'hA6; B = 8'hAA; #100;
A = 8'hA6; B = 8'hAB; #100;
A = 8'hA6; B = 8'hAC; #100;
A = 8'hA6; B = 8'hAD; #100;
A = 8'hA6; B = 8'hAE; #100;
A = 8'hA6; B = 8'hAF; #100;
A = 8'hA6; B = 8'hB0; #100;
A = 8'hA6; B = 8'hB1; #100;
A = 8'hA6; B = 8'hB2; #100;
A = 8'hA6; B = 8'hB3; #100;
A = 8'hA6; B = 8'hB4; #100;
A = 8'hA6; B = 8'hB5; #100;
A = 8'hA6; B = 8'hB6; #100;
A = 8'hA6; B = 8'hB7; #100;
A = 8'hA6; B = 8'hB8; #100;
A = 8'hA6; B = 8'hB9; #100;
A = 8'hA6; B = 8'hBA; #100;
A = 8'hA6; B = 8'hBB; #100;
A = 8'hA6; B = 8'hBC; #100;
A = 8'hA6; B = 8'hBD; #100;
A = 8'hA6; B = 8'hBE; #100;
A = 8'hA6; B = 8'hBF; #100;
A = 8'hA6; B = 8'hC0; #100;
A = 8'hA6; B = 8'hC1; #100;
A = 8'hA6; B = 8'hC2; #100;
A = 8'hA6; B = 8'hC3; #100;
A = 8'hA6; B = 8'hC4; #100;
A = 8'hA6; B = 8'hC5; #100;
A = 8'hA6; B = 8'hC6; #100;
A = 8'hA6; B = 8'hC7; #100;
A = 8'hA6; B = 8'hC8; #100;
A = 8'hA6; B = 8'hC9; #100;
A = 8'hA6; B = 8'hCA; #100;
A = 8'hA6; B = 8'hCB; #100;
A = 8'hA6; B = 8'hCC; #100;
A = 8'hA6; B = 8'hCD; #100;
A = 8'hA6; B = 8'hCE; #100;
A = 8'hA6; B = 8'hCF; #100;
A = 8'hA6; B = 8'hD0; #100;
A = 8'hA6; B = 8'hD1; #100;
A = 8'hA6; B = 8'hD2; #100;
A = 8'hA6; B = 8'hD3; #100;
A = 8'hA6; B = 8'hD4; #100;
A = 8'hA6; B = 8'hD5; #100;
A = 8'hA6; B = 8'hD6; #100;
A = 8'hA6; B = 8'hD7; #100;
A = 8'hA6; B = 8'hD8; #100;
A = 8'hA6; B = 8'hD9; #100;
A = 8'hA6; B = 8'hDA; #100;
A = 8'hA6; B = 8'hDB; #100;
A = 8'hA6; B = 8'hDC; #100;
A = 8'hA6; B = 8'hDD; #100;
A = 8'hA6; B = 8'hDE; #100;
A = 8'hA6; B = 8'hDF; #100;
A = 8'hA6; B = 8'hE0; #100;
A = 8'hA6; B = 8'hE1; #100;
A = 8'hA6; B = 8'hE2; #100;
A = 8'hA6; B = 8'hE3; #100;
A = 8'hA6; B = 8'hE4; #100;
A = 8'hA6; B = 8'hE5; #100;
A = 8'hA6; B = 8'hE6; #100;
A = 8'hA6; B = 8'hE7; #100;
A = 8'hA6; B = 8'hE8; #100;
A = 8'hA6; B = 8'hE9; #100;
A = 8'hA6; B = 8'hEA; #100;
A = 8'hA6; B = 8'hEB; #100;
A = 8'hA6; B = 8'hEC; #100;
A = 8'hA6; B = 8'hED; #100;
A = 8'hA6; B = 8'hEE; #100;
A = 8'hA6; B = 8'hEF; #100;
A = 8'hA6; B = 8'hF0; #100;
A = 8'hA6; B = 8'hF1; #100;
A = 8'hA6; B = 8'hF2; #100;
A = 8'hA6; B = 8'hF3; #100;
A = 8'hA6; B = 8'hF4; #100;
A = 8'hA6; B = 8'hF5; #100;
A = 8'hA6; B = 8'hF6; #100;
A = 8'hA6; B = 8'hF7; #100;
A = 8'hA6; B = 8'hF8; #100;
A = 8'hA6; B = 8'hF9; #100;
A = 8'hA6; B = 8'hFA; #100;
A = 8'hA6; B = 8'hFB; #100;
A = 8'hA6; B = 8'hFC; #100;
A = 8'hA6; B = 8'hFD; #100;
A = 8'hA6; B = 8'hFE; #100;
A = 8'hA6; B = 8'hFF; #100;
A = 8'hA7; B = 8'h0; #100;
A = 8'hA7; B = 8'h1; #100;
A = 8'hA7; B = 8'h2; #100;
A = 8'hA7; B = 8'h3; #100;
A = 8'hA7; B = 8'h4; #100;
A = 8'hA7; B = 8'h5; #100;
A = 8'hA7; B = 8'h6; #100;
A = 8'hA7; B = 8'h7; #100;
A = 8'hA7; B = 8'h8; #100;
A = 8'hA7; B = 8'h9; #100;
A = 8'hA7; B = 8'hA; #100;
A = 8'hA7; B = 8'hB; #100;
A = 8'hA7; B = 8'hC; #100;
A = 8'hA7; B = 8'hD; #100;
A = 8'hA7; B = 8'hE; #100;
A = 8'hA7; B = 8'hF; #100;
A = 8'hA7; B = 8'h10; #100;
A = 8'hA7; B = 8'h11; #100;
A = 8'hA7; B = 8'h12; #100;
A = 8'hA7; B = 8'h13; #100;
A = 8'hA7; B = 8'h14; #100;
A = 8'hA7; B = 8'h15; #100;
A = 8'hA7; B = 8'h16; #100;
A = 8'hA7; B = 8'h17; #100;
A = 8'hA7; B = 8'h18; #100;
A = 8'hA7; B = 8'h19; #100;
A = 8'hA7; B = 8'h1A; #100;
A = 8'hA7; B = 8'h1B; #100;
A = 8'hA7; B = 8'h1C; #100;
A = 8'hA7; B = 8'h1D; #100;
A = 8'hA7; B = 8'h1E; #100;
A = 8'hA7; B = 8'h1F; #100;
A = 8'hA7; B = 8'h20; #100;
A = 8'hA7; B = 8'h21; #100;
A = 8'hA7; B = 8'h22; #100;
A = 8'hA7; B = 8'h23; #100;
A = 8'hA7; B = 8'h24; #100;
A = 8'hA7; B = 8'h25; #100;
A = 8'hA7; B = 8'h26; #100;
A = 8'hA7; B = 8'h27; #100;
A = 8'hA7; B = 8'h28; #100;
A = 8'hA7; B = 8'h29; #100;
A = 8'hA7; B = 8'h2A; #100;
A = 8'hA7; B = 8'h2B; #100;
A = 8'hA7; B = 8'h2C; #100;
A = 8'hA7; B = 8'h2D; #100;
A = 8'hA7; B = 8'h2E; #100;
A = 8'hA7; B = 8'h2F; #100;
A = 8'hA7; B = 8'h30; #100;
A = 8'hA7; B = 8'h31; #100;
A = 8'hA7; B = 8'h32; #100;
A = 8'hA7; B = 8'h33; #100;
A = 8'hA7; B = 8'h34; #100;
A = 8'hA7; B = 8'h35; #100;
A = 8'hA7; B = 8'h36; #100;
A = 8'hA7; B = 8'h37; #100;
A = 8'hA7; B = 8'h38; #100;
A = 8'hA7; B = 8'h39; #100;
A = 8'hA7; B = 8'h3A; #100;
A = 8'hA7; B = 8'h3B; #100;
A = 8'hA7; B = 8'h3C; #100;
A = 8'hA7; B = 8'h3D; #100;
A = 8'hA7; B = 8'h3E; #100;
A = 8'hA7; B = 8'h3F; #100;
A = 8'hA7; B = 8'h40; #100;
A = 8'hA7; B = 8'h41; #100;
A = 8'hA7; B = 8'h42; #100;
A = 8'hA7; B = 8'h43; #100;
A = 8'hA7; B = 8'h44; #100;
A = 8'hA7; B = 8'h45; #100;
A = 8'hA7; B = 8'h46; #100;
A = 8'hA7; B = 8'h47; #100;
A = 8'hA7; B = 8'h48; #100;
A = 8'hA7; B = 8'h49; #100;
A = 8'hA7; B = 8'h4A; #100;
A = 8'hA7; B = 8'h4B; #100;
A = 8'hA7; B = 8'h4C; #100;
A = 8'hA7; B = 8'h4D; #100;
A = 8'hA7; B = 8'h4E; #100;
A = 8'hA7; B = 8'h4F; #100;
A = 8'hA7; B = 8'h50; #100;
A = 8'hA7; B = 8'h51; #100;
A = 8'hA7; B = 8'h52; #100;
A = 8'hA7; B = 8'h53; #100;
A = 8'hA7; B = 8'h54; #100;
A = 8'hA7; B = 8'h55; #100;
A = 8'hA7; B = 8'h56; #100;
A = 8'hA7; B = 8'h57; #100;
A = 8'hA7; B = 8'h58; #100;
A = 8'hA7; B = 8'h59; #100;
A = 8'hA7; B = 8'h5A; #100;
A = 8'hA7; B = 8'h5B; #100;
A = 8'hA7; B = 8'h5C; #100;
A = 8'hA7; B = 8'h5D; #100;
A = 8'hA7; B = 8'h5E; #100;
A = 8'hA7; B = 8'h5F; #100;
A = 8'hA7; B = 8'h60; #100;
A = 8'hA7; B = 8'h61; #100;
A = 8'hA7; B = 8'h62; #100;
A = 8'hA7; B = 8'h63; #100;
A = 8'hA7; B = 8'h64; #100;
A = 8'hA7; B = 8'h65; #100;
A = 8'hA7; B = 8'h66; #100;
A = 8'hA7; B = 8'h67; #100;
A = 8'hA7; B = 8'h68; #100;
A = 8'hA7; B = 8'h69; #100;
A = 8'hA7; B = 8'h6A; #100;
A = 8'hA7; B = 8'h6B; #100;
A = 8'hA7; B = 8'h6C; #100;
A = 8'hA7; B = 8'h6D; #100;
A = 8'hA7; B = 8'h6E; #100;
A = 8'hA7; B = 8'h6F; #100;
A = 8'hA7; B = 8'h70; #100;
A = 8'hA7; B = 8'h71; #100;
A = 8'hA7; B = 8'h72; #100;
A = 8'hA7; B = 8'h73; #100;
A = 8'hA7; B = 8'h74; #100;
A = 8'hA7; B = 8'h75; #100;
A = 8'hA7; B = 8'h76; #100;
A = 8'hA7; B = 8'h77; #100;
A = 8'hA7; B = 8'h78; #100;
A = 8'hA7; B = 8'h79; #100;
A = 8'hA7; B = 8'h7A; #100;
A = 8'hA7; B = 8'h7B; #100;
A = 8'hA7; B = 8'h7C; #100;
A = 8'hA7; B = 8'h7D; #100;
A = 8'hA7; B = 8'h7E; #100;
A = 8'hA7; B = 8'h7F; #100;
A = 8'hA7; B = 8'h80; #100;
A = 8'hA7; B = 8'h81; #100;
A = 8'hA7; B = 8'h82; #100;
A = 8'hA7; B = 8'h83; #100;
A = 8'hA7; B = 8'h84; #100;
A = 8'hA7; B = 8'h85; #100;
A = 8'hA7; B = 8'h86; #100;
A = 8'hA7; B = 8'h87; #100;
A = 8'hA7; B = 8'h88; #100;
A = 8'hA7; B = 8'h89; #100;
A = 8'hA7; B = 8'h8A; #100;
A = 8'hA7; B = 8'h8B; #100;
A = 8'hA7; B = 8'h8C; #100;
A = 8'hA7; B = 8'h8D; #100;
A = 8'hA7; B = 8'h8E; #100;
A = 8'hA7; B = 8'h8F; #100;
A = 8'hA7; B = 8'h90; #100;
A = 8'hA7; B = 8'h91; #100;
A = 8'hA7; B = 8'h92; #100;
A = 8'hA7; B = 8'h93; #100;
A = 8'hA7; B = 8'h94; #100;
A = 8'hA7; B = 8'h95; #100;
A = 8'hA7; B = 8'h96; #100;
A = 8'hA7; B = 8'h97; #100;
A = 8'hA7; B = 8'h98; #100;
A = 8'hA7; B = 8'h99; #100;
A = 8'hA7; B = 8'h9A; #100;
A = 8'hA7; B = 8'h9B; #100;
A = 8'hA7; B = 8'h9C; #100;
A = 8'hA7; B = 8'h9D; #100;
A = 8'hA7; B = 8'h9E; #100;
A = 8'hA7; B = 8'h9F; #100;
A = 8'hA7; B = 8'hA0; #100;
A = 8'hA7; B = 8'hA1; #100;
A = 8'hA7; B = 8'hA2; #100;
A = 8'hA7; B = 8'hA3; #100;
A = 8'hA7; B = 8'hA4; #100;
A = 8'hA7; B = 8'hA5; #100;
A = 8'hA7; B = 8'hA6; #100;
A = 8'hA7; B = 8'hA7; #100;
A = 8'hA7; B = 8'hA8; #100;
A = 8'hA7; B = 8'hA9; #100;
A = 8'hA7; B = 8'hAA; #100;
A = 8'hA7; B = 8'hAB; #100;
A = 8'hA7; B = 8'hAC; #100;
A = 8'hA7; B = 8'hAD; #100;
A = 8'hA7; B = 8'hAE; #100;
A = 8'hA7; B = 8'hAF; #100;
A = 8'hA7; B = 8'hB0; #100;
A = 8'hA7; B = 8'hB1; #100;
A = 8'hA7; B = 8'hB2; #100;
A = 8'hA7; B = 8'hB3; #100;
A = 8'hA7; B = 8'hB4; #100;
A = 8'hA7; B = 8'hB5; #100;
A = 8'hA7; B = 8'hB6; #100;
A = 8'hA7; B = 8'hB7; #100;
A = 8'hA7; B = 8'hB8; #100;
A = 8'hA7; B = 8'hB9; #100;
A = 8'hA7; B = 8'hBA; #100;
A = 8'hA7; B = 8'hBB; #100;
A = 8'hA7; B = 8'hBC; #100;
A = 8'hA7; B = 8'hBD; #100;
A = 8'hA7; B = 8'hBE; #100;
A = 8'hA7; B = 8'hBF; #100;
A = 8'hA7; B = 8'hC0; #100;
A = 8'hA7; B = 8'hC1; #100;
A = 8'hA7; B = 8'hC2; #100;
A = 8'hA7; B = 8'hC3; #100;
A = 8'hA7; B = 8'hC4; #100;
A = 8'hA7; B = 8'hC5; #100;
A = 8'hA7; B = 8'hC6; #100;
A = 8'hA7; B = 8'hC7; #100;
A = 8'hA7; B = 8'hC8; #100;
A = 8'hA7; B = 8'hC9; #100;
A = 8'hA7; B = 8'hCA; #100;
A = 8'hA7; B = 8'hCB; #100;
A = 8'hA7; B = 8'hCC; #100;
A = 8'hA7; B = 8'hCD; #100;
A = 8'hA7; B = 8'hCE; #100;
A = 8'hA7; B = 8'hCF; #100;
A = 8'hA7; B = 8'hD0; #100;
A = 8'hA7; B = 8'hD1; #100;
A = 8'hA7; B = 8'hD2; #100;
A = 8'hA7; B = 8'hD3; #100;
A = 8'hA7; B = 8'hD4; #100;
A = 8'hA7; B = 8'hD5; #100;
A = 8'hA7; B = 8'hD6; #100;
A = 8'hA7; B = 8'hD7; #100;
A = 8'hA7; B = 8'hD8; #100;
A = 8'hA7; B = 8'hD9; #100;
A = 8'hA7; B = 8'hDA; #100;
A = 8'hA7; B = 8'hDB; #100;
A = 8'hA7; B = 8'hDC; #100;
A = 8'hA7; B = 8'hDD; #100;
A = 8'hA7; B = 8'hDE; #100;
A = 8'hA7; B = 8'hDF; #100;
A = 8'hA7; B = 8'hE0; #100;
A = 8'hA7; B = 8'hE1; #100;
A = 8'hA7; B = 8'hE2; #100;
A = 8'hA7; B = 8'hE3; #100;
A = 8'hA7; B = 8'hE4; #100;
A = 8'hA7; B = 8'hE5; #100;
A = 8'hA7; B = 8'hE6; #100;
A = 8'hA7; B = 8'hE7; #100;
A = 8'hA7; B = 8'hE8; #100;
A = 8'hA7; B = 8'hE9; #100;
A = 8'hA7; B = 8'hEA; #100;
A = 8'hA7; B = 8'hEB; #100;
A = 8'hA7; B = 8'hEC; #100;
A = 8'hA7; B = 8'hED; #100;
A = 8'hA7; B = 8'hEE; #100;
A = 8'hA7; B = 8'hEF; #100;
A = 8'hA7; B = 8'hF0; #100;
A = 8'hA7; B = 8'hF1; #100;
A = 8'hA7; B = 8'hF2; #100;
A = 8'hA7; B = 8'hF3; #100;
A = 8'hA7; B = 8'hF4; #100;
A = 8'hA7; B = 8'hF5; #100;
A = 8'hA7; B = 8'hF6; #100;
A = 8'hA7; B = 8'hF7; #100;
A = 8'hA7; B = 8'hF8; #100;
A = 8'hA7; B = 8'hF9; #100;
A = 8'hA7; B = 8'hFA; #100;
A = 8'hA7; B = 8'hFB; #100;
A = 8'hA7; B = 8'hFC; #100;
A = 8'hA7; B = 8'hFD; #100;
A = 8'hA7; B = 8'hFE; #100;
A = 8'hA7; B = 8'hFF; #100;
A = 8'hA8; B = 8'h0; #100;
A = 8'hA8; B = 8'h1; #100;
A = 8'hA8; B = 8'h2; #100;
A = 8'hA8; B = 8'h3; #100;
A = 8'hA8; B = 8'h4; #100;
A = 8'hA8; B = 8'h5; #100;
A = 8'hA8; B = 8'h6; #100;
A = 8'hA8; B = 8'h7; #100;
A = 8'hA8; B = 8'h8; #100;
A = 8'hA8; B = 8'h9; #100;
A = 8'hA8; B = 8'hA; #100;
A = 8'hA8; B = 8'hB; #100;
A = 8'hA8; B = 8'hC; #100;
A = 8'hA8; B = 8'hD; #100;
A = 8'hA8; B = 8'hE; #100;
A = 8'hA8; B = 8'hF; #100;
A = 8'hA8; B = 8'h10; #100;
A = 8'hA8; B = 8'h11; #100;
A = 8'hA8; B = 8'h12; #100;
A = 8'hA8; B = 8'h13; #100;
A = 8'hA8; B = 8'h14; #100;
A = 8'hA8; B = 8'h15; #100;
A = 8'hA8; B = 8'h16; #100;
A = 8'hA8; B = 8'h17; #100;
A = 8'hA8; B = 8'h18; #100;
A = 8'hA8; B = 8'h19; #100;
A = 8'hA8; B = 8'h1A; #100;
A = 8'hA8; B = 8'h1B; #100;
A = 8'hA8; B = 8'h1C; #100;
A = 8'hA8; B = 8'h1D; #100;
A = 8'hA8; B = 8'h1E; #100;
A = 8'hA8; B = 8'h1F; #100;
A = 8'hA8; B = 8'h20; #100;
A = 8'hA8; B = 8'h21; #100;
A = 8'hA8; B = 8'h22; #100;
A = 8'hA8; B = 8'h23; #100;
A = 8'hA8; B = 8'h24; #100;
A = 8'hA8; B = 8'h25; #100;
A = 8'hA8; B = 8'h26; #100;
A = 8'hA8; B = 8'h27; #100;
A = 8'hA8; B = 8'h28; #100;
A = 8'hA8; B = 8'h29; #100;
A = 8'hA8; B = 8'h2A; #100;
A = 8'hA8; B = 8'h2B; #100;
A = 8'hA8; B = 8'h2C; #100;
A = 8'hA8; B = 8'h2D; #100;
A = 8'hA8; B = 8'h2E; #100;
A = 8'hA8; B = 8'h2F; #100;
A = 8'hA8; B = 8'h30; #100;
A = 8'hA8; B = 8'h31; #100;
A = 8'hA8; B = 8'h32; #100;
A = 8'hA8; B = 8'h33; #100;
A = 8'hA8; B = 8'h34; #100;
A = 8'hA8; B = 8'h35; #100;
A = 8'hA8; B = 8'h36; #100;
A = 8'hA8; B = 8'h37; #100;
A = 8'hA8; B = 8'h38; #100;
A = 8'hA8; B = 8'h39; #100;
A = 8'hA8; B = 8'h3A; #100;
A = 8'hA8; B = 8'h3B; #100;
A = 8'hA8; B = 8'h3C; #100;
A = 8'hA8; B = 8'h3D; #100;
A = 8'hA8; B = 8'h3E; #100;
A = 8'hA8; B = 8'h3F; #100;
A = 8'hA8; B = 8'h40; #100;
A = 8'hA8; B = 8'h41; #100;
A = 8'hA8; B = 8'h42; #100;
A = 8'hA8; B = 8'h43; #100;
A = 8'hA8; B = 8'h44; #100;
A = 8'hA8; B = 8'h45; #100;
A = 8'hA8; B = 8'h46; #100;
A = 8'hA8; B = 8'h47; #100;
A = 8'hA8; B = 8'h48; #100;
A = 8'hA8; B = 8'h49; #100;
A = 8'hA8; B = 8'h4A; #100;
A = 8'hA8; B = 8'h4B; #100;
A = 8'hA8; B = 8'h4C; #100;
A = 8'hA8; B = 8'h4D; #100;
A = 8'hA8; B = 8'h4E; #100;
A = 8'hA8; B = 8'h4F; #100;
A = 8'hA8; B = 8'h50; #100;
A = 8'hA8; B = 8'h51; #100;
A = 8'hA8; B = 8'h52; #100;
A = 8'hA8; B = 8'h53; #100;
A = 8'hA8; B = 8'h54; #100;
A = 8'hA8; B = 8'h55; #100;
A = 8'hA8; B = 8'h56; #100;
A = 8'hA8; B = 8'h57; #100;
A = 8'hA8; B = 8'h58; #100;
A = 8'hA8; B = 8'h59; #100;
A = 8'hA8; B = 8'h5A; #100;
A = 8'hA8; B = 8'h5B; #100;
A = 8'hA8; B = 8'h5C; #100;
A = 8'hA8; B = 8'h5D; #100;
A = 8'hA8; B = 8'h5E; #100;
A = 8'hA8; B = 8'h5F; #100;
A = 8'hA8; B = 8'h60; #100;
A = 8'hA8; B = 8'h61; #100;
A = 8'hA8; B = 8'h62; #100;
A = 8'hA8; B = 8'h63; #100;
A = 8'hA8; B = 8'h64; #100;
A = 8'hA8; B = 8'h65; #100;
A = 8'hA8; B = 8'h66; #100;
A = 8'hA8; B = 8'h67; #100;
A = 8'hA8; B = 8'h68; #100;
A = 8'hA8; B = 8'h69; #100;
A = 8'hA8; B = 8'h6A; #100;
A = 8'hA8; B = 8'h6B; #100;
A = 8'hA8; B = 8'h6C; #100;
A = 8'hA8; B = 8'h6D; #100;
A = 8'hA8; B = 8'h6E; #100;
A = 8'hA8; B = 8'h6F; #100;
A = 8'hA8; B = 8'h70; #100;
A = 8'hA8; B = 8'h71; #100;
A = 8'hA8; B = 8'h72; #100;
A = 8'hA8; B = 8'h73; #100;
A = 8'hA8; B = 8'h74; #100;
A = 8'hA8; B = 8'h75; #100;
A = 8'hA8; B = 8'h76; #100;
A = 8'hA8; B = 8'h77; #100;
A = 8'hA8; B = 8'h78; #100;
A = 8'hA8; B = 8'h79; #100;
A = 8'hA8; B = 8'h7A; #100;
A = 8'hA8; B = 8'h7B; #100;
A = 8'hA8; B = 8'h7C; #100;
A = 8'hA8; B = 8'h7D; #100;
A = 8'hA8; B = 8'h7E; #100;
A = 8'hA8; B = 8'h7F; #100;
A = 8'hA8; B = 8'h80; #100;
A = 8'hA8; B = 8'h81; #100;
A = 8'hA8; B = 8'h82; #100;
A = 8'hA8; B = 8'h83; #100;
A = 8'hA8; B = 8'h84; #100;
A = 8'hA8; B = 8'h85; #100;
A = 8'hA8; B = 8'h86; #100;
A = 8'hA8; B = 8'h87; #100;
A = 8'hA8; B = 8'h88; #100;
A = 8'hA8; B = 8'h89; #100;
A = 8'hA8; B = 8'h8A; #100;
A = 8'hA8; B = 8'h8B; #100;
A = 8'hA8; B = 8'h8C; #100;
A = 8'hA8; B = 8'h8D; #100;
A = 8'hA8; B = 8'h8E; #100;
A = 8'hA8; B = 8'h8F; #100;
A = 8'hA8; B = 8'h90; #100;
A = 8'hA8; B = 8'h91; #100;
A = 8'hA8; B = 8'h92; #100;
A = 8'hA8; B = 8'h93; #100;
A = 8'hA8; B = 8'h94; #100;
A = 8'hA8; B = 8'h95; #100;
A = 8'hA8; B = 8'h96; #100;
A = 8'hA8; B = 8'h97; #100;
A = 8'hA8; B = 8'h98; #100;
A = 8'hA8; B = 8'h99; #100;
A = 8'hA8; B = 8'h9A; #100;
A = 8'hA8; B = 8'h9B; #100;
A = 8'hA8; B = 8'h9C; #100;
A = 8'hA8; B = 8'h9D; #100;
A = 8'hA8; B = 8'h9E; #100;
A = 8'hA8; B = 8'h9F; #100;
A = 8'hA8; B = 8'hA0; #100;
A = 8'hA8; B = 8'hA1; #100;
A = 8'hA8; B = 8'hA2; #100;
A = 8'hA8; B = 8'hA3; #100;
A = 8'hA8; B = 8'hA4; #100;
A = 8'hA8; B = 8'hA5; #100;
A = 8'hA8; B = 8'hA6; #100;
A = 8'hA8; B = 8'hA7; #100;
A = 8'hA8; B = 8'hA8; #100;
A = 8'hA8; B = 8'hA9; #100;
A = 8'hA8; B = 8'hAA; #100;
A = 8'hA8; B = 8'hAB; #100;
A = 8'hA8; B = 8'hAC; #100;
A = 8'hA8; B = 8'hAD; #100;
A = 8'hA8; B = 8'hAE; #100;
A = 8'hA8; B = 8'hAF; #100;
A = 8'hA8; B = 8'hB0; #100;
A = 8'hA8; B = 8'hB1; #100;
A = 8'hA8; B = 8'hB2; #100;
A = 8'hA8; B = 8'hB3; #100;
A = 8'hA8; B = 8'hB4; #100;
A = 8'hA8; B = 8'hB5; #100;
A = 8'hA8; B = 8'hB6; #100;
A = 8'hA8; B = 8'hB7; #100;
A = 8'hA8; B = 8'hB8; #100;
A = 8'hA8; B = 8'hB9; #100;
A = 8'hA8; B = 8'hBA; #100;
A = 8'hA8; B = 8'hBB; #100;
A = 8'hA8; B = 8'hBC; #100;
A = 8'hA8; B = 8'hBD; #100;
A = 8'hA8; B = 8'hBE; #100;
A = 8'hA8; B = 8'hBF; #100;
A = 8'hA8; B = 8'hC0; #100;
A = 8'hA8; B = 8'hC1; #100;
A = 8'hA8; B = 8'hC2; #100;
A = 8'hA8; B = 8'hC3; #100;
A = 8'hA8; B = 8'hC4; #100;
A = 8'hA8; B = 8'hC5; #100;
A = 8'hA8; B = 8'hC6; #100;
A = 8'hA8; B = 8'hC7; #100;
A = 8'hA8; B = 8'hC8; #100;
A = 8'hA8; B = 8'hC9; #100;
A = 8'hA8; B = 8'hCA; #100;
A = 8'hA8; B = 8'hCB; #100;
A = 8'hA8; B = 8'hCC; #100;
A = 8'hA8; B = 8'hCD; #100;
A = 8'hA8; B = 8'hCE; #100;
A = 8'hA8; B = 8'hCF; #100;
A = 8'hA8; B = 8'hD0; #100;
A = 8'hA8; B = 8'hD1; #100;
A = 8'hA8; B = 8'hD2; #100;
A = 8'hA8; B = 8'hD3; #100;
A = 8'hA8; B = 8'hD4; #100;
A = 8'hA8; B = 8'hD5; #100;
A = 8'hA8; B = 8'hD6; #100;
A = 8'hA8; B = 8'hD7; #100;
A = 8'hA8; B = 8'hD8; #100;
A = 8'hA8; B = 8'hD9; #100;
A = 8'hA8; B = 8'hDA; #100;
A = 8'hA8; B = 8'hDB; #100;
A = 8'hA8; B = 8'hDC; #100;
A = 8'hA8; B = 8'hDD; #100;
A = 8'hA8; B = 8'hDE; #100;
A = 8'hA8; B = 8'hDF; #100;
A = 8'hA8; B = 8'hE0; #100;
A = 8'hA8; B = 8'hE1; #100;
A = 8'hA8; B = 8'hE2; #100;
A = 8'hA8; B = 8'hE3; #100;
A = 8'hA8; B = 8'hE4; #100;
A = 8'hA8; B = 8'hE5; #100;
A = 8'hA8; B = 8'hE6; #100;
A = 8'hA8; B = 8'hE7; #100;
A = 8'hA8; B = 8'hE8; #100;
A = 8'hA8; B = 8'hE9; #100;
A = 8'hA8; B = 8'hEA; #100;
A = 8'hA8; B = 8'hEB; #100;
A = 8'hA8; B = 8'hEC; #100;
A = 8'hA8; B = 8'hED; #100;
A = 8'hA8; B = 8'hEE; #100;
A = 8'hA8; B = 8'hEF; #100;
A = 8'hA8; B = 8'hF0; #100;
A = 8'hA8; B = 8'hF1; #100;
A = 8'hA8; B = 8'hF2; #100;
A = 8'hA8; B = 8'hF3; #100;
A = 8'hA8; B = 8'hF4; #100;
A = 8'hA8; B = 8'hF5; #100;
A = 8'hA8; B = 8'hF6; #100;
A = 8'hA8; B = 8'hF7; #100;
A = 8'hA8; B = 8'hF8; #100;
A = 8'hA8; B = 8'hF9; #100;
A = 8'hA8; B = 8'hFA; #100;
A = 8'hA8; B = 8'hFB; #100;
A = 8'hA8; B = 8'hFC; #100;
A = 8'hA8; B = 8'hFD; #100;
A = 8'hA8; B = 8'hFE; #100;
A = 8'hA8; B = 8'hFF; #100;
A = 8'hA9; B = 8'h0; #100;
A = 8'hA9; B = 8'h1; #100;
A = 8'hA9; B = 8'h2; #100;
A = 8'hA9; B = 8'h3; #100;
A = 8'hA9; B = 8'h4; #100;
A = 8'hA9; B = 8'h5; #100;
A = 8'hA9; B = 8'h6; #100;
A = 8'hA9; B = 8'h7; #100;
A = 8'hA9; B = 8'h8; #100;
A = 8'hA9; B = 8'h9; #100;
A = 8'hA9; B = 8'hA; #100;
A = 8'hA9; B = 8'hB; #100;
A = 8'hA9; B = 8'hC; #100;
A = 8'hA9; B = 8'hD; #100;
A = 8'hA9; B = 8'hE; #100;
A = 8'hA9; B = 8'hF; #100;
A = 8'hA9; B = 8'h10; #100;
A = 8'hA9; B = 8'h11; #100;
A = 8'hA9; B = 8'h12; #100;
A = 8'hA9; B = 8'h13; #100;
A = 8'hA9; B = 8'h14; #100;
A = 8'hA9; B = 8'h15; #100;
A = 8'hA9; B = 8'h16; #100;
A = 8'hA9; B = 8'h17; #100;
A = 8'hA9; B = 8'h18; #100;
A = 8'hA9; B = 8'h19; #100;
A = 8'hA9; B = 8'h1A; #100;
A = 8'hA9; B = 8'h1B; #100;
A = 8'hA9; B = 8'h1C; #100;
A = 8'hA9; B = 8'h1D; #100;
A = 8'hA9; B = 8'h1E; #100;
A = 8'hA9; B = 8'h1F; #100;
A = 8'hA9; B = 8'h20; #100;
A = 8'hA9; B = 8'h21; #100;
A = 8'hA9; B = 8'h22; #100;
A = 8'hA9; B = 8'h23; #100;
A = 8'hA9; B = 8'h24; #100;
A = 8'hA9; B = 8'h25; #100;
A = 8'hA9; B = 8'h26; #100;
A = 8'hA9; B = 8'h27; #100;
A = 8'hA9; B = 8'h28; #100;
A = 8'hA9; B = 8'h29; #100;
A = 8'hA9; B = 8'h2A; #100;
A = 8'hA9; B = 8'h2B; #100;
A = 8'hA9; B = 8'h2C; #100;
A = 8'hA9; B = 8'h2D; #100;
A = 8'hA9; B = 8'h2E; #100;
A = 8'hA9; B = 8'h2F; #100;
A = 8'hA9; B = 8'h30; #100;
A = 8'hA9; B = 8'h31; #100;
A = 8'hA9; B = 8'h32; #100;
A = 8'hA9; B = 8'h33; #100;
A = 8'hA9; B = 8'h34; #100;
A = 8'hA9; B = 8'h35; #100;
A = 8'hA9; B = 8'h36; #100;
A = 8'hA9; B = 8'h37; #100;
A = 8'hA9; B = 8'h38; #100;
A = 8'hA9; B = 8'h39; #100;
A = 8'hA9; B = 8'h3A; #100;
A = 8'hA9; B = 8'h3B; #100;
A = 8'hA9; B = 8'h3C; #100;
A = 8'hA9; B = 8'h3D; #100;
A = 8'hA9; B = 8'h3E; #100;
A = 8'hA9; B = 8'h3F; #100;
A = 8'hA9; B = 8'h40; #100;
A = 8'hA9; B = 8'h41; #100;
A = 8'hA9; B = 8'h42; #100;
A = 8'hA9; B = 8'h43; #100;
A = 8'hA9; B = 8'h44; #100;
A = 8'hA9; B = 8'h45; #100;
A = 8'hA9; B = 8'h46; #100;
A = 8'hA9; B = 8'h47; #100;
A = 8'hA9; B = 8'h48; #100;
A = 8'hA9; B = 8'h49; #100;
A = 8'hA9; B = 8'h4A; #100;
A = 8'hA9; B = 8'h4B; #100;
A = 8'hA9; B = 8'h4C; #100;
A = 8'hA9; B = 8'h4D; #100;
A = 8'hA9; B = 8'h4E; #100;
A = 8'hA9; B = 8'h4F; #100;
A = 8'hA9; B = 8'h50; #100;
A = 8'hA9; B = 8'h51; #100;
A = 8'hA9; B = 8'h52; #100;
A = 8'hA9; B = 8'h53; #100;
A = 8'hA9; B = 8'h54; #100;
A = 8'hA9; B = 8'h55; #100;
A = 8'hA9; B = 8'h56; #100;
A = 8'hA9; B = 8'h57; #100;
A = 8'hA9; B = 8'h58; #100;
A = 8'hA9; B = 8'h59; #100;
A = 8'hA9; B = 8'h5A; #100;
A = 8'hA9; B = 8'h5B; #100;
A = 8'hA9; B = 8'h5C; #100;
A = 8'hA9; B = 8'h5D; #100;
A = 8'hA9; B = 8'h5E; #100;
A = 8'hA9; B = 8'h5F; #100;
A = 8'hA9; B = 8'h60; #100;
A = 8'hA9; B = 8'h61; #100;
A = 8'hA9; B = 8'h62; #100;
A = 8'hA9; B = 8'h63; #100;
A = 8'hA9; B = 8'h64; #100;
A = 8'hA9; B = 8'h65; #100;
A = 8'hA9; B = 8'h66; #100;
A = 8'hA9; B = 8'h67; #100;
A = 8'hA9; B = 8'h68; #100;
A = 8'hA9; B = 8'h69; #100;
A = 8'hA9; B = 8'h6A; #100;
A = 8'hA9; B = 8'h6B; #100;
A = 8'hA9; B = 8'h6C; #100;
A = 8'hA9; B = 8'h6D; #100;
A = 8'hA9; B = 8'h6E; #100;
A = 8'hA9; B = 8'h6F; #100;
A = 8'hA9; B = 8'h70; #100;
A = 8'hA9; B = 8'h71; #100;
A = 8'hA9; B = 8'h72; #100;
A = 8'hA9; B = 8'h73; #100;
A = 8'hA9; B = 8'h74; #100;
A = 8'hA9; B = 8'h75; #100;
A = 8'hA9; B = 8'h76; #100;
A = 8'hA9; B = 8'h77; #100;
A = 8'hA9; B = 8'h78; #100;
A = 8'hA9; B = 8'h79; #100;
A = 8'hA9; B = 8'h7A; #100;
A = 8'hA9; B = 8'h7B; #100;
A = 8'hA9; B = 8'h7C; #100;
A = 8'hA9; B = 8'h7D; #100;
A = 8'hA9; B = 8'h7E; #100;
A = 8'hA9; B = 8'h7F; #100;
A = 8'hA9; B = 8'h80; #100;
A = 8'hA9; B = 8'h81; #100;
A = 8'hA9; B = 8'h82; #100;
A = 8'hA9; B = 8'h83; #100;
A = 8'hA9; B = 8'h84; #100;
A = 8'hA9; B = 8'h85; #100;
A = 8'hA9; B = 8'h86; #100;
A = 8'hA9; B = 8'h87; #100;
A = 8'hA9; B = 8'h88; #100;
A = 8'hA9; B = 8'h89; #100;
A = 8'hA9; B = 8'h8A; #100;
A = 8'hA9; B = 8'h8B; #100;
A = 8'hA9; B = 8'h8C; #100;
A = 8'hA9; B = 8'h8D; #100;
A = 8'hA9; B = 8'h8E; #100;
A = 8'hA9; B = 8'h8F; #100;
A = 8'hA9; B = 8'h90; #100;
A = 8'hA9; B = 8'h91; #100;
A = 8'hA9; B = 8'h92; #100;
A = 8'hA9; B = 8'h93; #100;
A = 8'hA9; B = 8'h94; #100;
A = 8'hA9; B = 8'h95; #100;
A = 8'hA9; B = 8'h96; #100;
A = 8'hA9; B = 8'h97; #100;
A = 8'hA9; B = 8'h98; #100;
A = 8'hA9; B = 8'h99; #100;
A = 8'hA9; B = 8'h9A; #100;
A = 8'hA9; B = 8'h9B; #100;
A = 8'hA9; B = 8'h9C; #100;
A = 8'hA9; B = 8'h9D; #100;
A = 8'hA9; B = 8'h9E; #100;
A = 8'hA9; B = 8'h9F; #100;
A = 8'hA9; B = 8'hA0; #100;
A = 8'hA9; B = 8'hA1; #100;
A = 8'hA9; B = 8'hA2; #100;
A = 8'hA9; B = 8'hA3; #100;
A = 8'hA9; B = 8'hA4; #100;
A = 8'hA9; B = 8'hA5; #100;
A = 8'hA9; B = 8'hA6; #100;
A = 8'hA9; B = 8'hA7; #100;
A = 8'hA9; B = 8'hA8; #100;
A = 8'hA9; B = 8'hA9; #100;
A = 8'hA9; B = 8'hAA; #100;
A = 8'hA9; B = 8'hAB; #100;
A = 8'hA9; B = 8'hAC; #100;
A = 8'hA9; B = 8'hAD; #100;
A = 8'hA9; B = 8'hAE; #100;
A = 8'hA9; B = 8'hAF; #100;
A = 8'hA9; B = 8'hB0; #100;
A = 8'hA9; B = 8'hB1; #100;
A = 8'hA9; B = 8'hB2; #100;
A = 8'hA9; B = 8'hB3; #100;
A = 8'hA9; B = 8'hB4; #100;
A = 8'hA9; B = 8'hB5; #100;
A = 8'hA9; B = 8'hB6; #100;
A = 8'hA9; B = 8'hB7; #100;
A = 8'hA9; B = 8'hB8; #100;
A = 8'hA9; B = 8'hB9; #100;
A = 8'hA9; B = 8'hBA; #100;
A = 8'hA9; B = 8'hBB; #100;
A = 8'hA9; B = 8'hBC; #100;
A = 8'hA9; B = 8'hBD; #100;
A = 8'hA9; B = 8'hBE; #100;
A = 8'hA9; B = 8'hBF; #100;
A = 8'hA9; B = 8'hC0; #100;
A = 8'hA9; B = 8'hC1; #100;
A = 8'hA9; B = 8'hC2; #100;
A = 8'hA9; B = 8'hC3; #100;
A = 8'hA9; B = 8'hC4; #100;
A = 8'hA9; B = 8'hC5; #100;
A = 8'hA9; B = 8'hC6; #100;
A = 8'hA9; B = 8'hC7; #100;
A = 8'hA9; B = 8'hC8; #100;
A = 8'hA9; B = 8'hC9; #100;
A = 8'hA9; B = 8'hCA; #100;
A = 8'hA9; B = 8'hCB; #100;
A = 8'hA9; B = 8'hCC; #100;
A = 8'hA9; B = 8'hCD; #100;
A = 8'hA9; B = 8'hCE; #100;
A = 8'hA9; B = 8'hCF; #100;
A = 8'hA9; B = 8'hD0; #100;
A = 8'hA9; B = 8'hD1; #100;
A = 8'hA9; B = 8'hD2; #100;
A = 8'hA9; B = 8'hD3; #100;
A = 8'hA9; B = 8'hD4; #100;
A = 8'hA9; B = 8'hD5; #100;
A = 8'hA9; B = 8'hD6; #100;
A = 8'hA9; B = 8'hD7; #100;
A = 8'hA9; B = 8'hD8; #100;
A = 8'hA9; B = 8'hD9; #100;
A = 8'hA9; B = 8'hDA; #100;
A = 8'hA9; B = 8'hDB; #100;
A = 8'hA9; B = 8'hDC; #100;
A = 8'hA9; B = 8'hDD; #100;
A = 8'hA9; B = 8'hDE; #100;
A = 8'hA9; B = 8'hDF; #100;
A = 8'hA9; B = 8'hE0; #100;
A = 8'hA9; B = 8'hE1; #100;
A = 8'hA9; B = 8'hE2; #100;
A = 8'hA9; B = 8'hE3; #100;
A = 8'hA9; B = 8'hE4; #100;
A = 8'hA9; B = 8'hE5; #100;
A = 8'hA9; B = 8'hE6; #100;
A = 8'hA9; B = 8'hE7; #100;
A = 8'hA9; B = 8'hE8; #100;
A = 8'hA9; B = 8'hE9; #100;
A = 8'hA9; B = 8'hEA; #100;
A = 8'hA9; B = 8'hEB; #100;
A = 8'hA9; B = 8'hEC; #100;
A = 8'hA9; B = 8'hED; #100;
A = 8'hA9; B = 8'hEE; #100;
A = 8'hA9; B = 8'hEF; #100;
A = 8'hA9; B = 8'hF0; #100;
A = 8'hA9; B = 8'hF1; #100;
A = 8'hA9; B = 8'hF2; #100;
A = 8'hA9; B = 8'hF3; #100;
A = 8'hA9; B = 8'hF4; #100;
A = 8'hA9; B = 8'hF5; #100;
A = 8'hA9; B = 8'hF6; #100;
A = 8'hA9; B = 8'hF7; #100;
A = 8'hA9; B = 8'hF8; #100;
A = 8'hA9; B = 8'hF9; #100;
A = 8'hA9; B = 8'hFA; #100;
A = 8'hA9; B = 8'hFB; #100;
A = 8'hA9; B = 8'hFC; #100;
A = 8'hA9; B = 8'hFD; #100;
A = 8'hA9; B = 8'hFE; #100;
A = 8'hA9; B = 8'hFF; #100;
A = 8'hAA; B = 8'h0; #100;
A = 8'hAA; B = 8'h1; #100;
A = 8'hAA; B = 8'h2; #100;
A = 8'hAA; B = 8'h3; #100;
A = 8'hAA; B = 8'h4; #100;
A = 8'hAA; B = 8'h5; #100;
A = 8'hAA; B = 8'h6; #100;
A = 8'hAA; B = 8'h7; #100;
A = 8'hAA; B = 8'h8; #100;
A = 8'hAA; B = 8'h9; #100;
A = 8'hAA; B = 8'hA; #100;
A = 8'hAA; B = 8'hB; #100;
A = 8'hAA; B = 8'hC; #100;
A = 8'hAA; B = 8'hD; #100;
A = 8'hAA; B = 8'hE; #100;
A = 8'hAA; B = 8'hF; #100;
A = 8'hAA; B = 8'h10; #100;
A = 8'hAA; B = 8'h11; #100;
A = 8'hAA; B = 8'h12; #100;
A = 8'hAA; B = 8'h13; #100;
A = 8'hAA; B = 8'h14; #100;
A = 8'hAA; B = 8'h15; #100;
A = 8'hAA; B = 8'h16; #100;
A = 8'hAA; B = 8'h17; #100;
A = 8'hAA; B = 8'h18; #100;
A = 8'hAA; B = 8'h19; #100;
A = 8'hAA; B = 8'h1A; #100;
A = 8'hAA; B = 8'h1B; #100;
A = 8'hAA; B = 8'h1C; #100;
A = 8'hAA; B = 8'h1D; #100;
A = 8'hAA; B = 8'h1E; #100;
A = 8'hAA; B = 8'h1F; #100;
A = 8'hAA; B = 8'h20; #100;
A = 8'hAA; B = 8'h21; #100;
A = 8'hAA; B = 8'h22; #100;
A = 8'hAA; B = 8'h23; #100;
A = 8'hAA; B = 8'h24; #100;
A = 8'hAA; B = 8'h25; #100;
A = 8'hAA; B = 8'h26; #100;
A = 8'hAA; B = 8'h27; #100;
A = 8'hAA; B = 8'h28; #100;
A = 8'hAA; B = 8'h29; #100;
A = 8'hAA; B = 8'h2A; #100;
A = 8'hAA; B = 8'h2B; #100;
A = 8'hAA; B = 8'h2C; #100;
A = 8'hAA; B = 8'h2D; #100;
A = 8'hAA; B = 8'h2E; #100;
A = 8'hAA; B = 8'h2F; #100;
A = 8'hAA; B = 8'h30; #100;
A = 8'hAA; B = 8'h31; #100;
A = 8'hAA; B = 8'h32; #100;
A = 8'hAA; B = 8'h33; #100;
A = 8'hAA; B = 8'h34; #100;
A = 8'hAA; B = 8'h35; #100;
A = 8'hAA; B = 8'h36; #100;
A = 8'hAA; B = 8'h37; #100;
A = 8'hAA; B = 8'h38; #100;
A = 8'hAA; B = 8'h39; #100;
A = 8'hAA; B = 8'h3A; #100;
A = 8'hAA; B = 8'h3B; #100;
A = 8'hAA; B = 8'h3C; #100;
A = 8'hAA; B = 8'h3D; #100;
A = 8'hAA; B = 8'h3E; #100;
A = 8'hAA; B = 8'h3F; #100;
A = 8'hAA; B = 8'h40; #100;
A = 8'hAA; B = 8'h41; #100;
A = 8'hAA; B = 8'h42; #100;
A = 8'hAA; B = 8'h43; #100;
A = 8'hAA; B = 8'h44; #100;
A = 8'hAA; B = 8'h45; #100;
A = 8'hAA; B = 8'h46; #100;
A = 8'hAA; B = 8'h47; #100;
A = 8'hAA; B = 8'h48; #100;
A = 8'hAA; B = 8'h49; #100;
A = 8'hAA; B = 8'h4A; #100;
A = 8'hAA; B = 8'h4B; #100;
A = 8'hAA; B = 8'h4C; #100;
A = 8'hAA; B = 8'h4D; #100;
A = 8'hAA; B = 8'h4E; #100;
A = 8'hAA; B = 8'h4F; #100;
A = 8'hAA; B = 8'h50; #100;
A = 8'hAA; B = 8'h51; #100;
A = 8'hAA; B = 8'h52; #100;
A = 8'hAA; B = 8'h53; #100;
A = 8'hAA; B = 8'h54; #100;
A = 8'hAA; B = 8'h55; #100;
A = 8'hAA; B = 8'h56; #100;
A = 8'hAA; B = 8'h57; #100;
A = 8'hAA; B = 8'h58; #100;
A = 8'hAA; B = 8'h59; #100;
A = 8'hAA; B = 8'h5A; #100;
A = 8'hAA; B = 8'h5B; #100;
A = 8'hAA; B = 8'h5C; #100;
A = 8'hAA; B = 8'h5D; #100;
A = 8'hAA; B = 8'h5E; #100;
A = 8'hAA; B = 8'h5F; #100;
A = 8'hAA; B = 8'h60; #100;
A = 8'hAA; B = 8'h61; #100;
A = 8'hAA; B = 8'h62; #100;
A = 8'hAA; B = 8'h63; #100;
A = 8'hAA; B = 8'h64; #100;
A = 8'hAA; B = 8'h65; #100;
A = 8'hAA; B = 8'h66; #100;
A = 8'hAA; B = 8'h67; #100;
A = 8'hAA; B = 8'h68; #100;
A = 8'hAA; B = 8'h69; #100;
A = 8'hAA; B = 8'h6A; #100;
A = 8'hAA; B = 8'h6B; #100;
A = 8'hAA; B = 8'h6C; #100;
A = 8'hAA; B = 8'h6D; #100;
A = 8'hAA; B = 8'h6E; #100;
A = 8'hAA; B = 8'h6F; #100;
A = 8'hAA; B = 8'h70; #100;
A = 8'hAA; B = 8'h71; #100;
A = 8'hAA; B = 8'h72; #100;
A = 8'hAA; B = 8'h73; #100;
A = 8'hAA; B = 8'h74; #100;
A = 8'hAA; B = 8'h75; #100;
A = 8'hAA; B = 8'h76; #100;
A = 8'hAA; B = 8'h77; #100;
A = 8'hAA; B = 8'h78; #100;
A = 8'hAA; B = 8'h79; #100;
A = 8'hAA; B = 8'h7A; #100;
A = 8'hAA; B = 8'h7B; #100;
A = 8'hAA; B = 8'h7C; #100;
A = 8'hAA; B = 8'h7D; #100;
A = 8'hAA; B = 8'h7E; #100;
A = 8'hAA; B = 8'h7F; #100;
A = 8'hAA; B = 8'h80; #100;
A = 8'hAA; B = 8'h81; #100;
A = 8'hAA; B = 8'h82; #100;
A = 8'hAA; B = 8'h83; #100;
A = 8'hAA; B = 8'h84; #100;
A = 8'hAA; B = 8'h85; #100;
A = 8'hAA; B = 8'h86; #100;
A = 8'hAA; B = 8'h87; #100;
A = 8'hAA; B = 8'h88; #100;
A = 8'hAA; B = 8'h89; #100;
A = 8'hAA; B = 8'h8A; #100;
A = 8'hAA; B = 8'h8B; #100;
A = 8'hAA; B = 8'h8C; #100;
A = 8'hAA; B = 8'h8D; #100;
A = 8'hAA; B = 8'h8E; #100;
A = 8'hAA; B = 8'h8F; #100;
A = 8'hAA; B = 8'h90; #100;
A = 8'hAA; B = 8'h91; #100;
A = 8'hAA; B = 8'h92; #100;
A = 8'hAA; B = 8'h93; #100;
A = 8'hAA; B = 8'h94; #100;
A = 8'hAA; B = 8'h95; #100;
A = 8'hAA; B = 8'h96; #100;
A = 8'hAA; B = 8'h97; #100;
A = 8'hAA; B = 8'h98; #100;
A = 8'hAA; B = 8'h99; #100;
A = 8'hAA; B = 8'h9A; #100;
A = 8'hAA; B = 8'h9B; #100;
A = 8'hAA; B = 8'h9C; #100;
A = 8'hAA; B = 8'h9D; #100;
A = 8'hAA; B = 8'h9E; #100;
A = 8'hAA; B = 8'h9F; #100;
A = 8'hAA; B = 8'hA0; #100;
A = 8'hAA; B = 8'hA1; #100;
A = 8'hAA; B = 8'hA2; #100;
A = 8'hAA; B = 8'hA3; #100;
A = 8'hAA; B = 8'hA4; #100;
A = 8'hAA; B = 8'hA5; #100;
A = 8'hAA; B = 8'hA6; #100;
A = 8'hAA; B = 8'hA7; #100;
A = 8'hAA; B = 8'hA8; #100;
A = 8'hAA; B = 8'hA9; #100;
A = 8'hAA; B = 8'hAA; #100;
A = 8'hAA; B = 8'hAB; #100;
A = 8'hAA; B = 8'hAC; #100;
A = 8'hAA; B = 8'hAD; #100;
A = 8'hAA; B = 8'hAE; #100;
A = 8'hAA; B = 8'hAF; #100;
A = 8'hAA; B = 8'hB0; #100;
A = 8'hAA; B = 8'hB1; #100;
A = 8'hAA; B = 8'hB2; #100;
A = 8'hAA; B = 8'hB3; #100;
A = 8'hAA; B = 8'hB4; #100;
A = 8'hAA; B = 8'hB5; #100;
A = 8'hAA; B = 8'hB6; #100;
A = 8'hAA; B = 8'hB7; #100;
A = 8'hAA; B = 8'hB8; #100;
A = 8'hAA; B = 8'hB9; #100;
A = 8'hAA; B = 8'hBA; #100;
A = 8'hAA; B = 8'hBB; #100;
A = 8'hAA; B = 8'hBC; #100;
A = 8'hAA; B = 8'hBD; #100;
A = 8'hAA; B = 8'hBE; #100;
A = 8'hAA; B = 8'hBF; #100;
A = 8'hAA; B = 8'hC0; #100;
A = 8'hAA; B = 8'hC1; #100;
A = 8'hAA; B = 8'hC2; #100;
A = 8'hAA; B = 8'hC3; #100;
A = 8'hAA; B = 8'hC4; #100;
A = 8'hAA; B = 8'hC5; #100;
A = 8'hAA; B = 8'hC6; #100;
A = 8'hAA; B = 8'hC7; #100;
A = 8'hAA; B = 8'hC8; #100;
A = 8'hAA; B = 8'hC9; #100;
A = 8'hAA; B = 8'hCA; #100;
A = 8'hAA; B = 8'hCB; #100;
A = 8'hAA; B = 8'hCC; #100;
A = 8'hAA; B = 8'hCD; #100;
A = 8'hAA; B = 8'hCE; #100;
A = 8'hAA; B = 8'hCF; #100;
A = 8'hAA; B = 8'hD0; #100;
A = 8'hAA; B = 8'hD1; #100;
A = 8'hAA; B = 8'hD2; #100;
A = 8'hAA; B = 8'hD3; #100;
A = 8'hAA; B = 8'hD4; #100;
A = 8'hAA; B = 8'hD5; #100;
A = 8'hAA; B = 8'hD6; #100;
A = 8'hAA; B = 8'hD7; #100;
A = 8'hAA; B = 8'hD8; #100;
A = 8'hAA; B = 8'hD9; #100;
A = 8'hAA; B = 8'hDA; #100;
A = 8'hAA; B = 8'hDB; #100;
A = 8'hAA; B = 8'hDC; #100;
A = 8'hAA; B = 8'hDD; #100;
A = 8'hAA; B = 8'hDE; #100;
A = 8'hAA; B = 8'hDF; #100;
A = 8'hAA; B = 8'hE0; #100;
A = 8'hAA; B = 8'hE1; #100;
A = 8'hAA; B = 8'hE2; #100;
A = 8'hAA; B = 8'hE3; #100;
A = 8'hAA; B = 8'hE4; #100;
A = 8'hAA; B = 8'hE5; #100;
A = 8'hAA; B = 8'hE6; #100;
A = 8'hAA; B = 8'hE7; #100;
A = 8'hAA; B = 8'hE8; #100;
A = 8'hAA; B = 8'hE9; #100;
A = 8'hAA; B = 8'hEA; #100;
A = 8'hAA; B = 8'hEB; #100;
A = 8'hAA; B = 8'hEC; #100;
A = 8'hAA; B = 8'hED; #100;
A = 8'hAA; B = 8'hEE; #100;
A = 8'hAA; B = 8'hEF; #100;
A = 8'hAA; B = 8'hF0; #100;
A = 8'hAA; B = 8'hF1; #100;
A = 8'hAA; B = 8'hF2; #100;
A = 8'hAA; B = 8'hF3; #100;
A = 8'hAA; B = 8'hF4; #100;
A = 8'hAA; B = 8'hF5; #100;
A = 8'hAA; B = 8'hF6; #100;
A = 8'hAA; B = 8'hF7; #100;
A = 8'hAA; B = 8'hF8; #100;
A = 8'hAA; B = 8'hF9; #100;
A = 8'hAA; B = 8'hFA; #100;
A = 8'hAA; B = 8'hFB; #100;
A = 8'hAA; B = 8'hFC; #100;
A = 8'hAA; B = 8'hFD; #100;
A = 8'hAA; B = 8'hFE; #100;
A = 8'hAA; B = 8'hFF; #100;
A = 8'hAB; B = 8'h0; #100;
A = 8'hAB; B = 8'h1; #100;
A = 8'hAB; B = 8'h2; #100;
A = 8'hAB; B = 8'h3; #100;
A = 8'hAB; B = 8'h4; #100;
A = 8'hAB; B = 8'h5; #100;
A = 8'hAB; B = 8'h6; #100;
A = 8'hAB; B = 8'h7; #100;
A = 8'hAB; B = 8'h8; #100;
A = 8'hAB; B = 8'h9; #100;
A = 8'hAB; B = 8'hA; #100;
A = 8'hAB; B = 8'hB; #100;
A = 8'hAB; B = 8'hC; #100;
A = 8'hAB; B = 8'hD; #100;
A = 8'hAB; B = 8'hE; #100;
A = 8'hAB; B = 8'hF; #100;
A = 8'hAB; B = 8'h10; #100;
A = 8'hAB; B = 8'h11; #100;
A = 8'hAB; B = 8'h12; #100;
A = 8'hAB; B = 8'h13; #100;
A = 8'hAB; B = 8'h14; #100;
A = 8'hAB; B = 8'h15; #100;
A = 8'hAB; B = 8'h16; #100;
A = 8'hAB; B = 8'h17; #100;
A = 8'hAB; B = 8'h18; #100;
A = 8'hAB; B = 8'h19; #100;
A = 8'hAB; B = 8'h1A; #100;
A = 8'hAB; B = 8'h1B; #100;
A = 8'hAB; B = 8'h1C; #100;
A = 8'hAB; B = 8'h1D; #100;
A = 8'hAB; B = 8'h1E; #100;
A = 8'hAB; B = 8'h1F; #100;
A = 8'hAB; B = 8'h20; #100;
A = 8'hAB; B = 8'h21; #100;
A = 8'hAB; B = 8'h22; #100;
A = 8'hAB; B = 8'h23; #100;
A = 8'hAB; B = 8'h24; #100;
A = 8'hAB; B = 8'h25; #100;
A = 8'hAB; B = 8'h26; #100;
A = 8'hAB; B = 8'h27; #100;
A = 8'hAB; B = 8'h28; #100;
A = 8'hAB; B = 8'h29; #100;
A = 8'hAB; B = 8'h2A; #100;
A = 8'hAB; B = 8'h2B; #100;
A = 8'hAB; B = 8'h2C; #100;
A = 8'hAB; B = 8'h2D; #100;
A = 8'hAB; B = 8'h2E; #100;
A = 8'hAB; B = 8'h2F; #100;
A = 8'hAB; B = 8'h30; #100;
A = 8'hAB; B = 8'h31; #100;
A = 8'hAB; B = 8'h32; #100;
A = 8'hAB; B = 8'h33; #100;
A = 8'hAB; B = 8'h34; #100;
A = 8'hAB; B = 8'h35; #100;
A = 8'hAB; B = 8'h36; #100;
A = 8'hAB; B = 8'h37; #100;
A = 8'hAB; B = 8'h38; #100;
A = 8'hAB; B = 8'h39; #100;
A = 8'hAB; B = 8'h3A; #100;
A = 8'hAB; B = 8'h3B; #100;
A = 8'hAB; B = 8'h3C; #100;
A = 8'hAB; B = 8'h3D; #100;
A = 8'hAB; B = 8'h3E; #100;
A = 8'hAB; B = 8'h3F; #100;
A = 8'hAB; B = 8'h40; #100;
A = 8'hAB; B = 8'h41; #100;
A = 8'hAB; B = 8'h42; #100;
A = 8'hAB; B = 8'h43; #100;
A = 8'hAB; B = 8'h44; #100;
A = 8'hAB; B = 8'h45; #100;
A = 8'hAB; B = 8'h46; #100;
A = 8'hAB; B = 8'h47; #100;
A = 8'hAB; B = 8'h48; #100;
A = 8'hAB; B = 8'h49; #100;
A = 8'hAB; B = 8'h4A; #100;
A = 8'hAB; B = 8'h4B; #100;
A = 8'hAB; B = 8'h4C; #100;
A = 8'hAB; B = 8'h4D; #100;
A = 8'hAB; B = 8'h4E; #100;
A = 8'hAB; B = 8'h4F; #100;
A = 8'hAB; B = 8'h50; #100;
A = 8'hAB; B = 8'h51; #100;
A = 8'hAB; B = 8'h52; #100;
A = 8'hAB; B = 8'h53; #100;
A = 8'hAB; B = 8'h54; #100;
A = 8'hAB; B = 8'h55; #100;
A = 8'hAB; B = 8'h56; #100;
A = 8'hAB; B = 8'h57; #100;
A = 8'hAB; B = 8'h58; #100;
A = 8'hAB; B = 8'h59; #100;
A = 8'hAB; B = 8'h5A; #100;
A = 8'hAB; B = 8'h5B; #100;
A = 8'hAB; B = 8'h5C; #100;
A = 8'hAB; B = 8'h5D; #100;
A = 8'hAB; B = 8'h5E; #100;
A = 8'hAB; B = 8'h5F; #100;
A = 8'hAB; B = 8'h60; #100;
A = 8'hAB; B = 8'h61; #100;
A = 8'hAB; B = 8'h62; #100;
A = 8'hAB; B = 8'h63; #100;
A = 8'hAB; B = 8'h64; #100;
A = 8'hAB; B = 8'h65; #100;
A = 8'hAB; B = 8'h66; #100;
A = 8'hAB; B = 8'h67; #100;
A = 8'hAB; B = 8'h68; #100;
A = 8'hAB; B = 8'h69; #100;
A = 8'hAB; B = 8'h6A; #100;
A = 8'hAB; B = 8'h6B; #100;
A = 8'hAB; B = 8'h6C; #100;
A = 8'hAB; B = 8'h6D; #100;
A = 8'hAB; B = 8'h6E; #100;
A = 8'hAB; B = 8'h6F; #100;
A = 8'hAB; B = 8'h70; #100;
A = 8'hAB; B = 8'h71; #100;
A = 8'hAB; B = 8'h72; #100;
A = 8'hAB; B = 8'h73; #100;
A = 8'hAB; B = 8'h74; #100;
A = 8'hAB; B = 8'h75; #100;
A = 8'hAB; B = 8'h76; #100;
A = 8'hAB; B = 8'h77; #100;
A = 8'hAB; B = 8'h78; #100;
A = 8'hAB; B = 8'h79; #100;
A = 8'hAB; B = 8'h7A; #100;
A = 8'hAB; B = 8'h7B; #100;
A = 8'hAB; B = 8'h7C; #100;
A = 8'hAB; B = 8'h7D; #100;
A = 8'hAB; B = 8'h7E; #100;
A = 8'hAB; B = 8'h7F; #100;
A = 8'hAB; B = 8'h80; #100;
A = 8'hAB; B = 8'h81; #100;
A = 8'hAB; B = 8'h82; #100;
A = 8'hAB; B = 8'h83; #100;
A = 8'hAB; B = 8'h84; #100;
A = 8'hAB; B = 8'h85; #100;
A = 8'hAB; B = 8'h86; #100;
A = 8'hAB; B = 8'h87; #100;
A = 8'hAB; B = 8'h88; #100;
A = 8'hAB; B = 8'h89; #100;
A = 8'hAB; B = 8'h8A; #100;
A = 8'hAB; B = 8'h8B; #100;
A = 8'hAB; B = 8'h8C; #100;
A = 8'hAB; B = 8'h8D; #100;
A = 8'hAB; B = 8'h8E; #100;
A = 8'hAB; B = 8'h8F; #100;
A = 8'hAB; B = 8'h90; #100;
A = 8'hAB; B = 8'h91; #100;
A = 8'hAB; B = 8'h92; #100;
A = 8'hAB; B = 8'h93; #100;
A = 8'hAB; B = 8'h94; #100;
A = 8'hAB; B = 8'h95; #100;
A = 8'hAB; B = 8'h96; #100;
A = 8'hAB; B = 8'h97; #100;
A = 8'hAB; B = 8'h98; #100;
A = 8'hAB; B = 8'h99; #100;
A = 8'hAB; B = 8'h9A; #100;
A = 8'hAB; B = 8'h9B; #100;
A = 8'hAB; B = 8'h9C; #100;
A = 8'hAB; B = 8'h9D; #100;
A = 8'hAB; B = 8'h9E; #100;
A = 8'hAB; B = 8'h9F; #100;
A = 8'hAB; B = 8'hA0; #100;
A = 8'hAB; B = 8'hA1; #100;
A = 8'hAB; B = 8'hA2; #100;
A = 8'hAB; B = 8'hA3; #100;
A = 8'hAB; B = 8'hA4; #100;
A = 8'hAB; B = 8'hA5; #100;
A = 8'hAB; B = 8'hA6; #100;
A = 8'hAB; B = 8'hA7; #100;
A = 8'hAB; B = 8'hA8; #100;
A = 8'hAB; B = 8'hA9; #100;
A = 8'hAB; B = 8'hAA; #100;
A = 8'hAB; B = 8'hAB; #100;
A = 8'hAB; B = 8'hAC; #100;
A = 8'hAB; B = 8'hAD; #100;
A = 8'hAB; B = 8'hAE; #100;
A = 8'hAB; B = 8'hAF; #100;
A = 8'hAB; B = 8'hB0; #100;
A = 8'hAB; B = 8'hB1; #100;
A = 8'hAB; B = 8'hB2; #100;
A = 8'hAB; B = 8'hB3; #100;
A = 8'hAB; B = 8'hB4; #100;
A = 8'hAB; B = 8'hB5; #100;
A = 8'hAB; B = 8'hB6; #100;
A = 8'hAB; B = 8'hB7; #100;
A = 8'hAB; B = 8'hB8; #100;
A = 8'hAB; B = 8'hB9; #100;
A = 8'hAB; B = 8'hBA; #100;
A = 8'hAB; B = 8'hBB; #100;
A = 8'hAB; B = 8'hBC; #100;
A = 8'hAB; B = 8'hBD; #100;
A = 8'hAB; B = 8'hBE; #100;
A = 8'hAB; B = 8'hBF; #100;
A = 8'hAB; B = 8'hC0; #100;
A = 8'hAB; B = 8'hC1; #100;
A = 8'hAB; B = 8'hC2; #100;
A = 8'hAB; B = 8'hC3; #100;
A = 8'hAB; B = 8'hC4; #100;
A = 8'hAB; B = 8'hC5; #100;
A = 8'hAB; B = 8'hC6; #100;
A = 8'hAB; B = 8'hC7; #100;
A = 8'hAB; B = 8'hC8; #100;
A = 8'hAB; B = 8'hC9; #100;
A = 8'hAB; B = 8'hCA; #100;
A = 8'hAB; B = 8'hCB; #100;
A = 8'hAB; B = 8'hCC; #100;
A = 8'hAB; B = 8'hCD; #100;
A = 8'hAB; B = 8'hCE; #100;
A = 8'hAB; B = 8'hCF; #100;
A = 8'hAB; B = 8'hD0; #100;
A = 8'hAB; B = 8'hD1; #100;
A = 8'hAB; B = 8'hD2; #100;
A = 8'hAB; B = 8'hD3; #100;
A = 8'hAB; B = 8'hD4; #100;
A = 8'hAB; B = 8'hD5; #100;
A = 8'hAB; B = 8'hD6; #100;
A = 8'hAB; B = 8'hD7; #100;
A = 8'hAB; B = 8'hD8; #100;
A = 8'hAB; B = 8'hD9; #100;
A = 8'hAB; B = 8'hDA; #100;
A = 8'hAB; B = 8'hDB; #100;
A = 8'hAB; B = 8'hDC; #100;
A = 8'hAB; B = 8'hDD; #100;
A = 8'hAB; B = 8'hDE; #100;
A = 8'hAB; B = 8'hDF; #100;
A = 8'hAB; B = 8'hE0; #100;
A = 8'hAB; B = 8'hE1; #100;
A = 8'hAB; B = 8'hE2; #100;
A = 8'hAB; B = 8'hE3; #100;
A = 8'hAB; B = 8'hE4; #100;
A = 8'hAB; B = 8'hE5; #100;
A = 8'hAB; B = 8'hE6; #100;
A = 8'hAB; B = 8'hE7; #100;
A = 8'hAB; B = 8'hE8; #100;
A = 8'hAB; B = 8'hE9; #100;
A = 8'hAB; B = 8'hEA; #100;
A = 8'hAB; B = 8'hEB; #100;
A = 8'hAB; B = 8'hEC; #100;
A = 8'hAB; B = 8'hED; #100;
A = 8'hAB; B = 8'hEE; #100;
A = 8'hAB; B = 8'hEF; #100;
A = 8'hAB; B = 8'hF0; #100;
A = 8'hAB; B = 8'hF1; #100;
A = 8'hAB; B = 8'hF2; #100;
A = 8'hAB; B = 8'hF3; #100;
A = 8'hAB; B = 8'hF4; #100;
A = 8'hAB; B = 8'hF5; #100;
A = 8'hAB; B = 8'hF6; #100;
A = 8'hAB; B = 8'hF7; #100;
A = 8'hAB; B = 8'hF8; #100;
A = 8'hAB; B = 8'hF9; #100;
A = 8'hAB; B = 8'hFA; #100;
A = 8'hAB; B = 8'hFB; #100;
A = 8'hAB; B = 8'hFC; #100;
A = 8'hAB; B = 8'hFD; #100;
A = 8'hAB; B = 8'hFE; #100;
A = 8'hAB; B = 8'hFF; #100;
A = 8'hAC; B = 8'h0; #100;
A = 8'hAC; B = 8'h1; #100;
A = 8'hAC; B = 8'h2; #100;
A = 8'hAC; B = 8'h3; #100;
A = 8'hAC; B = 8'h4; #100;
A = 8'hAC; B = 8'h5; #100;
A = 8'hAC; B = 8'h6; #100;
A = 8'hAC; B = 8'h7; #100;
A = 8'hAC; B = 8'h8; #100;
A = 8'hAC; B = 8'h9; #100;
A = 8'hAC; B = 8'hA; #100;
A = 8'hAC; B = 8'hB; #100;
A = 8'hAC; B = 8'hC; #100;
A = 8'hAC; B = 8'hD; #100;
A = 8'hAC; B = 8'hE; #100;
A = 8'hAC; B = 8'hF; #100;
A = 8'hAC; B = 8'h10; #100;
A = 8'hAC; B = 8'h11; #100;
A = 8'hAC; B = 8'h12; #100;
A = 8'hAC; B = 8'h13; #100;
A = 8'hAC; B = 8'h14; #100;
A = 8'hAC; B = 8'h15; #100;
A = 8'hAC; B = 8'h16; #100;
A = 8'hAC; B = 8'h17; #100;
A = 8'hAC; B = 8'h18; #100;
A = 8'hAC; B = 8'h19; #100;
A = 8'hAC; B = 8'h1A; #100;
A = 8'hAC; B = 8'h1B; #100;
A = 8'hAC; B = 8'h1C; #100;
A = 8'hAC; B = 8'h1D; #100;
A = 8'hAC; B = 8'h1E; #100;
A = 8'hAC; B = 8'h1F; #100;
A = 8'hAC; B = 8'h20; #100;
A = 8'hAC; B = 8'h21; #100;
A = 8'hAC; B = 8'h22; #100;
A = 8'hAC; B = 8'h23; #100;
A = 8'hAC; B = 8'h24; #100;
A = 8'hAC; B = 8'h25; #100;
A = 8'hAC; B = 8'h26; #100;
A = 8'hAC; B = 8'h27; #100;
A = 8'hAC; B = 8'h28; #100;
A = 8'hAC; B = 8'h29; #100;
A = 8'hAC; B = 8'h2A; #100;
A = 8'hAC; B = 8'h2B; #100;
A = 8'hAC; B = 8'h2C; #100;
A = 8'hAC; B = 8'h2D; #100;
A = 8'hAC; B = 8'h2E; #100;
A = 8'hAC; B = 8'h2F; #100;
A = 8'hAC; B = 8'h30; #100;
A = 8'hAC; B = 8'h31; #100;
A = 8'hAC; B = 8'h32; #100;
A = 8'hAC; B = 8'h33; #100;
A = 8'hAC; B = 8'h34; #100;
A = 8'hAC; B = 8'h35; #100;
A = 8'hAC; B = 8'h36; #100;
A = 8'hAC; B = 8'h37; #100;
A = 8'hAC; B = 8'h38; #100;
A = 8'hAC; B = 8'h39; #100;
A = 8'hAC; B = 8'h3A; #100;
A = 8'hAC; B = 8'h3B; #100;
A = 8'hAC; B = 8'h3C; #100;
A = 8'hAC; B = 8'h3D; #100;
A = 8'hAC; B = 8'h3E; #100;
A = 8'hAC; B = 8'h3F; #100;
A = 8'hAC; B = 8'h40; #100;
A = 8'hAC; B = 8'h41; #100;
A = 8'hAC; B = 8'h42; #100;
A = 8'hAC; B = 8'h43; #100;
A = 8'hAC; B = 8'h44; #100;
A = 8'hAC; B = 8'h45; #100;
A = 8'hAC; B = 8'h46; #100;
A = 8'hAC; B = 8'h47; #100;
A = 8'hAC; B = 8'h48; #100;
A = 8'hAC; B = 8'h49; #100;
A = 8'hAC; B = 8'h4A; #100;
A = 8'hAC; B = 8'h4B; #100;
A = 8'hAC; B = 8'h4C; #100;
A = 8'hAC; B = 8'h4D; #100;
A = 8'hAC; B = 8'h4E; #100;
A = 8'hAC; B = 8'h4F; #100;
A = 8'hAC; B = 8'h50; #100;
A = 8'hAC; B = 8'h51; #100;
A = 8'hAC; B = 8'h52; #100;
A = 8'hAC; B = 8'h53; #100;
A = 8'hAC; B = 8'h54; #100;
A = 8'hAC; B = 8'h55; #100;
A = 8'hAC; B = 8'h56; #100;
A = 8'hAC; B = 8'h57; #100;
A = 8'hAC; B = 8'h58; #100;
A = 8'hAC; B = 8'h59; #100;
A = 8'hAC; B = 8'h5A; #100;
A = 8'hAC; B = 8'h5B; #100;
A = 8'hAC; B = 8'h5C; #100;
A = 8'hAC; B = 8'h5D; #100;
A = 8'hAC; B = 8'h5E; #100;
A = 8'hAC; B = 8'h5F; #100;
A = 8'hAC; B = 8'h60; #100;
A = 8'hAC; B = 8'h61; #100;
A = 8'hAC; B = 8'h62; #100;
A = 8'hAC; B = 8'h63; #100;
A = 8'hAC; B = 8'h64; #100;
A = 8'hAC; B = 8'h65; #100;
A = 8'hAC; B = 8'h66; #100;
A = 8'hAC; B = 8'h67; #100;
A = 8'hAC; B = 8'h68; #100;
A = 8'hAC; B = 8'h69; #100;
A = 8'hAC; B = 8'h6A; #100;
A = 8'hAC; B = 8'h6B; #100;
A = 8'hAC; B = 8'h6C; #100;
A = 8'hAC; B = 8'h6D; #100;
A = 8'hAC; B = 8'h6E; #100;
A = 8'hAC; B = 8'h6F; #100;
A = 8'hAC; B = 8'h70; #100;
A = 8'hAC; B = 8'h71; #100;
A = 8'hAC; B = 8'h72; #100;
A = 8'hAC; B = 8'h73; #100;
A = 8'hAC; B = 8'h74; #100;
A = 8'hAC; B = 8'h75; #100;
A = 8'hAC; B = 8'h76; #100;
A = 8'hAC; B = 8'h77; #100;
A = 8'hAC; B = 8'h78; #100;
A = 8'hAC; B = 8'h79; #100;
A = 8'hAC; B = 8'h7A; #100;
A = 8'hAC; B = 8'h7B; #100;
A = 8'hAC; B = 8'h7C; #100;
A = 8'hAC; B = 8'h7D; #100;
A = 8'hAC; B = 8'h7E; #100;
A = 8'hAC; B = 8'h7F; #100;
A = 8'hAC; B = 8'h80; #100;
A = 8'hAC; B = 8'h81; #100;
A = 8'hAC; B = 8'h82; #100;
A = 8'hAC; B = 8'h83; #100;
A = 8'hAC; B = 8'h84; #100;
A = 8'hAC; B = 8'h85; #100;
A = 8'hAC; B = 8'h86; #100;
A = 8'hAC; B = 8'h87; #100;
A = 8'hAC; B = 8'h88; #100;
A = 8'hAC; B = 8'h89; #100;
A = 8'hAC; B = 8'h8A; #100;
A = 8'hAC; B = 8'h8B; #100;
A = 8'hAC; B = 8'h8C; #100;
A = 8'hAC; B = 8'h8D; #100;
A = 8'hAC; B = 8'h8E; #100;
A = 8'hAC; B = 8'h8F; #100;
A = 8'hAC; B = 8'h90; #100;
A = 8'hAC; B = 8'h91; #100;
A = 8'hAC; B = 8'h92; #100;
A = 8'hAC; B = 8'h93; #100;
A = 8'hAC; B = 8'h94; #100;
A = 8'hAC; B = 8'h95; #100;
A = 8'hAC; B = 8'h96; #100;
A = 8'hAC; B = 8'h97; #100;
A = 8'hAC; B = 8'h98; #100;
A = 8'hAC; B = 8'h99; #100;
A = 8'hAC; B = 8'h9A; #100;
A = 8'hAC; B = 8'h9B; #100;
A = 8'hAC; B = 8'h9C; #100;
A = 8'hAC; B = 8'h9D; #100;
A = 8'hAC; B = 8'h9E; #100;
A = 8'hAC; B = 8'h9F; #100;
A = 8'hAC; B = 8'hA0; #100;
A = 8'hAC; B = 8'hA1; #100;
A = 8'hAC; B = 8'hA2; #100;
A = 8'hAC; B = 8'hA3; #100;
A = 8'hAC; B = 8'hA4; #100;
A = 8'hAC; B = 8'hA5; #100;
A = 8'hAC; B = 8'hA6; #100;
A = 8'hAC; B = 8'hA7; #100;
A = 8'hAC; B = 8'hA8; #100;
A = 8'hAC; B = 8'hA9; #100;
A = 8'hAC; B = 8'hAA; #100;
A = 8'hAC; B = 8'hAB; #100;
A = 8'hAC; B = 8'hAC; #100;
A = 8'hAC; B = 8'hAD; #100;
A = 8'hAC; B = 8'hAE; #100;
A = 8'hAC; B = 8'hAF; #100;
A = 8'hAC; B = 8'hB0; #100;
A = 8'hAC; B = 8'hB1; #100;
A = 8'hAC; B = 8'hB2; #100;
A = 8'hAC; B = 8'hB3; #100;
A = 8'hAC; B = 8'hB4; #100;
A = 8'hAC; B = 8'hB5; #100;
A = 8'hAC; B = 8'hB6; #100;
A = 8'hAC; B = 8'hB7; #100;
A = 8'hAC; B = 8'hB8; #100;
A = 8'hAC; B = 8'hB9; #100;
A = 8'hAC; B = 8'hBA; #100;
A = 8'hAC; B = 8'hBB; #100;
A = 8'hAC; B = 8'hBC; #100;
A = 8'hAC; B = 8'hBD; #100;
A = 8'hAC; B = 8'hBE; #100;
A = 8'hAC; B = 8'hBF; #100;
A = 8'hAC; B = 8'hC0; #100;
A = 8'hAC; B = 8'hC1; #100;
A = 8'hAC; B = 8'hC2; #100;
A = 8'hAC; B = 8'hC3; #100;
A = 8'hAC; B = 8'hC4; #100;
A = 8'hAC; B = 8'hC5; #100;
A = 8'hAC; B = 8'hC6; #100;
A = 8'hAC; B = 8'hC7; #100;
A = 8'hAC; B = 8'hC8; #100;
A = 8'hAC; B = 8'hC9; #100;
A = 8'hAC; B = 8'hCA; #100;
A = 8'hAC; B = 8'hCB; #100;
A = 8'hAC; B = 8'hCC; #100;
A = 8'hAC; B = 8'hCD; #100;
A = 8'hAC; B = 8'hCE; #100;
A = 8'hAC; B = 8'hCF; #100;
A = 8'hAC; B = 8'hD0; #100;
A = 8'hAC; B = 8'hD1; #100;
A = 8'hAC; B = 8'hD2; #100;
A = 8'hAC; B = 8'hD3; #100;
A = 8'hAC; B = 8'hD4; #100;
A = 8'hAC; B = 8'hD5; #100;
A = 8'hAC; B = 8'hD6; #100;
A = 8'hAC; B = 8'hD7; #100;
A = 8'hAC; B = 8'hD8; #100;
A = 8'hAC; B = 8'hD9; #100;
A = 8'hAC; B = 8'hDA; #100;
A = 8'hAC; B = 8'hDB; #100;
A = 8'hAC; B = 8'hDC; #100;
A = 8'hAC; B = 8'hDD; #100;
A = 8'hAC; B = 8'hDE; #100;
A = 8'hAC; B = 8'hDF; #100;
A = 8'hAC; B = 8'hE0; #100;
A = 8'hAC; B = 8'hE1; #100;
A = 8'hAC; B = 8'hE2; #100;
A = 8'hAC; B = 8'hE3; #100;
A = 8'hAC; B = 8'hE4; #100;
A = 8'hAC; B = 8'hE5; #100;
A = 8'hAC; B = 8'hE6; #100;
A = 8'hAC; B = 8'hE7; #100;
A = 8'hAC; B = 8'hE8; #100;
A = 8'hAC; B = 8'hE9; #100;
A = 8'hAC; B = 8'hEA; #100;
A = 8'hAC; B = 8'hEB; #100;
A = 8'hAC; B = 8'hEC; #100;
A = 8'hAC; B = 8'hED; #100;
A = 8'hAC; B = 8'hEE; #100;
A = 8'hAC; B = 8'hEF; #100;
A = 8'hAC; B = 8'hF0; #100;
A = 8'hAC; B = 8'hF1; #100;
A = 8'hAC; B = 8'hF2; #100;
A = 8'hAC; B = 8'hF3; #100;
A = 8'hAC; B = 8'hF4; #100;
A = 8'hAC; B = 8'hF5; #100;
A = 8'hAC; B = 8'hF6; #100;
A = 8'hAC; B = 8'hF7; #100;
A = 8'hAC; B = 8'hF8; #100;
A = 8'hAC; B = 8'hF9; #100;
A = 8'hAC; B = 8'hFA; #100;
A = 8'hAC; B = 8'hFB; #100;
A = 8'hAC; B = 8'hFC; #100;
A = 8'hAC; B = 8'hFD; #100;
A = 8'hAC; B = 8'hFE; #100;
A = 8'hAC; B = 8'hFF; #100;
A = 8'hAD; B = 8'h0; #100;
A = 8'hAD; B = 8'h1; #100;
A = 8'hAD; B = 8'h2; #100;
A = 8'hAD; B = 8'h3; #100;
A = 8'hAD; B = 8'h4; #100;
A = 8'hAD; B = 8'h5; #100;
A = 8'hAD; B = 8'h6; #100;
A = 8'hAD; B = 8'h7; #100;
A = 8'hAD; B = 8'h8; #100;
A = 8'hAD; B = 8'h9; #100;
A = 8'hAD; B = 8'hA; #100;
A = 8'hAD; B = 8'hB; #100;
A = 8'hAD; B = 8'hC; #100;
A = 8'hAD; B = 8'hD; #100;
A = 8'hAD; B = 8'hE; #100;
A = 8'hAD; B = 8'hF; #100;
A = 8'hAD; B = 8'h10; #100;
A = 8'hAD; B = 8'h11; #100;
A = 8'hAD; B = 8'h12; #100;
A = 8'hAD; B = 8'h13; #100;
A = 8'hAD; B = 8'h14; #100;
A = 8'hAD; B = 8'h15; #100;
A = 8'hAD; B = 8'h16; #100;
A = 8'hAD; B = 8'h17; #100;
A = 8'hAD; B = 8'h18; #100;
A = 8'hAD; B = 8'h19; #100;
A = 8'hAD; B = 8'h1A; #100;
A = 8'hAD; B = 8'h1B; #100;
A = 8'hAD; B = 8'h1C; #100;
A = 8'hAD; B = 8'h1D; #100;
A = 8'hAD; B = 8'h1E; #100;
A = 8'hAD; B = 8'h1F; #100;
A = 8'hAD; B = 8'h20; #100;
A = 8'hAD; B = 8'h21; #100;
A = 8'hAD; B = 8'h22; #100;
A = 8'hAD; B = 8'h23; #100;
A = 8'hAD; B = 8'h24; #100;
A = 8'hAD; B = 8'h25; #100;
A = 8'hAD; B = 8'h26; #100;
A = 8'hAD; B = 8'h27; #100;
A = 8'hAD; B = 8'h28; #100;
A = 8'hAD; B = 8'h29; #100;
A = 8'hAD; B = 8'h2A; #100;
A = 8'hAD; B = 8'h2B; #100;
A = 8'hAD; B = 8'h2C; #100;
A = 8'hAD; B = 8'h2D; #100;
A = 8'hAD; B = 8'h2E; #100;
A = 8'hAD; B = 8'h2F; #100;
A = 8'hAD; B = 8'h30; #100;
A = 8'hAD; B = 8'h31; #100;
A = 8'hAD; B = 8'h32; #100;
A = 8'hAD; B = 8'h33; #100;
A = 8'hAD; B = 8'h34; #100;
A = 8'hAD; B = 8'h35; #100;
A = 8'hAD; B = 8'h36; #100;
A = 8'hAD; B = 8'h37; #100;
A = 8'hAD; B = 8'h38; #100;
A = 8'hAD; B = 8'h39; #100;
A = 8'hAD; B = 8'h3A; #100;
A = 8'hAD; B = 8'h3B; #100;
A = 8'hAD; B = 8'h3C; #100;
A = 8'hAD; B = 8'h3D; #100;
A = 8'hAD; B = 8'h3E; #100;
A = 8'hAD; B = 8'h3F; #100;
A = 8'hAD; B = 8'h40; #100;
A = 8'hAD; B = 8'h41; #100;
A = 8'hAD; B = 8'h42; #100;
A = 8'hAD; B = 8'h43; #100;
A = 8'hAD; B = 8'h44; #100;
A = 8'hAD; B = 8'h45; #100;
A = 8'hAD; B = 8'h46; #100;
A = 8'hAD; B = 8'h47; #100;
A = 8'hAD; B = 8'h48; #100;
A = 8'hAD; B = 8'h49; #100;
A = 8'hAD; B = 8'h4A; #100;
A = 8'hAD; B = 8'h4B; #100;
A = 8'hAD; B = 8'h4C; #100;
A = 8'hAD; B = 8'h4D; #100;
A = 8'hAD; B = 8'h4E; #100;
A = 8'hAD; B = 8'h4F; #100;
A = 8'hAD; B = 8'h50; #100;
A = 8'hAD; B = 8'h51; #100;
A = 8'hAD; B = 8'h52; #100;
A = 8'hAD; B = 8'h53; #100;
A = 8'hAD; B = 8'h54; #100;
A = 8'hAD; B = 8'h55; #100;
A = 8'hAD; B = 8'h56; #100;
A = 8'hAD; B = 8'h57; #100;
A = 8'hAD; B = 8'h58; #100;
A = 8'hAD; B = 8'h59; #100;
A = 8'hAD; B = 8'h5A; #100;
A = 8'hAD; B = 8'h5B; #100;
A = 8'hAD; B = 8'h5C; #100;
A = 8'hAD; B = 8'h5D; #100;
A = 8'hAD; B = 8'h5E; #100;
A = 8'hAD; B = 8'h5F; #100;
A = 8'hAD; B = 8'h60; #100;
A = 8'hAD; B = 8'h61; #100;
A = 8'hAD; B = 8'h62; #100;
A = 8'hAD; B = 8'h63; #100;
A = 8'hAD; B = 8'h64; #100;
A = 8'hAD; B = 8'h65; #100;
A = 8'hAD; B = 8'h66; #100;
A = 8'hAD; B = 8'h67; #100;
A = 8'hAD; B = 8'h68; #100;
A = 8'hAD; B = 8'h69; #100;
A = 8'hAD; B = 8'h6A; #100;
A = 8'hAD; B = 8'h6B; #100;
A = 8'hAD; B = 8'h6C; #100;
A = 8'hAD; B = 8'h6D; #100;
A = 8'hAD; B = 8'h6E; #100;
A = 8'hAD; B = 8'h6F; #100;
A = 8'hAD; B = 8'h70; #100;
A = 8'hAD; B = 8'h71; #100;
A = 8'hAD; B = 8'h72; #100;
A = 8'hAD; B = 8'h73; #100;
A = 8'hAD; B = 8'h74; #100;
A = 8'hAD; B = 8'h75; #100;
A = 8'hAD; B = 8'h76; #100;
A = 8'hAD; B = 8'h77; #100;
A = 8'hAD; B = 8'h78; #100;
A = 8'hAD; B = 8'h79; #100;
A = 8'hAD; B = 8'h7A; #100;
A = 8'hAD; B = 8'h7B; #100;
A = 8'hAD; B = 8'h7C; #100;
A = 8'hAD; B = 8'h7D; #100;
A = 8'hAD; B = 8'h7E; #100;
A = 8'hAD; B = 8'h7F; #100;
A = 8'hAD; B = 8'h80; #100;
A = 8'hAD; B = 8'h81; #100;
A = 8'hAD; B = 8'h82; #100;
A = 8'hAD; B = 8'h83; #100;
A = 8'hAD; B = 8'h84; #100;
A = 8'hAD; B = 8'h85; #100;
A = 8'hAD; B = 8'h86; #100;
A = 8'hAD; B = 8'h87; #100;
A = 8'hAD; B = 8'h88; #100;
A = 8'hAD; B = 8'h89; #100;
A = 8'hAD; B = 8'h8A; #100;
A = 8'hAD; B = 8'h8B; #100;
A = 8'hAD; B = 8'h8C; #100;
A = 8'hAD; B = 8'h8D; #100;
A = 8'hAD; B = 8'h8E; #100;
A = 8'hAD; B = 8'h8F; #100;
A = 8'hAD; B = 8'h90; #100;
A = 8'hAD; B = 8'h91; #100;
A = 8'hAD; B = 8'h92; #100;
A = 8'hAD; B = 8'h93; #100;
A = 8'hAD; B = 8'h94; #100;
A = 8'hAD; B = 8'h95; #100;
A = 8'hAD; B = 8'h96; #100;
A = 8'hAD; B = 8'h97; #100;
A = 8'hAD; B = 8'h98; #100;
A = 8'hAD; B = 8'h99; #100;
A = 8'hAD; B = 8'h9A; #100;
A = 8'hAD; B = 8'h9B; #100;
A = 8'hAD; B = 8'h9C; #100;
A = 8'hAD; B = 8'h9D; #100;
A = 8'hAD; B = 8'h9E; #100;
A = 8'hAD; B = 8'h9F; #100;
A = 8'hAD; B = 8'hA0; #100;
A = 8'hAD; B = 8'hA1; #100;
A = 8'hAD; B = 8'hA2; #100;
A = 8'hAD; B = 8'hA3; #100;
A = 8'hAD; B = 8'hA4; #100;
A = 8'hAD; B = 8'hA5; #100;
A = 8'hAD; B = 8'hA6; #100;
A = 8'hAD; B = 8'hA7; #100;
A = 8'hAD; B = 8'hA8; #100;
A = 8'hAD; B = 8'hA9; #100;
A = 8'hAD; B = 8'hAA; #100;
A = 8'hAD; B = 8'hAB; #100;
A = 8'hAD; B = 8'hAC; #100;
A = 8'hAD; B = 8'hAD; #100;
A = 8'hAD; B = 8'hAE; #100;
A = 8'hAD; B = 8'hAF; #100;
A = 8'hAD; B = 8'hB0; #100;
A = 8'hAD; B = 8'hB1; #100;
A = 8'hAD; B = 8'hB2; #100;
A = 8'hAD; B = 8'hB3; #100;
A = 8'hAD; B = 8'hB4; #100;
A = 8'hAD; B = 8'hB5; #100;
A = 8'hAD; B = 8'hB6; #100;
A = 8'hAD; B = 8'hB7; #100;
A = 8'hAD; B = 8'hB8; #100;
A = 8'hAD; B = 8'hB9; #100;
A = 8'hAD; B = 8'hBA; #100;
A = 8'hAD; B = 8'hBB; #100;
A = 8'hAD; B = 8'hBC; #100;
A = 8'hAD; B = 8'hBD; #100;
A = 8'hAD; B = 8'hBE; #100;
A = 8'hAD; B = 8'hBF; #100;
A = 8'hAD; B = 8'hC0; #100;
A = 8'hAD; B = 8'hC1; #100;
A = 8'hAD; B = 8'hC2; #100;
A = 8'hAD; B = 8'hC3; #100;
A = 8'hAD; B = 8'hC4; #100;
A = 8'hAD; B = 8'hC5; #100;
A = 8'hAD; B = 8'hC6; #100;
A = 8'hAD; B = 8'hC7; #100;
A = 8'hAD; B = 8'hC8; #100;
A = 8'hAD; B = 8'hC9; #100;
A = 8'hAD; B = 8'hCA; #100;
A = 8'hAD; B = 8'hCB; #100;
A = 8'hAD; B = 8'hCC; #100;
A = 8'hAD; B = 8'hCD; #100;
A = 8'hAD; B = 8'hCE; #100;
A = 8'hAD; B = 8'hCF; #100;
A = 8'hAD; B = 8'hD0; #100;
A = 8'hAD; B = 8'hD1; #100;
A = 8'hAD; B = 8'hD2; #100;
A = 8'hAD; B = 8'hD3; #100;
A = 8'hAD; B = 8'hD4; #100;
A = 8'hAD; B = 8'hD5; #100;
A = 8'hAD; B = 8'hD6; #100;
A = 8'hAD; B = 8'hD7; #100;
A = 8'hAD; B = 8'hD8; #100;
A = 8'hAD; B = 8'hD9; #100;
A = 8'hAD; B = 8'hDA; #100;
A = 8'hAD; B = 8'hDB; #100;
A = 8'hAD; B = 8'hDC; #100;
A = 8'hAD; B = 8'hDD; #100;
A = 8'hAD; B = 8'hDE; #100;
A = 8'hAD; B = 8'hDF; #100;
A = 8'hAD; B = 8'hE0; #100;
A = 8'hAD; B = 8'hE1; #100;
A = 8'hAD; B = 8'hE2; #100;
A = 8'hAD; B = 8'hE3; #100;
A = 8'hAD; B = 8'hE4; #100;
A = 8'hAD; B = 8'hE5; #100;
A = 8'hAD; B = 8'hE6; #100;
A = 8'hAD; B = 8'hE7; #100;
A = 8'hAD; B = 8'hE8; #100;
A = 8'hAD; B = 8'hE9; #100;
A = 8'hAD; B = 8'hEA; #100;
A = 8'hAD; B = 8'hEB; #100;
A = 8'hAD; B = 8'hEC; #100;
A = 8'hAD; B = 8'hED; #100;
A = 8'hAD; B = 8'hEE; #100;
A = 8'hAD; B = 8'hEF; #100;
A = 8'hAD; B = 8'hF0; #100;
A = 8'hAD; B = 8'hF1; #100;
A = 8'hAD; B = 8'hF2; #100;
A = 8'hAD; B = 8'hF3; #100;
A = 8'hAD; B = 8'hF4; #100;
A = 8'hAD; B = 8'hF5; #100;
A = 8'hAD; B = 8'hF6; #100;
A = 8'hAD; B = 8'hF7; #100;
A = 8'hAD; B = 8'hF8; #100;
A = 8'hAD; B = 8'hF9; #100;
A = 8'hAD; B = 8'hFA; #100;
A = 8'hAD; B = 8'hFB; #100;
A = 8'hAD; B = 8'hFC; #100;
A = 8'hAD; B = 8'hFD; #100;
A = 8'hAD; B = 8'hFE; #100;
A = 8'hAD; B = 8'hFF; #100;
A = 8'hAE; B = 8'h0; #100;
A = 8'hAE; B = 8'h1; #100;
A = 8'hAE; B = 8'h2; #100;
A = 8'hAE; B = 8'h3; #100;
A = 8'hAE; B = 8'h4; #100;
A = 8'hAE; B = 8'h5; #100;
A = 8'hAE; B = 8'h6; #100;
A = 8'hAE; B = 8'h7; #100;
A = 8'hAE; B = 8'h8; #100;
A = 8'hAE; B = 8'h9; #100;
A = 8'hAE; B = 8'hA; #100;
A = 8'hAE; B = 8'hB; #100;
A = 8'hAE; B = 8'hC; #100;
A = 8'hAE; B = 8'hD; #100;
A = 8'hAE; B = 8'hE; #100;
A = 8'hAE; B = 8'hF; #100;
A = 8'hAE; B = 8'h10; #100;
A = 8'hAE; B = 8'h11; #100;
A = 8'hAE; B = 8'h12; #100;
A = 8'hAE; B = 8'h13; #100;
A = 8'hAE; B = 8'h14; #100;
A = 8'hAE; B = 8'h15; #100;
A = 8'hAE; B = 8'h16; #100;
A = 8'hAE; B = 8'h17; #100;
A = 8'hAE; B = 8'h18; #100;
A = 8'hAE; B = 8'h19; #100;
A = 8'hAE; B = 8'h1A; #100;
A = 8'hAE; B = 8'h1B; #100;
A = 8'hAE; B = 8'h1C; #100;
A = 8'hAE; B = 8'h1D; #100;
A = 8'hAE; B = 8'h1E; #100;
A = 8'hAE; B = 8'h1F; #100;
A = 8'hAE; B = 8'h20; #100;
A = 8'hAE; B = 8'h21; #100;
A = 8'hAE; B = 8'h22; #100;
A = 8'hAE; B = 8'h23; #100;
A = 8'hAE; B = 8'h24; #100;
A = 8'hAE; B = 8'h25; #100;
A = 8'hAE; B = 8'h26; #100;
A = 8'hAE; B = 8'h27; #100;
A = 8'hAE; B = 8'h28; #100;
A = 8'hAE; B = 8'h29; #100;
A = 8'hAE; B = 8'h2A; #100;
A = 8'hAE; B = 8'h2B; #100;
A = 8'hAE; B = 8'h2C; #100;
A = 8'hAE; B = 8'h2D; #100;
A = 8'hAE; B = 8'h2E; #100;
A = 8'hAE; B = 8'h2F; #100;
A = 8'hAE; B = 8'h30; #100;
A = 8'hAE; B = 8'h31; #100;
A = 8'hAE; B = 8'h32; #100;
A = 8'hAE; B = 8'h33; #100;
A = 8'hAE; B = 8'h34; #100;
A = 8'hAE; B = 8'h35; #100;
A = 8'hAE; B = 8'h36; #100;
A = 8'hAE; B = 8'h37; #100;
A = 8'hAE; B = 8'h38; #100;
A = 8'hAE; B = 8'h39; #100;
A = 8'hAE; B = 8'h3A; #100;
A = 8'hAE; B = 8'h3B; #100;
A = 8'hAE; B = 8'h3C; #100;
A = 8'hAE; B = 8'h3D; #100;
A = 8'hAE; B = 8'h3E; #100;
A = 8'hAE; B = 8'h3F; #100;
A = 8'hAE; B = 8'h40; #100;
A = 8'hAE; B = 8'h41; #100;
A = 8'hAE; B = 8'h42; #100;
A = 8'hAE; B = 8'h43; #100;
A = 8'hAE; B = 8'h44; #100;
A = 8'hAE; B = 8'h45; #100;
A = 8'hAE; B = 8'h46; #100;
A = 8'hAE; B = 8'h47; #100;
A = 8'hAE; B = 8'h48; #100;
A = 8'hAE; B = 8'h49; #100;
A = 8'hAE; B = 8'h4A; #100;
A = 8'hAE; B = 8'h4B; #100;
A = 8'hAE; B = 8'h4C; #100;
A = 8'hAE; B = 8'h4D; #100;
A = 8'hAE; B = 8'h4E; #100;
A = 8'hAE; B = 8'h4F; #100;
A = 8'hAE; B = 8'h50; #100;
A = 8'hAE; B = 8'h51; #100;
A = 8'hAE; B = 8'h52; #100;
A = 8'hAE; B = 8'h53; #100;
A = 8'hAE; B = 8'h54; #100;
A = 8'hAE; B = 8'h55; #100;
A = 8'hAE; B = 8'h56; #100;
A = 8'hAE; B = 8'h57; #100;
A = 8'hAE; B = 8'h58; #100;
A = 8'hAE; B = 8'h59; #100;
A = 8'hAE; B = 8'h5A; #100;
A = 8'hAE; B = 8'h5B; #100;
A = 8'hAE; B = 8'h5C; #100;
A = 8'hAE; B = 8'h5D; #100;
A = 8'hAE; B = 8'h5E; #100;
A = 8'hAE; B = 8'h5F; #100;
A = 8'hAE; B = 8'h60; #100;
A = 8'hAE; B = 8'h61; #100;
A = 8'hAE; B = 8'h62; #100;
A = 8'hAE; B = 8'h63; #100;
A = 8'hAE; B = 8'h64; #100;
A = 8'hAE; B = 8'h65; #100;
A = 8'hAE; B = 8'h66; #100;
A = 8'hAE; B = 8'h67; #100;
A = 8'hAE; B = 8'h68; #100;
A = 8'hAE; B = 8'h69; #100;
A = 8'hAE; B = 8'h6A; #100;
A = 8'hAE; B = 8'h6B; #100;
A = 8'hAE; B = 8'h6C; #100;
A = 8'hAE; B = 8'h6D; #100;
A = 8'hAE; B = 8'h6E; #100;
A = 8'hAE; B = 8'h6F; #100;
A = 8'hAE; B = 8'h70; #100;
A = 8'hAE; B = 8'h71; #100;
A = 8'hAE; B = 8'h72; #100;
A = 8'hAE; B = 8'h73; #100;
A = 8'hAE; B = 8'h74; #100;
A = 8'hAE; B = 8'h75; #100;
A = 8'hAE; B = 8'h76; #100;
A = 8'hAE; B = 8'h77; #100;
A = 8'hAE; B = 8'h78; #100;
A = 8'hAE; B = 8'h79; #100;
A = 8'hAE; B = 8'h7A; #100;
A = 8'hAE; B = 8'h7B; #100;
A = 8'hAE; B = 8'h7C; #100;
A = 8'hAE; B = 8'h7D; #100;
A = 8'hAE; B = 8'h7E; #100;
A = 8'hAE; B = 8'h7F; #100;
A = 8'hAE; B = 8'h80; #100;
A = 8'hAE; B = 8'h81; #100;
A = 8'hAE; B = 8'h82; #100;
A = 8'hAE; B = 8'h83; #100;
A = 8'hAE; B = 8'h84; #100;
A = 8'hAE; B = 8'h85; #100;
A = 8'hAE; B = 8'h86; #100;
A = 8'hAE; B = 8'h87; #100;
A = 8'hAE; B = 8'h88; #100;
A = 8'hAE; B = 8'h89; #100;
A = 8'hAE; B = 8'h8A; #100;
A = 8'hAE; B = 8'h8B; #100;
A = 8'hAE; B = 8'h8C; #100;
A = 8'hAE; B = 8'h8D; #100;
A = 8'hAE; B = 8'h8E; #100;
A = 8'hAE; B = 8'h8F; #100;
A = 8'hAE; B = 8'h90; #100;
A = 8'hAE; B = 8'h91; #100;
A = 8'hAE; B = 8'h92; #100;
A = 8'hAE; B = 8'h93; #100;
A = 8'hAE; B = 8'h94; #100;
A = 8'hAE; B = 8'h95; #100;
A = 8'hAE; B = 8'h96; #100;
A = 8'hAE; B = 8'h97; #100;
A = 8'hAE; B = 8'h98; #100;
A = 8'hAE; B = 8'h99; #100;
A = 8'hAE; B = 8'h9A; #100;
A = 8'hAE; B = 8'h9B; #100;
A = 8'hAE; B = 8'h9C; #100;
A = 8'hAE; B = 8'h9D; #100;
A = 8'hAE; B = 8'h9E; #100;
A = 8'hAE; B = 8'h9F; #100;
A = 8'hAE; B = 8'hA0; #100;
A = 8'hAE; B = 8'hA1; #100;
A = 8'hAE; B = 8'hA2; #100;
A = 8'hAE; B = 8'hA3; #100;
A = 8'hAE; B = 8'hA4; #100;
A = 8'hAE; B = 8'hA5; #100;
A = 8'hAE; B = 8'hA6; #100;
A = 8'hAE; B = 8'hA7; #100;
A = 8'hAE; B = 8'hA8; #100;
A = 8'hAE; B = 8'hA9; #100;
A = 8'hAE; B = 8'hAA; #100;
A = 8'hAE; B = 8'hAB; #100;
A = 8'hAE; B = 8'hAC; #100;
A = 8'hAE; B = 8'hAD; #100;
A = 8'hAE; B = 8'hAE; #100;
A = 8'hAE; B = 8'hAF; #100;
A = 8'hAE; B = 8'hB0; #100;
A = 8'hAE; B = 8'hB1; #100;
A = 8'hAE; B = 8'hB2; #100;
A = 8'hAE; B = 8'hB3; #100;
A = 8'hAE; B = 8'hB4; #100;
A = 8'hAE; B = 8'hB5; #100;
A = 8'hAE; B = 8'hB6; #100;
A = 8'hAE; B = 8'hB7; #100;
A = 8'hAE; B = 8'hB8; #100;
A = 8'hAE; B = 8'hB9; #100;
A = 8'hAE; B = 8'hBA; #100;
A = 8'hAE; B = 8'hBB; #100;
A = 8'hAE; B = 8'hBC; #100;
A = 8'hAE; B = 8'hBD; #100;
A = 8'hAE; B = 8'hBE; #100;
A = 8'hAE; B = 8'hBF; #100;
A = 8'hAE; B = 8'hC0; #100;
A = 8'hAE; B = 8'hC1; #100;
A = 8'hAE; B = 8'hC2; #100;
A = 8'hAE; B = 8'hC3; #100;
A = 8'hAE; B = 8'hC4; #100;
A = 8'hAE; B = 8'hC5; #100;
A = 8'hAE; B = 8'hC6; #100;
A = 8'hAE; B = 8'hC7; #100;
A = 8'hAE; B = 8'hC8; #100;
A = 8'hAE; B = 8'hC9; #100;
A = 8'hAE; B = 8'hCA; #100;
A = 8'hAE; B = 8'hCB; #100;
A = 8'hAE; B = 8'hCC; #100;
A = 8'hAE; B = 8'hCD; #100;
A = 8'hAE; B = 8'hCE; #100;
A = 8'hAE; B = 8'hCF; #100;
A = 8'hAE; B = 8'hD0; #100;
A = 8'hAE; B = 8'hD1; #100;
A = 8'hAE; B = 8'hD2; #100;
A = 8'hAE; B = 8'hD3; #100;
A = 8'hAE; B = 8'hD4; #100;
A = 8'hAE; B = 8'hD5; #100;
A = 8'hAE; B = 8'hD6; #100;
A = 8'hAE; B = 8'hD7; #100;
A = 8'hAE; B = 8'hD8; #100;
A = 8'hAE; B = 8'hD9; #100;
A = 8'hAE; B = 8'hDA; #100;
A = 8'hAE; B = 8'hDB; #100;
A = 8'hAE; B = 8'hDC; #100;
A = 8'hAE; B = 8'hDD; #100;
A = 8'hAE; B = 8'hDE; #100;
A = 8'hAE; B = 8'hDF; #100;
A = 8'hAE; B = 8'hE0; #100;
A = 8'hAE; B = 8'hE1; #100;
A = 8'hAE; B = 8'hE2; #100;
A = 8'hAE; B = 8'hE3; #100;
A = 8'hAE; B = 8'hE4; #100;
A = 8'hAE; B = 8'hE5; #100;
A = 8'hAE; B = 8'hE6; #100;
A = 8'hAE; B = 8'hE7; #100;
A = 8'hAE; B = 8'hE8; #100;
A = 8'hAE; B = 8'hE9; #100;
A = 8'hAE; B = 8'hEA; #100;
A = 8'hAE; B = 8'hEB; #100;
A = 8'hAE; B = 8'hEC; #100;
A = 8'hAE; B = 8'hED; #100;
A = 8'hAE; B = 8'hEE; #100;
A = 8'hAE; B = 8'hEF; #100;
A = 8'hAE; B = 8'hF0; #100;
A = 8'hAE; B = 8'hF1; #100;
A = 8'hAE; B = 8'hF2; #100;
A = 8'hAE; B = 8'hF3; #100;
A = 8'hAE; B = 8'hF4; #100;
A = 8'hAE; B = 8'hF5; #100;
A = 8'hAE; B = 8'hF6; #100;
A = 8'hAE; B = 8'hF7; #100;
A = 8'hAE; B = 8'hF8; #100;
A = 8'hAE; B = 8'hF9; #100;
A = 8'hAE; B = 8'hFA; #100;
A = 8'hAE; B = 8'hFB; #100;
A = 8'hAE; B = 8'hFC; #100;
A = 8'hAE; B = 8'hFD; #100;
A = 8'hAE; B = 8'hFE; #100;
A = 8'hAE; B = 8'hFF; #100;
A = 8'hAF; B = 8'h0; #100;
A = 8'hAF; B = 8'h1; #100;
A = 8'hAF; B = 8'h2; #100;
A = 8'hAF; B = 8'h3; #100;
A = 8'hAF; B = 8'h4; #100;
A = 8'hAF; B = 8'h5; #100;
A = 8'hAF; B = 8'h6; #100;
A = 8'hAF; B = 8'h7; #100;
A = 8'hAF; B = 8'h8; #100;
A = 8'hAF; B = 8'h9; #100;
A = 8'hAF; B = 8'hA; #100;
A = 8'hAF; B = 8'hB; #100;
A = 8'hAF; B = 8'hC; #100;
A = 8'hAF; B = 8'hD; #100;
A = 8'hAF; B = 8'hE; #100;
A = 8'hAF; B = 8'hF; #100;
A = 8'hAF; B = 8'h10; #100;
A = 8'hAF; B = 8'h11; #100;
A = 8'hAF; B = 8'h12; #100;
A = 8'hAF; B = 8'h13; #100;
A = 8'hAF; B = 8'h14; #100;
A = 8'hAF; B = 8'h15; #100;
A = 8'hAF; B = 8'h16; #100;
A = 8'hAF; B = 8'h17; #100;
A = 8'hAF; B = 8'h18; #100;
A = 8'hAF; B = 8'h19; #100;
A = 8'hAF; B = 8'h1A; #100;
A = 8'hAF; B = 8'h1B; #100;
A = 8'hAF; B = 8'h1C; #100;
A = 8'hAF; B = 8'h1D; #100;
A = 8'hAF; B = 8'h1E; #100;
A = 8'hAF; B = 8'h1F; #100;
A = 8'hAF; B = 8'h20; #100;
A = 8'hAF; B = 8'h21; #100;
A = 8'hAF; B = 8'h22; #100;
A = 8'hAF; B = 8'h23; #100;
A = 8'hAF; B = 8'h24; #100;
A = 8'hAF; B = 8'h25; #100;
A = 8'hAF; B = 8'h26; #100;
A = 8'hAF; B = 8'h27; #100;
A = 8'hAF; B = 8'h28; #100;
A = 8'hAF; B = 8'h29; #100;
A = 8'hAF; B = 8'h2A; #100;
A = 8'hAF; B = 8'h2B; #100;
A = 8'hAF; B = 8'h2C; #100;
A = 8'hAF; B = 8'h2D; #100;
A = 8'hAF; B = 8'h2E; #100;
A = 8'hAF; B = 8'h2F; #100;
A = 8'hAF; B = 8'h30; #100;
A = 8'hAF; B = 8'h31; #100;
A = 8'hAF; B = 8'h32; #100;
A = 8'hAF; B = 8'h33; #100;
A = 8'hAF; B = 8'h34; #100;
A = 8'hAF; B = 8'h35; #100;
A = 8'hAF; B = 8'h36; #100;
A = 8'hAF; B = 8'h37; #100;
A = 8'hAF; B = 8'h38; #100;
A = 8'hAF; B = 8'h39; #100;
A = 8'hAF; B = 8'h3A; #100;
A = 8'hAF; B = 8'h3B; #100;
A = 8'hAF; B = 8'h3C; #100;
A = 8'hAF; B = 8'h3D; #100;
A = 8'hAF; B = 8'h3E; #100;
A = 8'hAF; B = 8'h3F; #100;
A = 8'hAF; B = 8'h40; #100;
A = 8'hAF; B = 8'h41; #100;
A = 8'hAF; B = 8'h42; #100;
A = 8'hAF; B = 8'h43; #100;
A = 8'hAF; B = 8'h44; #100;
A = 8'hAF; B = 8'h45; #100;
A = 8'hAF; B = 8'h46; #100;
A = 8'hAF; B = 8'h47; #100;
A = 8'hAF; B = 8'h48; #100;
A = 8'hAF; B = 8'h49; #100;
A = 8'hAF; B = 8'h4A; #100;
A = 8'hAF; B = 8'h4B; #100;
A = 8'hAF; B = 8'h4C; #100;
A = 8'hAF; B = 8'h4D; #100;
A = 8'hAF; B = 8'h4E; #100;
A = 8'hAF; B = 8'h4F; #100;
A = 8'hAF; B = 8'h50; #100;
A = 8'hAF; B = 8'h51; #100;
A = 8'hAF; B = 8'h52; #100;
A = 8'hAF; B = 8'h53; #100;
A = 8'hAF; B = 8'h54; #100;
A = 8'hAF; B = 8'h55; #100;
A = 8'hAF; B = 8'h56; #100;
A = 8'hAF; B = 8'h57; #100;
A = 8'hAF; B = 8'h58; #100;
A = 8'hAF; B = 8'h59; #100;
A = 8'hAF; B = 8'h5A; #100;
A = 8'hAF; B = 8'h5B; #100;
A = 8'hAF; B = 8'h5C; #100;
A = 8'hAF; B = 8'h5D; #100;
A = 8'hAF; B = 8'h5E; #100;
A = 8'hAF; B = 8'h5F; #100;
A = 8'hAF; B = 8'h60; #100;
A = 8'hAF; B = 8'h61; #100;
A = 8'hAF; B = 8'h62; #100;
A = 8'hAF; B = 8'h63; #100;
A = 8'hAF; B = 8'h64; #100;
A = 8'hAF; B = 8'h65; #100;
A = 8'hAF; B = 8'h66; #100;
A = 8'hAF; B = 8'h67; #100;
A = 8'hAF; B = 8'h68; #100;
A = 8'hAF; B = 8'h69; #100;
A = 8'hAF; B = 8'h6A; #100;
A = 8'hAF; B = 8'h6B; #100;
A = 8'hAF; B = 8'h6C; #100;
A = 8'hAF; B = 8'h6D; #100;
A = 8'hAF; B = 8'h6E; #100;
A = 8'hAF; B = 8'h6F; #100;
A = 8'hAF; B = 8'h70; #100;
A = 8'hAF; B = 8'h71; #100;
A = 8'hAF; B = 8'h72; #100;
A = 8'hAF; B = 8'h73; #100;
A = 8'hAF; B = 8'h74; #100;
A = 8'hAF; B = 8'h75; #100;
A = 8'hAF; B = 8'h76; #100;
A = 8'hAF; B = 8'h77; #100;
A = 8'hAF; B = 8'h78; #100;
A = 8'hAF; B = 8'h79; #100;
A = 8'hAF; B = 8'h7A; #100;
A = 8'hAF; B = 8'h7B; #100;
A = 8'hAF; B = 8'h7C; #100;
A = 8'hAF; B = 8'h7D; #100;
A = 8'hAF; B = 8'h7E; #100;
A = 8'hAF; B = 8'h7F; #100;
A = 8'hAF; B = 8'h80; #100;
A = 8'hAF; B = 8'h81; #100;
A = 8'hAF; B = 8'h82; #100;
A = 8'hAF; B = 8'h83; #100;
A = 8'hAF; B = 8'h84; #100;
A = 8'hAF; B = 8'h85; #100;
A = 8'hAF; B = 8'h86; #100;
A = 8'hAF; B = 8'h87; #100;
A = 8'hAF; B = 8'h88; #100;
A = 8'hAF; B = 8'h89; #100;
A = 8'hAF; B = 8'h8A; #100;
A = 8'hAF; B = 8'h8B; #100;
A = 8'hAF; B = 8'h8C; #100;
A = 8'hAF; B = 8'h8D; #100;
A = 8'hAF; B = 8'h8E; #100;
A = 8'hAF; B = 8'h8F; #100;
A = 8'hAF; B = 8'h90; #100;
A = 8'hAF; B = 8'h91; #100;
A = 8'hAF; B = 8'h92; #100;
A = 8'hAF; B = 8'h93; #100;
A = 8'hAF; B = 8'h94; #100;
A = 8'hAF; B = 8'h95; #100;
A = 8'hAF; B = 8'h96; #100;
A = 8'hAF; B = 8'h97; #100;
A = 8'hAF; B = 8'h98; #100;
A = 8'hAF; B = 8'h99; #100;
A = 8'hAF; B = 8'h9A; #100;
A = 8'hAF; B = 8'h9B; #100;
A = 8'hAF; B = 8'h9C; #100;
A = 8'hAF; B = 8'h9D; #100;
A = 8'hAF; B = 8'h9E; #100;
A = 8'hAF; B = 8'h9F; #100;
A = 8'hAF; B = 8'hA0; #100;
A = 8'hAF; B = 8'hA1; #100;
A = 8'hAF; B = 8'hA2; #100;
A = 8'hAF; B = 8'hA3; #100;
A = 8'hAF; B = 8'hA4; #100;
A = 8'hAF; B = 8'hA5; #100;
A = 8'hAF; B = 8'hA6; #100;
A = 8'hAF; B = 8'hA7; #100;
A = 8'hAF; B = 8'hA8; #100;
A = 8'hAF; B = 8'hA9; #100;
A = 8'hAF; B = 8'hAA; #100;
A = 8'hAF; B = 8'hAB; #100;
A = 8'hAF; B = 8'hAC; #100;
A = 8'hAF; B = 8'hAD; #100;
A = 8'hAF; B = 8'hAE; #100;
A = 8'hAF; B = 8'hAF; #100;
A = 8'hAF; B = 8'hB0; #100;
A = 8'hAF; B = 8'hB1; #100;
A = 8'hAF; B = 8'hB2; #100;
A = 8'hAF; B = 8'hB3; #100;
A = 8'hAF; B = 8'hB4; #100;
A = 8'hAF; B = 8'hB5; #100;
A = 8'hAF; B = 8'hB6; #100;
A = 8'hAF; B = 8'hB7; #100;
A = 8'hAF; B = 8'hB8; #100;
A = 8'hAF; B = 8'hB9; #100;
A = 8'hAF; B = 8'hBA; #100;
A = 8'hAF; B = 8'hBB; #100;
A = 8'hAF; B = 8'hBC; #100;
A = 8'hAF; B = 8'hBD; #100;
A = 8'hAF; B = 8'hBE; #100;
A = 8'hAF; B = 8'hBF; #100;
A = 8'hAF; B = 8'hC0; #100;
A = 8'hAF; B = 8'hC1; #100;
A = 8'hAF; B = 8'hC2; #100;
A = 8'hAF; B = 8'hC3; #100;
A = 8'hAF; B = 8'hC4; #100;
A = 8'hAF; B = 8'hC5; #100;
A = 8'hAF; B = 8'hC6; #100;
A = 8'hAF; B = 8'hC7; #100;
A = 8'hAF; B = 8'hC8; #100;
A = 8'hAF; B = 8'hC9; #100;
A = 8'hAF; B = 8'hCA; #100;
A = 8'hAF; B = 8'hCB; #100;
A = 8'hAF; B = 8'hCC; #100;
A = 8'hAF; B = 8'hCD; #100;
A = 8'hAF; B = 8'hCE; #100;
A = 8'hAF; B = 8'hCF; #100;
A = 8'hAF; B = 8'hD0; #100;
A = 8'hAF; B = 8'hD1; #100;
A = 8'hAF; B = 8'hD2; #100;
A = 8'hAF; B = 8'hD3; #100;
A = 8'hAF; B = 8'hD4; #100;
A = 8'hAF; B = 8'hD5; #100;
A = 8'hAF; B = 8'hD6; #100;
A = 8'hAF; B = 8'hD7; #100;
A = 8'hAF; B = 8'hD8; #100;
A = 8'hAF; B = 8'hD9; #100;
A = 8'hAF; B = 8'hDA; #100;
A = 8'hAF; B = 8'hDB; #100;
A = 8'hAF; B = 8'hDC; #100;
A = 8'hAF; B = 8'hDD; #100;
A = 8'hAF; B = 8'hDE; #100;
A = 8'hAF; B = 8'hDF; #100;
A = 8'hAF; B = 8'hE0; #100;
A = 8'hAF; B = 8'hE1; #100;
A = 8'hAF; B = 8'hE2; #100;
A = 8'hAF; B = 8'hE3; #100;
A = 8'hAF; B = 8'hE4; #100;
A = 8'hAF; B = 8'hE5; #100;
A = 8'hAF; B = 8'hE6; #100;
A = 8'hAF; B = 8'hE7; #100;
A = 8'hAF; B = 8'hE8; #100;
A = 8'hAF; B = 8'hE9; #100;
A = 8'hAF; B = 8'hEA; #100;
A = 8'hAF; B = 8'hEB; #100;
A = 8'hAF; B = 8'hEC; #100;
A = 8'hAF; B = 8'hED; #100;
A = 8'hAF; B = 8'hEE; #100;
A = 8'hAF; B = 8'hEF; #100;
A = 8'hAF; B = 8'hF0; #100;
A = 8'hAF; B = 8'hF1; #100;
A = 8'hAF; B = 8'hF2; #100;
A = 8'hAF; B = 8'hF3; #100;
A = 8'hAF; B = 8'hF4; #100;
A = 8'hAF; B = 8'hF5; #100;
A = 8'hAF; B = 8'hF6; #100;
A = 8'hAF; B = 8'hF7; #100;
A = 8'hAF; B = 8'hF8; #100;
A = 8'hAF; B = 8'hF9; #100;
A = 8'hAF; B = 8'hFA; #100;
A = 8'hAF; B = 8'hFB; #100;
A = 8'hAF; B = 8'hFC; #100;
A = 8'hAF; B = 8'hFD; #100;
A = 8'hAF; B = 8'hFE; #100;
A = 8'hAF; B = 8'hFF; #100;
A = 8'hB0; B = 8'h0; #100;
A = 8'hB0; B = 8'h1; #100;
A = 8'hB0; B = 8'h2; #100;
A = 8'hB0; B = 8'h3; #100;
A = 8'hB0; B = 8'h4; #100;
A = 8'hB0; B = 8'h5; #100;
A = 8'hB0; B = 8'h6; #100;
A = 8'hB0; B = 8'h7; #100;
A = 8'hB0; B = 8'h8; #100;
A = 8'hB0; B = 8'h9; #100;
A = 8'hB0; B = 8'hA; #100;
A = 8'hB0; B = 8'hB; #100;
A = 8'hB0; B = 8'hC; #100;
A = 8'hB0; B = 8'hD; #100;
A = 8'hB0; B = 8'hE; #100;
A = 8'hB0; B = 8'hF; #100;
A = 8'hB0; B = 8'h10; #100;
A = 8'hB0; B = 8'h11; #100;
A = 8'hB0; B = 8'h12; #100;
A = 8'hB0; B = 8'h13; #100;
A = 8'hB0; B = 8'h14; #100;
A = 8'hB0; B = 8'h15; #100;
A = 8'hB0; B = 8'h16; #100;
A = 8'hB0; B = 8'h17; #100;
A = 8'hB0; B = 8'h18; #100;
A = 8'hB0; B = 8'h19; #100;
A = 8'hB0; B = 8'h1A; #100;
A = 8'hB0; B = 8'h1B; #100;
A = 8'hB0; B = 8'h1C; #100;
A = 8'hB0; B = 8'h1D; #100;
A = 8'hB0; B = 8'h1E; #100;
A = 8'hB0; B = 8'h1F; #100;
A = 8'hB0; B = 8'h20; #100;
A = 8'hB0; B = 8'h21; #100;
A = 8'hB0; B = 8'h22; #100;
A = 8'hB0; B = 8'h23; #100;
A = 8'hB0; B = 8'h24; #100;
A = 8'hB0; B = 8'h25; #100;
A = 8'hB0; B = 8'h26; #100;
A = 8'hB0; B = 8'h27; #100;
A = 8'hB0; B = 8'h28; #100;
A = 8'hB0; B = 8'h29; #100;
A = 8'hB0; B = 8'h2A; #100;
A = 8'hB0; B = 8'h2B; #100;
A = 8'hB0; B = 8'h2C; #100;
A = 8'hB0; B = 8'h2D; #100;
A = 8'hB0; B = 8'h2E; #100;
A = 8'hB0; B = 8'h2F; #100;
A = 8'hB0; B = 8'h30; #100;
A = 8'hB0; B = 8'h31; #100;
A = 8'hB0; B = 8'h32; #100;
A = 8'hB0; B = 8'h33; #100;
A = 8'hB0; B = 8'h34; #100;
A = 8'hB0; B = 8'h35; #100;
A = 8'hB0; B = 8'h36; #100;
A = 8'hB0; B = 8'h37; #100;
A = 8'hB0; B = 8'h38; #100;
A = 8'hB0; B = 8'h39; #100;
A = 8'hB0; B = 8'h3A; #100;
A = 8'hB0; B = 8'h3B; #100;
A = 8'hB0; B = 8'h3C; #100;
A = 8'hB0; B = 8'h3D; #100;
A = 8'hB0; B = 8'h3E; #100;
A = 8'hB0; B = 8'h3F; #100;
A = 8'hB0; B = 8'h40; #100;
A = 8'hB0; B = 8'h41; #100;
A = 8'hB0; B = 8'h42; #100;
A = 8'hB0; B = 8'h43; #100;
A = 8'hB0; B = 8'h44; #100;
A = 8'hB0; B = 8'h45; #100;
A = 8'hB0; B = 8'h46; #100;
A = 8'hB0; B = 8'h47; #100;
A = 8'hB0; B = 8'h48; #100;
A = 8'hB0; B = 8'h49; #100;
A = 8'hB0; B = 8'h4A; #100;
A = 8'hB0; B = 8'h4B; #100;
A = 8'hB0; B = 8'h4C; #100;
A = 8'hB0; B = 8'h4D; #100;
A = 8'hB0; B = 8'h4E; #100;
A = 8'hB0; B = 8'h4F; #100;
A = 8'hB0; B = 8'h50; #100;
A = 8'hB0; B = 8'h51; #100;
A = 8'hB0; B = 8'h52; #100;
A = 8'hB0; B = 8'h53; #100;
A = 8'hB0; B = 8'h54; #100;
A = 8'hB0; B = 8'h55; #100;
A = 8'hB0; B = 8'h56; #100;
A = 8'hB0; B = 8'h57; #100;
A = 8'hB0; B = 8'h58; #100;
A = 8'hB0; B = 8'h59; #100;
A = 8'hB0; B = 8'h5A; #100;
A = 8'hB0; B = 8'h5B; #100;
A = 8'hB0; B = 8'h5C; #100;
A = 8'hB0; B = 8'h5D; #100;
A = 8'hB0; B = 8'h5E; #100;
A = 8'hB0; B = 8'h5F; #100;
A = 8'hB0; B = 8'h60; #100;
A = 8'hB0; B = 8'h61; #100;
A = 8'hB0; B = 8'h62; #100;
A = 8'hB0; B = 8'h63; #100;
A = 8'hB0; B = 8'h64; #100;
A = 8'hB0; B = 8'h65; #100;
A = 8'hB0; B = 8'h66; #100;
A = 8'hB0; B = 8'h67; #100;
A = 8'hB0; B = 8'h68; #100;
A = 8'hB0; B = 8'h69; #100;
A = 8'hB0; B = 8'h6A; #100;
A = 8'hB0; B = 8'h6B; #100;
A = 8'hB0; B = 8'h6C; #100;
A = 8'hB0; B = 8'h6D; #100;
A = 8'hB0; B = 8'h6E; #100;
A = 8'hB0; B = 8'h6F; #100;
A = 8'hB0; B = 8'h70; #100;
A = 8'hB0; B = 8'h71; #100;
A = 8'hB0; B = 8'h72; #100;
A = 8'hB0; B = 8'h73; #100;
A = 8'hB0; B = 8'h74; #100;
A = 8'hB0; B = 8'h75; #100;
A = 8'hB0; B = 8'h76; #100;
A = 8'hB0; B = 8'h77; #100;
A = 8'hB0; B = 8'h78; #100;
A = 8'hB0; B = 8'h79; #100;
A = 8'hB0; B = 8'h7A; #100;
A = 8'hB0; B = 8'h7B; #100;
A = 8'hB0; B = 8'h7C; #100;
A = 8'hB0; B = 8'h7D; #100;
A = 8'hB0; B = 8'h7E; #100;
A = 8'hB0; B = 8'h7F; #100;
A = 8'hB0; B = 8'h80; #100;
A = 8'hB0; B = 8'h81; #100;
A = 8'hB0; B = 8'h82; #100;
A = 8'hB0; B = 8'h83; #100;
A = 8'hB0; B = 8'h84; #100;
A = 8'hB0; B = 8'h85; #100;
A = 8'hB0; B = 8'h86; #100;
A = 8'hB0; B = 8'h87; #100;
A = 8'hB0; B = 8'h88; #100;
A = 8'hB0; B = 8'h89; #100;
A = 8'hB0; B = 8'h8A; #100;
A = 8'hB0; B = 8'h8B; #100;
A = 8'hB0; B = 8'h8C; #100;
A = 8'hB0; B = 8'h8D; #100;
A = 8'hB0; B = 8'h8E; #100;
A = 8'hB0; B = 8'h8F; #100;
A = 8'hB0; B = 8'h90; #100;
A = 8'hB0; B = 8'h91; #100;
A = 8'hB0; B = 8'h92; #100;
A = 8'hB0; B = 8'h93; #100;
A = 8'hB0; B = 8'h94; #100;
A = 8'hB0; B = 8'h95; #100;
A = 8'hB0; B = 8'h96; #100;
A = 8'hB0; B = 8'h97; #100;
A = 8'hB0; B = 8'h98; #100;
A = 8'hB0; B = 8'h99; #100;
A = 8'hB0; B = 8'h9A; #100;
A = 8'hB0; B = 8'h9B; #100;
A = 8'hB0; B = 8'h9C; #100;
A = 8'hB0; B = 8'h9D; #100;
A = 8'hB0; B = 8'h9E; #100;
A = 8'hB0; B = 8'h9F; #100;
A = 8'hB0; B = 8'hA0; #100;
A = 8'hB0; B = 8'hA1; #100;
A = 8'hB0; B = 8'hA2; #100;
A = 8'hB0; B = 8'hA3; #100;
A = 8'hB0; B = 8'hA4; #100;
A = 8'hB0; B = 8'hA5; #100;
A = 8'hB0; B = 8'hA6; #100;
A = 8'hB0; B = 8'hA7; #100;
A = 8'hB0; B = 8'hA8; #100;
A = 8'hB0; B = 8'hA9; #100;
A = 8'hB0; B = 8'hAA; #100;
A = 8'hB0; B = 8'hAB; #100;
A = 8'hB0; B = 8'hAC; #100;
A = 8'hB0; B = 8'hAD; #100;
A = 8'hB0; B = 8'hAE; #100;
A = 8'hB0; B = 8'hAF; #100;
A = 8'hB0; B = 8'hB0; #100;
A = 8'hB0; B = 8'hB1; #100;
A = 8'hB0; B = 8'hB2; #100;
A = 8'hB0; B = 8'hB3; #100;
A = 8'hB0; B = 8'hB4; #100;
A = 8'hB0; B = 8'hB5; #100;
A = 8'hB0; B = 8'hB6; #100;
A = 8'hB0; B = 8'hB7; #100;
A = 8'hB0; B = 8'hB8; #100;
A = 8'hB0; B = 8'hB9; #100;
A = 8'hB0; B = 8'hBA; #100;
A = 8'hB0; B = 8'hBB; #100;
A = 8'hB0; B = 8'hBC; #100;
A = 8'hB0; B = 8'hBD; #100;
A = 8'hB0; B = 8'hBE; #100;
A = 8'hB0; B = 8'hBF; #100;
A = 8'hB0; B = 8'hC0; #100;
A = 8'hB0; B = 8'hC1; #100;
A = 8'hB0; B = 8'hC2; #100;
A = 8'hB0; B = 8'hC3; #100;
A = 8'hB0; B = 8'hC4; #100;
A = 8'hB0; B = 8'hC5; #100;
A = 8'hB0; B = 8'hC6; #100;
A = 8'hB0; B = 8'hC7; #100;
A = 8'hB0; B = 8'hC8; #100;
A = 8'hB0; B = 8'hC9; #100;
A = 8'hB0; B = 8'hCA; #100;
A = 8'hB0; B = 8'hCB; #100;
A = 8'hB0; B = 8'hCC; #100;
A = 8'hB0; B = 8'hCD; #100;
A = 8'hB0; B = 8'hCE; #100;
A = 8'hB0; B = 8'hCF; #100;
A = 8'hB0; B = 8'hD0; #100;
A = 8'hB0; B = 8'hD1; #100;
A = 8'hB0; B = 8'hD2; #100;
A = 8'hB0; B = 8'hD3; #100;
A = 8'hB0; B = 8'hD4; #100;
A = 8'hB0; B = 8'hD5; #100;
A = 8'hB0; B = 8'hD6; #100;
A = 8'hB0; B = 8'hD7; #100;
A = 8'hB0; B = 8'hD8; #100;
A = 8'hB0; B = 8'hD9; #100;
A = 8'hB0; B = 8'hDA; #100;
A = 8'hB0; B = 8'hDB; #100;
A = 8'hB0; B = 8'hDC; #100;
A = 8'hB0; B = 8'hDD; #100;
A = 8'hB0; B = 8'hDE; #100;
A = 8'hB0; B = 8'hDF; #100;
A = 8'hB0; B = 8'hE0; #100;
A = 8'hB0; B = 8'hE1; #100;
A = 8'hB0; B = 8'hE2; #100;
A = 8'hB0; B = 8'hE3; #100;
A = 8'hB0; B = 8'hE4; #100;
A = 8'hB0; B = 8'hE5; #100;
A = 8'hB0; B = 8'hE6; #100;
A = 8'hB0; B = 8'hE7; #100;
A = 8'hB0; B = 8'hE8; #100;
A = 8'hB0; B = 8'hE9; #100;
A = 8'hB0; B = 8'hEA; #100;
A = 8'hB0; B = 8'hEB; #100;
A = 8'hB0; B = 8'hEC; #100;
A = 8'hB0; B = 8'hED; #100;
A = 8'hB0; B = 8'hEE; #100;
A = 8'hB0; B = 8'hEF; #100;
A = 8'hB0; B = 8'hF0; #100;
A = 8'hB0; B = 8'hF1; #100;
A = 8'hB0; B = 8'hF2; #100;
A = 8'hB0; B = 8'hF3; #100;
A = 8'hB0; B = 8'hF4; #100;
A = 8'hB0; B = 8'hF5; #100;
A = 8'hB0; B = 8'hF6; #100;
A = 8'hB0; B = 8'hF7; #100;
A = 8'hB0; B = 8'hF8; #100;
A = 8'hB0; B = 8'hF9; #100;
A = 8'hB0; B = 8'hFA; #100;
A = 8'hB0; B = 8'hFB; #100;
A = 8'hB0; B = 8'hFC; #100;
A = 8'hB0; B = 8'hFD; #100;
A = 8'hB0; B = 8'hFE; #100;
A = 8'hB0; B = 8'hFF; #100;
A = 8'hB1; B = 8'h0; #100;
A = 8'hB1; B = 8'h1; #100;
A = 8'hB1; B = 8'h2; #100;
A = 8'hB1; B = 8'h3; #100;
A = 8'hB1; B = 8'h4; #100;
A = 8'hB1; B = 8'h5; #100;
A = 8'hB1; B = 8'h6; #100;
A = 8'hB1; B = 8'h7; #100;
A = 8'hB1; B = 8'h8; #100;
A = 8'hB1; B = 8'h9; #100;
A = 8'hB1; B = 8'hA; #100;
A = 8'hB1; B = 8'hB; #100;
A = 8'hB1; B = 8'hC; #100;
A = 8'hB1; B = 8'hD; #100;
A = 8'hB1; B = 8'hE; #100;
A = 8'hB1; B = 8'hF; #100;
A = 8'hB1; B = 8'h10; #100;
A = 8'hB1; B = 8'h11; #100;
A = 8'hB1; B = 8'h12; #100;
A = 8'hB1; B = 8'h13; #100;
A = 8'hB1; B = 8'h14; #100;
A = 8'hB1; B = 8'h15; #100;
A = 8'hB1; B = 8'h16; #100;
A = 8'hB1; B = 8'h17; #100;
A = 8'hB1; B = 8'h18; #100;
A = 8'hB1; B = 8'h19; #100;
A = 8'hB1; B = 8'h1A; #100;
A = 8'hB1; B = 8'h1B; #100;
A = 8'hB1; B = 8'h1C; #100;
A = 8'hB1; B = 8'h1D; #100;
A = 8'hB1; B = 8'h1E; #100;
A = 8'hB1; B = 8'h1F; #100;
A = 8'hB1; B = 8'h20; #100;
A = 8'hB1; B = 8'h21; #100;
A = 8'hB1; B = 8'h22; #100;
A = 8'hB1; B = 8'h23; #100;
A = 8'hB1; B = 8'h24; #100;
A = 8'hB1; B = 8'h25; #100;
A = 8'hB1; B = 8'h26; #100;
A = 8'hB1; B = 8'h27; #100;
A = 8'hB1; B = 8'h28; #100;
A = 8'hB1; B = 8'h29; #100;
A = 8'hB1; B = 8'h2A; #100;
A = 8'hB1; B = 8'h2B; #100;
A = 8'hB1; B = 8'h2C; #100;
A = 8'hB1; B = 8'h2D; #100;
A = 8'hB1; B = 8'h2E; #100;
A = 8'hB1; B = 8'h2F; #100;
A = 8'hB1; B = 8'h30; #100;
A = 8'hB1; B = 8'h31; #100;
A = 8'hB1; B = 8'h32; #100;
A = 8'hB1; B = 8'h33; #100;
A = 8'hB1; B = 8'h34; #100;
A = 8'hB1; B = 8'h35; #100;
A = 8'hB1; B = 8'h36; #100;
A = 8'hB1; B = 8'h37; #100;
A = 8'hB1; B = 8'h38; #100;
A = 8'hB1; B = 8'h39; #100;
A = 8'hB1; B = 8'h3A; #100;
A = 8'hB1; B = 8'h3B; #100;
A = 8'hB1; B = 8'h3C; #100;
A = 8'hB1; B = 8'h3D; #100;
A = 8'hB1; B = 8'h3E; #100;
A = 8'hB1; B = 8'h3F; #100;
A = 8'hB1; B = 8'h40; #100;
A = 8'hB1; B = 8'h41; #100;
A = 8'hB1; B = 8'h42; #100;
A = 8'hB1; B = 8'h43; #100;
A = 8'hB1; B = 8'h44; #100;
A = 8'hB1; B = 8'h45; #100;
A = 8'hB1; B = 8'h46; #100;
A = 8'hB1; B = 8'h47; #100;
A = 8'hB1; B = 8'h48; #100;
A = 8'hB1; B = 8'h49; #100;
A = 8'hB1; B = 8'h4A; #100;
A = 8'hB1; B = 8'h4B; #100;
A = 8'hB1; B = 8'h4C; #100;
A = 8'hB1; B = 8'h4D; #100;
A = 8'hB1; B = 8'h4E; #100;
A = 8'hB1; B = 8'h4F; #100;
A = 8'hB1; B = 8'h50; #100;
A = 8'hB1; B = 8'h51; #100;
A = 8'hB1; B = 8'h52; #100;
A = 8'hB1; B = 8'h53; #100;
A = 8'hB1; B = 8'h54; #100;
A = 8'hB1; B = 8'h55; #100;
A = 8'hB1; B = 8'h56; #100;
A = 8'hB1; B = 8'h57; #100;
A = 8'hB1; B = 8'h58; #100;
A = 8'hB1; B = 8'h59; #100;
A = 8'hB1; B = 8'h5A; #100;
A = 8'hB1; B = 8'h5B; #100;
A = 8'hB1; B = 8'h5C; #100;
A = 8'hB1; B = 8'h5D; #100;
A = 8'hB1; B = 8'h5E; #100;
A = 8'hB1; B = 8'h5F; #100;
A = 8'hB1; B = 8'h60; #100;
A = 8'hB1; B = 8'h61; #100;
A = 8'hB1; B = 8'h62; #100;
A = 8'hB1; B = 8'h63; #100;
A = 8'hB1; B = 8'h64; #100;
A = 8'hB1; B = 8'h65; #100;
A = 8'hB1; B = 8'h66; #100;
A = 8'hB1; B = 8'h67; #100;
A = 8'hB1; B = 8'h68; #100;
A = 8'hB1; B = 8'h69; #100;
A = 8'hB1; B = 8'h6A; #100;
A = 8'hB1; B = 8'h6B; #100;
A = 8'hB1; B = 8'h6C; #100;
A = 8'hB1; B = 8'h6D; #100;
A = 8'hB1; B = 8'h6E; #100;
A = 8'hB1; B = 8'h6F; #100;
A = 8'hB1; B = 8'h70; #100;
A = 8'hB1; B = 8'h71; #100;
A = 8'hB1; B = 8'h72; #100;
A = 8'hB1; B = 8'h73; #100;
A = 8'hB1; B = 8'h74; #100;
A = 8'hB1; B = 8'h75; #100;
A = 8'hB1; B = 8'h76; #100;
A = 8'hB1; B = 8'h77; #100;
A = 8'hB1; B = 8'h78; #100;
A = 8'hB1; B = 8'h79; #100;
A = 8'hB1; B = 8'h7A; #100;
A = 8'hB1; B = 8'h7B; #100;
A = 8'hB1; B = 8'h7C; #100;
A = 8'hB1; B = 8'h7D; #100;
A = 8'hB1; B = 8'h7E; #100;
A = 8'hB1; B = 8'h7F; #100;
A = 8'hB1; B = 8'h80; #100;
A = 8'hB1; B = 8'h81; #100;
A = 8'hB1; B = 8'h82; #100;
A = 8'hB1; B = 8'h83; #100;
A = 8'hB1; B = 8'h84; #100;
A = 8'hB1; B = 8'h85; #100;
A = 8'hB1; B = 8'h86; #100;
A = 8'hB1; B = 8'h87; #100;
A = 8'hB1; B = 8'h88; #100;
A = 8'hB1; B = 8'h89; #100;
A = 8'hB1; B = 8'h8A; #100;
A = 8'hB1; B = 8'h8B; #100;
A = 8'hB1; B = 8'h8C; #100;
A = 8'hB1; B = 8'h8D; #100;
A = 8'hB1; B = 8'h8E; #100;
A = 8'hB1; B = 8'h8F; #100;
A = 8'hB1; B = 8'h90; #100;
A = 8'hB1; B = 8'h91; #100;
A = 8'hB1; B = 8'h92; #100;
A = 8'hB1; B = 8'h93; #100;
A = 8'hB1; B = 8'h94; #100;
A = 8'hB1; B = 8'h95; #100;
A = 8'hB1; B = 8'h96; #100;
A = 8'hB1; B = 8'h97; #100;
A = 8'hB1; B = 8'h98; #100;
A = 8'hB1; B = 8'h99; #100;
A = 8'hB1; B = 8'h9A; #100;
A = 8'hB1; B = 8'h9B; #100;
A = 8'hB1; B = 8'h9C; #100;
A = 8'hB1; B = 8'h9D; #100;
A = 8'hB1; B = 8'h9E; #100;
A = 8'hB1; B = 8'h9F; #100;
A = 8'hB1; B = 8'hA0; #100;
A = 8'hB1; B = 8'hA1; #100;
A = 8'hB1; B = 8'hA2; #100;
A = 8'hB1; B = 8'hA3; #100;
A = 8'hB1; B = 8'hA4; #100;
A = 8'hB1; B = 8'hA5; #100;
A = 8'hB1; B = 8'hA6; #100;
A = 8'hB1; B = 8'hA7; #100;
A = 8'hB1; B = 8'hA8; #100;
A = 8'hB1; B = 8'hA9; #100;
A = 8'hB1; B = 8'hAA; #100;
A = 8'hB1; B = 8'hAB; #100;
A = 8'hB1; B = 8'hAC; #100;
A = 8'hB1; B = 8'hAD; #100;
A = 8'hB1; B = 8'hAE; #100;
A = 8'hB1; B = 8'hAF; #100;
A = 8'hB1; B = 8'hB0; #100;
A = 8'hB1; B = 8'hB1; #100;
A = 8'hB1; B = 8'hB2; #100;
A = 8'hB1; B = 8'hB3; #100;
A = 8'hB1; B = 8'hB4; #100;
A = 8'hB1; B = 8'hB5; #100;
A = 8'hB1; B = 8'hB6; #100;
A = 8'hB1; B = 8'hB7; #100;
A = 8'hB1; B = 8'hB8; #100;
A = 8'hB1; B = 8'hB9; #100;
A = 8'hB1; B = 8'hBA; #100;
A = 8'hB1; B = 8'hBB; #100;
A = 8'hB1; B = 8'hBC; #100;
A = 8'hB1; B = 8'hBD; #100;
A = 8'hB1; B = 8'hBE; #100;
A = 8'hB1; B = 8'hBF; #100;
A = 8'hB1; B = 8'hC0; #100;
A = 8'hB1; B = 8'hC1; #100;
A = 8'hB1; B = 8'hC2; #100;
A = 8'hB1; B = 8'hC3; #100;
A = 8'hB1; B = 8'hC4; #100;
A = 8'hB1; B = 8'hC5; #100;
A = 8'hB1; B = 8'hC6; #100;
A = 8'hB1; B = 8'hC7; #100;
A = 8'hB1; B = 8'hC8; #100;
A = 8'hB1; B = 8'hC9; #100;
A = 8'hB1; B = 8'hCA; #100;
A = 8'hB1; B = 8'hCB; #100;
A = 8'hB1; B = 8'hCC; #100;
A = 8'hB1; B = 8'hCD; #100;
A = 8'hB1; B = 8'hCE; #100;
A = 8'hB1; B = 8'hCF; #100;
A = 8'hB1; B = 8'hD0; #100;
A = 8'hB1; B = 8'hD1; #100;
A = 8'hB1; B = 8'hD2; #100;
A = 8'hB1; B = 8'hD3; #100;
A = 8'hB1; B = 8'hD4; #100;
A = 8'hB1; B = 8'hD5; #100;
A = 8'hB1; B = 8'hD6; #100;
A = 8'hB1; B = 8'hD7; #100;
A = 8'hB1; B = 8'hD8; #100;
A = 8'hB1; B = 8'hD9; #100;
A = 8'hB1; B = 8'hDA; #100;
A = 8'hB1; B = 8'hDB; #100;
A = 8'hB1; B = 8'hDC; #100;
A = 8'hB1; B = 8'hDD; #100;
A = 8'hB1; B = 8'hDE; #100;
A = 8'hB1; B = 8'hDF; #100;
A = 8'hB1; B = 8'hE0; #100;
A = 8'hB1; B = 8'hE1; #100;
A = 8'hB1; B = 8'hE2; #100;
A = 8'hB1; B = 8'hE3; #100;
A = 8'hB1; B = 8'hE4; #100;
A = 8'hB1; B = 8'hE5; #100;
A = 8'hB1; B = 8'hE6; #100;
A = 8'hB1; B = 8'hE7; #100;
A = 8'hB1; B = 8'hE8; #100;
A = 8'hB1; B = 8'hE9; #100;
A = 8'hB1; B = 8'hEA; #100;
A = 8'hB1; B = 8'hEB; #100;
A = 8'hB1; B = 8'hEC; #100;
A = 8'hB1; B = 8'hED; #100;
A = 8'hB1; B = 8'hEE; #100;
A = 8'hB1; B = 8'hEF; #100;
A = 8'hB1; B = 8'hF0; #100;
A = 8'hB1; B = 8'hF1; #100;
A = 8'hB1; B = 8'hF2; #100;
A = 8'hB1; B = 8'hF3; #100;
A = 8'hB1; B = 8'hF4; #100;
A = 8'hB1; B = 8'hF5; #100;
A = 8'hB1; B = 8'hF6; #100;
A = 8'hB1; B = 8'hF7; #100;
A = 8'hB1; B = 8'hF8; #100;
A = 8'hB1; B = 8'hF9; #100;
A = 8'hB1; B = 8'hFA; #100;
A = 8'hB1; B = 8'hFB; #100;
A = 8'hB1; B = 8'hFC; #100;
A = 8'hB1; B = 8'hFD; #100;
A = 8'hB1; B = 8'hFE; #100;
A = 8'hB1; B = 8'hFF; #100;
A = 8'hB2; B = 8'h0; #100;
A = 8'hB2; B = 8'h1; #100;
A = 8'hB2; B = 8'h2; #100;
A = 8'hB2; B = 8'h3; #100;
A = 8'hB2; B = 8'h4; #100;
A = 8'hB2; B = 8'h5; #100;
A = 8'hB2; B = 8'h6; #100;
A = 8'hB2; B = 8'h7; #100;
A = 8'hB2; B = 8'h8; #100;
A = 8'hB2; B = 8'h9; #100;
A = 8'hB2; B = 8'hA; #100;
A = 8'hB2; B = 8'hB; #100;
A = 8'hB2; B = 8'hC; #100;
A = 8'hB2; B = 8'hD; #100;
A = 8'hB2; B = 8'hE; #100;
A = 8'hB2; B = 8'hF; #100;
A = 8'hB2; B = 8'h10; #100;
A = 8'hB2; B = 8'h11; #100;
A = 8'hB2; B = 8'h12; #100;
A = 8'hB2; B = 8'h13; #100;
A = 8'hB2; B = 8'h14; #100;
A = 8'hB2; B = 8'h15; #100;
A = 8'hB2; B = 8'h16; #100;
A = 8'hB2; B = 8'h17; #100;
A = 8'hB2; B = 8'h18; #100;
A = 8'hB2; B = 8'h19; #100;
A = 8'hB2; B = 8'h1A; #100;
A = 8'hB2; B = 8'h1B; #100;
A = 8'hB2; B = 8'h1C; #100;
A = 8'hB2; B = 8'h1D; #100;
A = 8'hB2; B = 8'h1E; #100;
A = 8'hB2; B = 8'h1F; #100;
A = 8'hB2; B = 8'h20; #100;
A = 8'hB2; B = 8'h21; #100;
A = 8'hB2; B = 8'h22; #100;
A = 8'hB2; B = 8'h23; #100;
A = 8'hB2; B = 8'h24; #100;
A = 8'hB2; B = 8'h25; #100;
A = 8'hB2; B = 8'h26; #100;
A = 8'hB2; B = 8'h27; #100;
A = 8'hB2; B = 8'h28; #100;
A = 8'hB2; B = 8'h29; #100;
A = 8'hB2; B = 8'h2A; #100;
A = 8'hB2; B = 8'h2B; #100;
A = 8'hB2; B = 8'h2C; #100;
A = 8'hB2; B = 8'h2D; #100;
A = 8'hB2; B = 8'h2E; #100;
A = 8'hB2; B = 8'h2F; #100;
A = 8'hB2; B = 8'h30; #100;
A = 8'hB2; B = 8'h31; #100;
A = 8'hB2; B = 8'h32; #100;
A = 8'hB2; B = 8'h33; #100;
A = 8'hB2; B = 8'h34; #100;
A = 8'hB2; B = 8'h35; #100;
A = 8'hB2; B = 8'h36; #100;
A = 8'hB2; B = 8'h37; #100;
A = 8'hB2; B = 8'h38; #100;
A = 8'hB2; B = 8'h39; #100;
A = 8'hB2; B = 8'h3A; #100;
A = 8'hB2; B = 8'h3B; #100;
A = 8'hB2; B = 8'h3C; #100;
A = 8'hB2; B = 8'h3D; #100;
A = 8'hB2; B = 8'h3E; #100;
A = 8'hB2; B = 8'h3F; #100;
A = 8'hB2; B = 8'h40; #100;
A = 8'hB2; B = 8'h41; #100;
A = 8'hB2; B = 8'h42; #100;
A = 8'hB2; B = 8'h43; #100;
A = 8'hB2; B = 8'h44; #100;
A = 8'hB2; B = 8'h45; #100;
A = 8'hB2; B = 8'h46; #100;
A = 8'hB2; B = 8'h47; #100;
A = 8'hB2; B = 8'h48; #100;
A = 8'hB2; B = 8'h49; #100;
A = 8'hB2; B = 8'h4A; #100;
A = 8'hB2; B = 8'h4B; #100;
A = 8'hB2; B = 8'h4C; #100;
A = 8'hB2; B = 8'h4D; #100;
A = 8'hB2; B = 8'h4E; #100;
A = 8'hB2; B = 8'h4F; #100;
A = 8'hB2; B = 8'h50; #100;
A = 8'hB2; B = 8'h51; #100;
A = 8'hB2; B = 8'h52; #100;
A = 8'hB2; B = 8'h53; #100;
A = 8'hB2; B = 8'h54; #100;
A = 8'hB2; B = 8'h55; #100;
A = 8'hB2; B = 8'h56; #100;
A = 8'hB2; B = 8'h57; #100;
A = 8'hB2; B = 8'h58; #100;
A = 8'hB2; B = 8'h59; #100;
A = 8'hB2; B = 8'h5A; #100;
A = 8'hB2; B = 8'h5B; #100;
A = 8'hB2; B = 8'h5C; #100;
A = 8'hB2; B = 8'h5D; #100;
A = 8'hB2; B = 8'h5E; #100;
A = 8'hB2; B = 8'h5F; #100;
A = 8'hB2; B = 8'h60; #100;
A = 8'hB2; B = 8'h61; #100;
A = 8'hB2; B = 8'h62; #100;
A = 8'hB2; B = 8'h63; #100;
A = 8'hB2; B = 8'h64; #100;
A = 8'hB2; B = 8'h65; #100;
A = 8'hB2; B = 8'h66; #100;
A = 8'hB2; B = 8'h67; #100;
A = 8'hB2; B = 8'h68; #100;
A = 8'hB2; B = 8'h69; #100;
A = 8'hB2; B = 8'h6A; #100;
A = 8'hB2; B = 8'h6B; #100;
A = 8'hB2; B = 8'h6C; #100;
A = 8'hB2; B = 8'h6D; #100;
A = 8'hB2; B = 8'h6E; #100;
A = 8'hB2; B = 8'h6F; #100;
A = 8'hB2; B = 8'h70; #100;
A = 8'hB2; B = 8'h71; #100;
A = 8'hB2; B = 8'h72; #100;
A = 8'hB2; B = 8'h73; #100;
A = 8'hB2; B = 8'h74; #100;
A = 8'hB2; B = 8'h75; #100;
A = 8'hB2; B = 8'h76; #100;
A = 8'hB2; B = 8'h77; #100;
A = 8'hB2; B = 8'h78; #100;
A = 8'hB2; B = 8'h79; #100;
A = 8'hB2; B = 8'h7A; #100;
A = 8'hB2; B = 8'h7B; #100;
A = 8'hB2; B = 8'h7C; #100;
A = 8'hB2; B = 8'h7D; #100;
A = 8'hB2; B = 8'h7E; #100;
A = 8'hB2; B = 8'h7F; #100;
A = 8'hB2; B = 8'h80; #100;
A = 8'hB2; B = 8'h81; #100;
A = 8'hB2; B = 8'h82; #100;
A = 8'hB2; B = 8'h83; #100;
A = 8'hB2; B = 8'h84; #100;
A = 8'hB2; B = 8'h85; #100;
A = 8'hB2; B = 8'h86; #100;
A = 8'hB2; B = 8'h87; #100;
A = 8'hB2; B = 8'h88; #100;
A = 8'hB2; B = 8'h89; #100;
A = 8'hB2; B = 8'h8A; #100;
A = 8'hB2; B = 8'h8B; #100;
A = 8'hB2; B = 8'h8C; #100;
A = 8'hB2; B = 8'h8D; #100;
A = 8'hB2; B = 8'h8E; #100;
A = 8'hB2; B = 8'h8F; #100;
A = 8'hB2; B = 8'h90; #100;
A = 8'hB2; B = 8'h91; #100;
A = 8'hB2; B = 8'h92; #100;
A = 8'hB2; B = 8'h93; #100;
A = 8'hB2; B = 8'h94; #100;
A = 8'hB2; B = 8'h95; #100;
A = 8'hB2; B = 8'h96; #100;
A = 8'hB2; B = 8'h97; #100;
A = 8'hB2; B = 8'h98; #100;
A = 8'hB2; B = 8'h99; #100;
A = 8'hB2; B = 8'h9A; #100;
A = 8'hB2; B = 8'h9B; #100;
A = 8'hB2; B = 8'h9C; #100;
A = 8'hB2; B = 8'h9D; #100;
A = 8'hB2; B = 8'h9E; #100;
A = 8'hB2; B = 8'h9F; #100;
A = 8'hB2; B = 8'hA0; #100;
A = 8'hB2; B = 8'hA1; #100;
A = 8'hB2; B = 8'hA2; #100;
A = 8'hB2; B = 8'hA3; #100;
A = 8'hB2; B = 8'hA4; #100;
A = 8'hB2; B = 8'hA5; #100;
A = 8'hB2; B = 8'hA6; #100;
A = 8'hB2; B = 8'hA7; #100;
A = 8'hB2; B = 8'hA8; #100;
A = 8'hB2; B = 8'hA9; #100;
A = 8'hB2; B = 8'hAA; #100;
A = 8'hB2; B = 8'hAB; #100;
A = 8'hB2; B = 8'hAC; #100;
A = 8'hB2; B = 8'hAD; #100;
A = 8'hB2; B = 8'hAE; #100;
A = 8'hB2; B = 8'hAF; #100;
A = 8'hB2; B = 8'hB0; #100;
A = 8'hB2; B = 8'hB1; #100;
A = 8'hB2; B = 8'hB2; #100;
A = 8'hB2; B = 8'hB3; #100;
A = 8'hB2; B = 8'hB4; #100;
A = 8'hB2; B = 8'hB5; #100;
A = 8'hB2; B = 8'hB6; #100;
A = 8'hB2; B = 8'hB7; #100;
A = 8'hB2; B = 8'hB8; #100;
A = 8'hB2; B = 8'hB9; #100;
A = 8'hB2; B = 8'hBA; #100;
A = 8'hB2; B = 8'hBB; #100;
A = 8'hB2; B = 8'hBC; #100;
A = 8'hB2; B = 8'hBD; #100;
A = 8'hB2; B = 8'hBE; #100;
A = 8'hB2; B = 8'hBF; #100;
A = 8'hB2; B = 8'hC0; #100;
A = 8'hB2; B = 8'hC1; #100;
A = 8'hB2; B = 8'hC2; #100;
A = 8'hB2; B = 8'hC3; #100;
A = 8'hB2; B = 8'hC4; #100;
A = 8'hB2; B = 8'hC5; #100;
A = 8'hB2; B = 8'hC6; #100;
A = 8'hB2; B = 8'hC7; #100;
A = 8'hB2; B = 8'hC8; #100;
A = 8'hB2; B = 8'hC9; #100;
A = 8'hB2; B = 8'hCA; #100;
A = 8'hB2; B = 8'hCB; #100;
A = 8'hB2; B = 8'hCC; #100;
A = 8'hB2; B = 8'hCD; #100;
A = 8'hB2; B = 8'hCE; #100;
A = 8'hB2; B = 8'hCF; #100;
A = 8'hB2; B = 8'hD0; #100;
A = 8'hB2; B = 8'hD1; #100;
A = 8'hB2; B = 8'hD2; #100;
A = 8'hB2; B = 8'hD3; #100;
A = 8'hB2; B = 8'hD4; #100;
A = 8'hB2; B = 8'hD5; #100;
A = 8'hB2; B = 8'hD6; #100;
A = 8'hB2; B = 8'hD7; #100;
A = 8'hB2; B = 8'hD8; #100;
A = 8'hB2; B = 8'hD9; #100;
A = 8'hB2; B = 8'hDA; #100;
A = 8'hB2; B = 8'hDB; #100;
A = 8'hB2; B = 8'hDC; #100;
A = 8'hB2; B = 8'hDD; #100;
A = 8'hB2; B = 8'hDE; #100;
A = 8'hB2; B = 8'hDF; #100;
A = 8'hB2; B = 8'hE0; #100;
A = 8'hB2; B = 8'hE1; #100;
A = 8'hB2; B = 8'hE2; #100;
A = 8'hB2; B = 8'hE3; #100;
A = 8'hB2; B = 8'hE4; #100;
A = 8'hB2; B = 8'hE5; #100;
A = 8'hB2; B = 8'hE6; #100;
A = 8'hB2; B = 8'hE7; #100;
A = 8'hB2; B = 8'hE8; #100;
A = 8'hB2; B = 8'hE9; #100;
A = 8'hB2; B = 8'hEA; #100;
A = 8'hB2; B = 8'hEB; #100;
A = 8'hB2; B = 8'hEC; #100;
A = 8'hB2; B = 8'hED; #100;
A = 8'hB2; B = 8'hEE; #100;
A = 8'hB2; B = 8'hEF; #100;
A = 8'hB2; B = 8'hF0; #100;
A = 8'hB2; B = 8'hF1; #100;
A = 8'hB2; B = 8'hF2; #100;
A = 8'hB2; B = 8'hF3; #100;
A = 8'hB2; B = 8'hF4; #100;
A = 8'hB2; B = 8'hF5; #100;
A = 8'hB2; B = 8'hF6; #100;
A = 8'hB2; B = 8'hF7; #100;
A = 8'hB2; B = 8'hF8; #100;
A = 8'hB2; B = 8'hF9; #100;
A = 8'hB2; B = 8'hFA; #100;
A = 8'hB2; B = 8'hFB; #100;
A = 8'hB2; B = 8'hFC; #100;
A = 8'hB2; B = 8'hFD; #100;
A = 8'hB2; B = 8'hFE; #100;
A = 8'hB2; B = 8'hFF; #100;
A = 8'hB3; B = 8'h0; #100;
A = 8'hB3; B = 8'h1; #100;
A = 8'hB3; B = 8'h2; #100;
A = 8'hB3; B = 8'h3; #100;
A = 8'hB3; B = 8'h4; #100;
A = 8'hB3; B = 8'h5; #100;
A = 8'hB3; B = 8'h6; #100;
A = 8'hB3; B = 8'h7; #100;
A = 8'hB3; B = 8'h8; #100;
A = 8'hB3; B = 8'h9; #100;
A = 8'hB3; B = 8'hA; #100;
A = 8'hB3; B = 8'hB; #100;
A = 8'hB3; B = 8'hC; #100;
A = 8'hB3; B = 8'hD; #100;
A = 8'hB3; B = 8'hE; #100;
A = 8'hB3; B = 8'hF; #100;
A = 8'hB3; B = 8'h10; #100;
A = 8'hB3; B = 8'h11; #100;
A = 8'hB3; B = 8'h12; #100;
A = 8'hB3; B = 8'h13; #100;
A = 8'hB3; B = 8'h14; #100;
A = 8'hB3; B = 8'h15; #100;
A = 8'hB3; B = 8'h16; #100;
A = 8'hB3; B = 8'h17; #100;
A = 8'hB3; B = 8'h18; #100;
A = 8'hB3; B = 8'h19; #100;
A = 8'hB3; B = 8'h1A; #100;
A = 8'hB3; B = 8'h1B; #100;
A = 8'hB3; B = 8'h1C; #100;
A = 8'hB3; B = 8'h1D; #100;
A = 8'hB3; B = 8'h1E; #100;
A = 8'hB3; B = 8'h1F; #100;
A = 8'hB3; B = 8'h20; #100;
A = 8'hB3; B = 8'h21; #100;
A = 8'hB3; B = 8'h22; #100;
A = 8'hB3; B = 8'h23; #100;
A = 8'hB3; B = 8'h24; #100;
A = 8'hB3; B = 8'h25; #100;
A = 8'hB3; B = 8'h26; #100;
A = 8'hB3; B = 8'h27; #100;
A = 8'hB3; B = 8'h28; #100;
A = 8'hB3; B = 8'h29; #100;
A = 8'hB3; B = 8'h2A; #100;
A = 8'hB3; B = 8'h2B; #100;
A = 8'hB3; B = 8'h2C; #100;
A = 8'hB3; B = 8'h2D; #100;
A = 8'hB3; B = 8'h2E; #100;
A = 8'hB3; B = 8'h2F; #100;
A = 8'hB3; B = 8'h30; #100;
A = 8'hB3; B = 8'h31; #100;
A = 8'hB3; B = 8'h32; #100;
A = 8'hB3; B = 8'h33; #100;
A = 8'hB3; B = 8'h34; #100;
A = 8'hB3; B = 8'h35; #100;
A = 8'hB3; B = 8'h36; #100;
A = 8'hB3; B = 8'h37; #100;
A = 8'hB3; B = 8'h38; #100;
A = 8'hB3; B = 8'h39; #100;
A = 8'hB3; B = 8'h3A; #100;
A = 8'hB3; B = 8'h3B; #100;
A = 8'hB3; B = 8'h3C; #100;
A = 8'hB3; B = 8'h3D; #100;
A = 8'hB3; B = 8'h3E; #100;
A = 8'hB3; B = 8'h3F; #100;
A = 8'hB3; B = 8'h40; #100;
A = 8'hB3; B = 8'h41; #100;
A = 8'hB3; B = 8'h42; #100;
A = 8'hB3; B = 8'h43; #100;
A = 8'hB3; B = 8'h44; #100;
A = 8'hB3; B = 8'h45; #100;
A = 8'hB3; B = 8'h46; #100;
A = 8'hB3; B = 8'h47; #100;
A = 8'hB3; B = 8'h48; #100;
A = 8'hB3; B = 8'h49; #100;
A = 8'hB3; B = 8'h4A; #100;
A = 8'hB3; B = 8'h4B; #100;
A = 8'hB3; B = 8'h4C; #100;
A = 8'hB3; B = 8'h4D; #100;
A = 8'hB3; B = 8'h4E; #100;
A = 8'hB3; B = 8'h4F; #100;
A = 8'hB3; B = 8'h50; #100;
A = 8'hB3; B = 8'h51; #100;
A = 8'hB3; B = 8'h52; #100;
A = 8'hB3; B = 8'h53; #100;
A = 8'hB3; B = 8'h54; #100;
A = 8'hB3; B = 8'h55; #100;
A = 8'hB3; B = 8'h56; #100;
A = 8'hB3; B = 8'h57; #100;
A = 8'hB3; B = 8'h58; #100;
A = 8'hB3; B = 8'h59; #100;
A = 8'hB3; B = 8'h5A; #100;
A = 8'hB3; B = 8'h5B; #100;
A = 8'hB3; B = 8'h5C; #100;
A = 8'hB3; B = 8'h5D; #100;
A = 8'hB3; B = 8'h5E; #100;
A = 8'hB3; B = 8'h5F; #100;
A = 8'hB3; B = 8'h60; #100;
A = 8'hB3; B = 8'h61; #100;
A = 8'hB3; B = 8'h62; #100;
A = 8'hB3; B = 8'h63; #100;
A = 8'hB3; B = 8'h64; #100;
A = 8'hB3; B = 8'h65; #100;
A = 8'hB3; B = 8'h66; #100;
A = 8'hB3; B = 8'h67; #100;
A = 8'hB3; B = 8'h68; #100;
A = 8'hB3; B = 8'h69; #100;
A = 8'hB3; B = 8'h6A; #100;
A = 8'hB3; B = 8'h6B; #100;
A = 8'hB3; B = 8'h6C; #100;
A = 8'hB3; B = 8'h6D; #100;
A = 8'hB3; B = 8'h6E; #100;
A = 8'hB3; B = 8'h6F; #100;
A = 8'hB3; B = 8'h70; #100;
A = 8'hB3; B = 8'h71; #100;
A = 8'hB3; B = 8'h72; #100;
A = 8'hB3; B = 8'h73; #100;
A = 8'hB3; B = 8'h74; #100;
A = 8'hB3; B = 8'h75; #100;
A = 8'hB3; B = 8'h76; #100;
A = 8'hB3; B = 8'h77; #100;
A = 8'hB3; B = 8'h78; #100;
A = 8'hB3; B = 8'h79; #100;
A = 8'hB3; B = 8'h7A; #100;
A = 8'hB3; B = 8'h7B; #100;
A = 8'hB3; B = 8'h7C; #100;
A = 8'hB3; B = 8'h7D; #100;
A = 8'hB3; B = 8'h7E; #100;
A = 8'hB3; B = 8'h7F; #100;
A = 8'hB3; B = 8'h80; #100;
A = 8'hB3; B = 8'h81; #100;
A = 8'hB3; B = 8'h82; #100;
A = 8'hB3; B = 8'h83; #100;
A = 8'hB3; B = 8'h84; #100;
A = 8'hB3; B = 8'h85; #100;
A = 8'hB3; B = 8'h86; #100;
A = 8'hB3; B = 8'h87; #100;
A = 8'hB3; B = 8'h88; #100;
A = 8'hB3; B = 8'h89; #100;
A = 8'hB3; B = 8'h8A; #100;
A = 8'hB3; B = 8'h8B; #100;
A = 8'hB3; B = 8'h8C; #100;
A = 8'hB3; B = 8'h8D; #100;
A = 8'hB3; B = 8'h8E; #100;
A = 8'hB3; B = 8'h8F; #100;
A = 8'hB3; B = 8'h90; #100;
A = 8'hB3; B = 8'h91; #100;
A = 8'hB3; B = 8'h92; #100;
A = 8'hB3; B = 8'h93; #100;
A = 8'hB3; B = 8'h94; #100;
A = 8'hB3; B = 8'h95; #100;
A = 8'hB3; B = 8'h96; #100;
A = 8'hB3; B = 8'h97; #100;
A = 8'hB3; B = 8'h98; #100;
A = 8'hB3; B = 8'h99; #100;
A = 8'hB3; B = 8'h9A; #100;
A = 8'hB3; B = 8'h9B; #100;
A = 8'hB3; B = 8'h9C; #100;
A = 8'hB3; B = 8'h9D; #100;
A = 8'hB3; B = 8'h9E; #100;
A = 8'hB3; B = 8'h9F; #100;
A = 8'hB3; B = 8'hA0; #100;
A = 8'hB3; B = 8'hA1; #100;
A = 8'hB3; B = 8'hA2; #100;
A = 8'hB3; B = 8'hA3; #100;
A = 8'hB3; B = 8'hA4; #100;
A = 8'hB3; B = 8'hA5; #100;
A = 8'hB3; B = 8'hA6; #100;
A = 8'hB3; B = 8'hA7; #100;
A = 8'hB3; B = 8'hA8; #100;
A = 8'hB3; B = 8'hA9; #100;
A = 8'hB3; B = 8'hAA; #100;
A = 8'hB3; B = 8'hAB; #100;
A = 8'hB3; B = 8'hAC; #100;
A = 8'hB3; B = 8'hAD; #100;
A = 8'hB3; B = 8'hAE; #100;
A = 8'hB3; B = 8'hAF; #100;
A = 8'hB3; B = 8'hB0; #100;
A = 8'hB3; B = 8'hB1; #100;
A = 8'hB3; B = 8'hB2; #100;
A = 8'hB3; B = 8'hB3; #100;
A = 8'hB3; B = 8'hB4; #100;
A = 8'hB3; B = 8'hB5; #100;
A = 8'hB3; B = 8'hB6; #100;
A = 8'hB3; B = 8'hB7; #100;
A = 8'hB3; B = 8'hB8; #100;
A = 8'hB3; B = 8'hB9; #100;
A = 8'hB3; B = 8'hBA; #100;
A = 8'hB3; B = 8'hBB; #100;
A = 8'hB3; B = 8'hBC; #100;
A = 8'hB3; B = 8'hBD; #100;
A = 8'hB3; B = 8'hBE; #100;
A = 8'hB3; B = 8'hBF; #100;
A = 8'hB3; B = 8'hC0; #100;
A = 8'hB3; B = 8'hC1; #100;
A = 8'hB3; B = 8'hC2; #100;
A = 8'hB3; B = 8'hC3; #100;
A = 8'hB3; B = 8'hC4; #100;
A = 8'hB3; B = 8'hC5; #100;
A = 8'hB3; B = 8'hC6; #100;
A = 8'hB3; B = 8'hC7; #100;
A = 8'hB3; B = 8'hC8; #100;
A = 8'hB3; B = 8'hC9; #100;
A = 8'hB3; B = 8'hCA; #100;
A = 8'hB3; B = 8'hCB; #100;
A = 8'hB3; B = 8'hCC; #100;
A = 8'hB3; B = 8'hCD; #100;
A = 8'hB3; B = 8'hCE; #100;
A = 8'hB3; B = 8'hCF; #100;
A = 8'hB3; B = 8'hD0; #100;
A = 8'hB3; B = 8'hD1; #100;
A = 8'hB3; B = 8'hD2; #100;
A = 8'hB3; B = 8'hD3; #100;
A = 8'hB3; B = 8'hD4; #100;
A = 8'hB3; B = 8'hD5; #100;
A = 8'hB3; B = 8'hD6; #100;
A = 8'hB3; B = 8'hD7; #100;
A = 8'hB3; B = 8'hD8; #100;
A = 8'hB3; B = 8'hD9; #100;
A = 8'hB3; B = 8'hDA; #100;
A = 8'hB3; B = 8'hDB; #100;
A = 8'hB3; B = 8'hDC; #100;
A = 8'hB3; B = 8'hDD; #100;
A = 8'hB3; B = 8'hDE; #100;
A = 8'hB3; B = 8'hDF; #100;
A = 8'hB3; B = 8'hE0; #100;
A = 8'hB3; B = 8'hE1; #100;
A = 8'hB3; B = 8'hE2; #100;
A = 8'hB3; B = 8'hE3; #100;
A = 8'hB3; B = 8'hE4; #100;
A = 8'hB3; B = 8'hE5; #100;
A = 8'hB3; B = 8'hE6; #100;
A = 8'hB3; B = 8'hE7; #100;
A = 8'hB3; B = 8'hE8; #100;
A = 8'hB3; B = 8'hE9; #100;
A = 8'hB3; B = 8'hEA; #100;
A = 8'hB3; B = 8'hEB; #100;
A = 8'hB3; B = 8'hEC; #100;
A = 8'hB3; B = 8'hED; #100;
A = 8'hB3; B = 8'hEE; #100;
A = 8'hB3; B = 8'hEF; #100;
A = 8'hB3; B = 8'hF0; #100;
A = 8'hB3; B = 8'hF1; #100;
A = 8'hB3; B = 8'hF2; #100;
A = 8'hB3; B = 8'hF3; #100;
A = 8'hB3; B = 8'hF4; #100;
A = 8'hB3; B = 8'hF5; #100;
A = 8'hB3; B = 8'hF6; #100;
A = 8'hB3; B = 8'hF7; #100;
A = 8'hB3; B = 8'hF8; #100;
A = 8'hB3; B = 8'hF9; #100;
A = 8'hB3; B = 8'hFA; #100;
A = 8'hB3; B = 8'hFB; #100;
A = 8'hB3; B = 8'hFC; #100;
A = 8'hB3; B = 8'hFD; #100;
A = 8'hB3; B = 8'hFE; #100;
A = 8'hB3; B = 8'hFF; #100;
A = 8'hB4; B = 8'h0; #100;
A = 8'hB4; B = 8'h1; #100;
A = 8'hB4; B = 8'h2; #100;
A = 8'hB4; B = 8'h3; #100;
A = 8'hB4; B = 8'h4; #100;
A = 8'hB4; B = 8'h5; #100;
A = 8'hB4; B = 8'h6; #100;
A = 8'hB4; B = 8'h7; #100;
A = 8'hB4; B = 8'h8; #100;
A = 8'hB4; B = 8'h9; #100;
A = 8'hB4; B = 8'hA; #100;
A = 8'hB4; B = 8'hB; #100;
A = 8'hB4; B = 8'hC; #100;
A = 8'hB4; B = 8'hD; #100;
A = 8'hB4; B = 8'hE; #100;
A = 8'hB4; B = 8'hF; #100;
A = 8'hB4; B = 8'h10; #100;
A = 8'hB4; B = 8'h11; #100;
A = 8'hB4; B = 8'h12; #100;
A = 8'hB4; B = 8'h13; #100;
A = 8'hB4; B = 8'h14; #100;
A = 8'hB4; B = 8'h15; #100;
A = 8'hB4; B = 8'h16; #100;
A = 8'hB4; B = 8'h17; #100;
A = 8'hB4; B = 8'h18; #100;
A = 8'hB4; B = 8'h19; #100;
A = 8'hB4; B = 8'h1A; #100;
A = 8'hB4; B = 8'h1B; #100;
A = 8'hB4; B = 8'h1C; #100;
A = 8'hB4; B = 8'h1D; #100;
A = 8'hB4; B = 8'h1E; #100;
A = 8'hB4; B = 8'h1F; #100;
A = 8'hB4; B = 8'h20; #100;
A = 8'hB4; B = 8'h21; #100;
A = 8'hB4; B = 8'h22; #100;
A = 8'hB4; B = 8'h23; #100;
A = 8'hB4; B = 8'h24; #100;
A = 8'hB4; B = 8'h25; #100;
A = 8'hB4; B = 8'h26; #100;
A = 8'hB4; B = 8'h27; #100;
A = 8'hB4; B = 8'h28; #100;
A = 8'hB4; B = 8'h29; #100;
A = 8'hB4; B = 8'h2A; #100;
A = 8'hB4; B = 8'h2B; #100;
A = 8'hB4; B = 8'h2C; #100;
A = 8'hB4; B = 8'h2D; #100;
A = 8'hB4; B = 8'h2E; #100;
A = 8'hB4; B = 8'h2F; #100;
A = 8'hB4; B = 8'h30; #100;
A = 8'hB4; B = 8'h31; #100;
A = 8'hB4; B = 8'h32; #100;
A = 8'hB4; B = 8'h33; #100;
A = 8'hB4; B = 8'h34; #100;
A = 8'hB4; B = 8'h35; #100;
A = 8'hB4; B = 8'h36; #100;
A = 8'hB4; B = 8'h37; #100;
A = 8'hB4; B = 8'h38; #100;
A = 8'hB4; B = 8'h39; #100;
A = 8'hB4; B = 8'h3A; #100;
A = 8'hB4; B = 8'h3B; #100;
A = 8'hB4; B = 8'h3C; #100;
A = 8'hB4; B = 8'h3D; #100;
A = 8'hB4; B = 8'h3E; #100;
A = 8'hB4; B = 8'h3F; #100;
A = 8'hB4; B = 8'h40; #100;
A = 8'hB4; B = 8'h41; #100;
A = 8'hB4; B = 8'h42; #100;
A = 8'hB4; B = 8'h43; #100;
A = 8'hB4; B = 8'h44; #100;
A = 8'hB4; B = 8'h45; #100;
A = 8'hB4; B = 8'h46; #100;
A = 8'hB4; B = 8'h47; #100;
A = 8'hB4; B = 8'h48; #100;
A = 8'hB4; B = 8'h49; #100;
A = 8'hB4; B = 8'h4A; #100;
A = 8'hB4; B = 8'h4B; #100;
A = 8'hB4; B = 8'h4C; #100;
A = 8'hB4; B = 8'h4D; #100;
A = 8'hB4; B = 8'h4E; #100;
A = 8'hB4; B = 8'h4F; #100;
A = 8'hB4; B = 8'h50; #100;
A = 8'hB4; B = 8'h51; #100;
A = 8'hB4; B = 8'h52; #100;
A = 8'hB4; B = 8'h53; #100;
A = 8'hB4; B = 8'h54; #100;
A = 8'hB4; B = 8'h55; #100;
A = 8'hB4; B = 8'h56; #100;
A = 8'hB4; B = 8'h57; #100;
A = 8'hB4; B = 8'h58; #100;
A = 8'hB4; B = 8'h59; #100;
A = 8'hB4; B = 8'h5A; #100;
A = 8'hB4; B = 8'h5B; #100;
A = 8'hB4; B = 8'h5C; #100;
A = 8'hB4; B = 8'h5D; #100;
A = 8'hB4; B = 8'h5E; #100;
A = 8'hB4; B = 8'h5F; #100;
A = 8'hB4; B = 8'h60; #100;
A = 8'hB4; B = 8'h61; #100;
A = 8'hB4; B = 8'h62; #100;
A = 8'hB4; B = 8'h63; #100;
A = 8'hB4; B = 8'h64; #100;
A = 8'hB4; B = 8'h65; #100;
A = 8'hB4; B = 8'h66; #100;
A = 8'hB4; B = 8'h67; #100;
A = 8'hB4; B = 8'h68; #100;
A = 8'hB4; B = 8'h69; #100;
A = 8'hB4; B = 8'h6A; #100;
A = 8'hB4; B = 8'h6B; #100;
A = 8'hB4; B = 8'h6C; #100;
A = 8'hB4; B = 8'h6D; #100;
A = 8'hB4; B = 8'h6E; #100;
A = 8'hB4; B = 8'h6F; #100;
A = 8'hB4; B = 8'h70; #100;
A = 8'hB4; B = 8'h71; #100;
A = 8'hB4; B = 8'h72; #100;
A = 8'hB4; B = 8'h73; #100;
A = 8'hB4; B = 8'h74; #100;
A = 8'hB4; B = 8'h75; #100;
A = 8'hB4; B = 8'h76; #100;
A = 8'hB4; B = 8'h77; #100;
A = 8'hB4; B = 8'h78; #100;
A = 8'hB4; B = 8'h79; #100;
A = 8'hB4; B = 8'h7A; #100;
A = 8'hB4; B = 8'h7B; #100;
A = 8'hB4; B = 8'h7C; #100;
A = 8'hB4; B = 8'h7D; #100;
A = 8'hB4; B = 8'h7E; #100;
A = 8'hB4; B = 8'h7F; #100;
A = 8'hB4; B = 8'h80; #100;
A = 8'hB4; B = 8'h81; #100;
A = 8'hB4; B = 8'h82; #100;
A = 8'hB4; B = 8'h83; #100;
A = 8'hB4; B = 8'h84; #100;
A = 8'hB4; B = 8'h85; #100;
A = 8'hB4; B = 8'h86; #100;
A = 8'hB4; B = 8'h87; #100;
A = 8'hB4; B = 8'h88; #100;
A = 8'hB4; B = 8'h89; #100;
A = 8'hB4; B = 8'h8A; #100;
A = 8'hB4; B = 8'h8B; #100;
A = 8'hB4; B = 8'h8C; #100;
A = 8'hB4; B = 8'h8D; #100;
A = 8'hB4; B = 8'h8E; #100;
A = 8'hB4; B = 8'h8F; #100;
A = 8'hB4; B = 8'h90; #100;
A = 8'hB4; B = 8'h91; #100;
A = 8'hB4; B = 8'h92; #100;
A = 8'hB4; B = 8'h93; #100;
A = 8'hB4; B = 8'h94; #100;
A = 8'hB4; B = 8'h95; #100;
A = 8'hB4; B = 8'h96; #100;
A = 8'hB4; B = 8'h97; #100;
A = 8'hB4; B = 8'h98; #100;
A = 8'hB4; B = 8'h99; #100;
A = 8'hB4; B = 8'h9A; #100;
A = 8'hB4; B = 8'h9B; #100;
A = 8'hB4; B = 8'h9C; #100;
A = 8'hB4; B = 8'h9D; #100;
A = 8'hB4; B = 8'h9E; #100;
A = 8'hB4; B = 8'h9F; #100;
A = 8'hB4; B = 8'hA0; #100;
A = 8'hB4; B = 8'hA1; #100;
A = 8'hB4; B = 8'hA2; #100;
A = 8'hB4; B = 8'hA3; #100;
A = 8'hB4; B = 8'hA4; #100;
A = 8'hB4; B = 8'hA5; #100;
A = 8'hB4; B = 8'hA6; #100;
A = 8'hB4; B = 8'hA7; #100;
A = 8'hB4; B = 8'hA8; #100;
A = 8'hB4; B = 8'hA9; #100;
A = 8'hB4; B = 8'hAA; #100;
A = 8'hB4; B = 8'hAB; #100;
A = 8'hB4; B = 8'hAC; #100;
A = 8'hB4; B = 8'hAD; #100;
A = 8'hB4; B = 8'hAE; #100;
A = 8'hB4; B = 8'hAF; #100;
A = 8'hB4; B = 8'hB0; #100;
A = 8'hB4; B = 8'hB1; #100;
A = 8'hB4; B = 8'hB2; #100;
A = 8'hB4; B = 8'hB3; #100;
A = 8'hB4; B = 8'hB4; #100;
A = 8'hB4; B = 8'hB5; #100;
A = 8'hB4; B = 8'hB6; #100;
A = 8'hB4; B = 8'hB7; #100;
A = 8'hB4; B = 8'hB8; #100;
A = 8'hB4; B = 8'hB9; #100;
A = 8'hB4; B = 8'hBA; #100;
A = 8'hB4; B = 8'hBB; #100;
A = 8'hB4; B = 8'hBC; #100;
A = 8'hB4; B = 8'hBD; #100;
A = 8'hB4; B = 8'hBE; #100;
A = 8'hB4; B = 8'hBF; #100;
A = 8'hB4; B = 8'hC0; #100;
A = 8'hB4; B = 8'hC1; #100;
A = 8'hB4; B = 8'hC2; #100;
A = 8'hB4; B = 8'hC3; #100;
A = 8'hB4; B = 8'hC4; #100;
A = 8'hB4; B = 8'hC5; #100;
A = 8'hB4; B = 8'hC6; #100;
A = 8'hB4; B = 8'hC7; #100;
A = 8'hB4; B = 8'hC8; #100;
A = 8'hB4; B = 8'hC9; #100;
A = 8'hB4; B = 8'hCA; #100;
A = 8'hB4; B = 8'hCB; #100;
A = 8'hB4; B = 8'hCC; #100;
A = 8'hB4; B = 8'hCD; #100;
A = 8'hB4; B = 8'hCE; #100;
A = 8'hB4; B = 8'hCF; #100;
A = 8'hB4; B = 8'hD0; #100;
A = 8'hB4; B = 8'hD1; #100;
A = 8'hB4; B = 8'hD2; #100;
A = 8'hB4; B = 8'hD3; #100;
A = 8'hB4; B = 8'hD4; #100;
A = 8'hB4; B = 8'hD5; #100;
A = 8'hB4; B = 8'hD6; #100;
A = 8'hB4; B = 8'hD7; #100;
A = 8'hB4; B = 8'hD8; #100;
A = 8'hB4; B = 8'hD9; #100;
A = 8'hB4; B = 8'hDA; #100;
A = 8'hB4; B = 8'hDB; #100;
A = 8'hB4; B = 8'hDC; #100;
A = 8'hB4; B = 8'hDD; #100;
A = 8'hB4; B = 8'hDE; #100;
A = 8'hB4; B = 8'hDF; #100;
A = 8'hB4; B = 8'hE0; #100;
A = 8'hB4; B = 8'hE1; #100;
A = 8'hB4; B = 8'hE2; #100;
A = 8'hB4; B = 8'hE3; #100;
A = 8'hB4; B = 8'hE4; #100;
A = 8'hB4; B = 8'hE5; #100;
A = 8'hB4; B = 8'hE6; #100;
A = 8'hB4; B = 8'hE7; #100;
A = 8'hB4; B = 8'hE8; #100;
A = 8'hB4; B = 8'hE9; #100;
A = 8'hB4; B = 8'hEA; #100;
A = 8'hB4; B = 8'hEB; #100;
A = 8'hB4; B = 8'hEC; #100;
A = 8'hB4; B = 8'hED; #100;
A = 8'hB4; B = 8'hEE; #100;
A = 8'hB4; B = 8'hEF; #100;
A = 8'hB4; B = 8'hF0; #100;
A = 8'hB4; B = 8'hF1; #100;
A = 8'hB4; B = 8'hF2; #100;
A = 8'hB4; B = 8'hF3; #100;
A = 8'hB4; B = 8'hF4; #100;
A = 8'hB4; B = 8'hF5; #100;
A = 8'hB4; B = 8'hF6; #100;
A = 8'hB4; B = 8'hF7; #100;
A = 8'hB4; B = 8'hF8; #100;
A = 8'hB4; B = 8'hF9; #100;
A = 8'hB4; B = 8'hFA; #100;
A = 8'hB4; B = 8'hFB; #100;
A = 8'hB4; B = 8'hFC; #100;
A = 8'hB4; B = 8'hFD; #100;
A = 8'hB4; B = 8'hFE; #100;
A = 8'hB4; B = 8'hFF; #100;
A = 8'hB5; B = 8'h0; #100;
A = 8'hB5; B = 8'h1; #100;
A = 8'hB5; B = 8'h2; #100;
A = 8'hB5; B = 8'h3; #100;
A = 8'hB5; B = 8'h4; #100;
A = 8'hB5; B = 8'h5; #100;
A = 8'hB5; B = 8'h6; #100;
A = 8'hB5; B = 8'h7; #100;
A = 8'hB5; B = 8'h8; #100;
A = 8'hB5; B = 8'h9; #100;
A = 8'hB5; B = 8'hA; #100;
A = 8'hB5; B = 8'hB; #100;
A = 8'hB5; B = 8'hC; #100;
A = 8'hB5; B = 8'hD; #100;
A = 8'hB5; B = 8'hE; #100;
A = 8'hB5; B = 8'hF; #100;
A = 8'hB5; B = 8'h10; #100;
A = 8'hB5; B = 8'h11; #100;
A = 8'hB5; B = 8'h12; #100;
A = 8'hB5; B = 8'h13; #100;
A = 8'hB5; B = 8'h14; #100;
A = 8'hB5; B = 8'h15; #100;
A = 8'hB5; B = 8'h16; #100;
A = 8'hB5; B = 8'h17; #100;
A = 8'hB5; B = 8'h18; #100;
A = 8'hB5; B = 8'h19; #100;
A = 8'hB5; B = 8'h1A; #100;
A = 8'hB5; B = 8'h1B; #100;
A = 8'hB5; B = 8'h1C; #100;
A = 8'hB5; B = 8'h1D; #100;
A = 8'hB5; B = 8'h1E; #100;
A = 8'hB5; B = 8'h1F; #100;
A = 8'hB5; B = 8'h20; #100;
A = 8'hB5; B = 8'h21; #100;
A = 8'hB5; B = 8'h22; #100;
A = 8'hB5; B = 8'h23; #100;
A = 8'hB5; B = 8'h24; #100;
A = 8'hB5; B = 8'h25; #100;
A = 8'hB5; B = 8'h26; #100;
A = 8'hB5; B = 8'h27; #100;
A = 8'hB5; B = 8'h28; #100;
A = 8'hB5; B = 8'h29; #100;
A = 8'hB5; B = 8'h2A; #100;
A = 8'hB5; B = 8'h2B; #100;
A = 8'hB5; B = 8'h2C; #100;
A = 8'hB5; B = 8'h2D; #100;
A = 8'hB5; B = 8'h2E; #100;
A = 8'hB5; B = 8'h2F; #100;
A = 8'hB5; B = 8'h30; #100;
A = 8'hB5; B = 8'h31; #100;
A = 8'hB5; B = 8'h32; #100;
A = 8'hB5; B = 8'h33; #100;
A = 8'hB5; B = 8'h34; #100;
A = 8'hB5; B = 8'h35; #100;
A = 8'hB5; B = 8'h36; #100;
A = 8'hB5; B = 8'h37; #100;
A = 8'hB5; B = 8'h38; #100;
A = 8'hB5; B = 8'h39; #100;
A = 8'hB5; B = 8'h3A; #100;
A = 8'hB5; B = 8'h3B; #100;
A = 8'hB5; B = 8'h3C; #100;
A = 8'hB5; B = 8'h3D; #100;
A = 8'hB5; B = 8'h3E; #100;
A = 8'hB5; B = 8'h3F; #100;
A = 8'hB5; B = 8'h40; #100;
A = 8'hB5; B = 8'h41; #100;
A = 8'hB5; B = 8'h42; #100;
A = 8'hB5; B = 8'h43; #100;
A = 8'hB5; B = 8'h44; #100;
A = 8'hB5; B = 8'h45; #100;
A = 8'hB5; B = 8'h46; #100;
A = 8'hB5; B = 8'h47; #100;
A = 8'hB5; B = 8'h48; #100;
A = 8'hB5; B = 8'h49; #100;
A = 8'hB5; B = 8'h4A; #100;
A = 8'hB5; B = 8'h4B; #100;
A = 8'hB5; B = 8'h4C; #100;
A = 8'hB5; B = 8'h4D; #100;
A = 8'hB5; B = 8'h4E; #100;
A = 8'hB5; B = 8'h4F; #100;
A = 8'hB5; B = 8'h50; #100;
A = 8'hB5; B = 8'h51; #100;
A = 8'hB5; B = 8'h52; #100;
A = 8'hB5; B = 8'h53; #100;
A = 8'hB5; B = 8'h54; #100;
A = 8'hB5; B = 8'h55; #100;
A = 8'hB5; B = 8'h56; #100;
A = 8'hB5; B = 8'h57; #100;
A = 8'hB5; B = 8'h58; #100;
A = 8'hB5; B = 8'h59; #100;
A = 8'hB5; B = 8'h5A; #100;
A = 8'hB5; B = 8'h5B; #100;
A = 8'hB5; B = 8'h5C; #100;
A = 8'hB5; B = 8'h5D; #100;
A = 8'hB5; B = 8'h5E; #100;
A = 8'hB5; B = 8'h5F; #100;
A = 8'hB5; B = 8'h60; #100;
A = 8'hB5; B = 8'h61; #100;
A = 8'hB5; B = 8'h62; #100;
A = 8'hB5; B = 8'h63; #100;
A = 8'hB5; B = 8'h64; #100;
A = 8'hB5; B = 8'h65; #100;
A = 8'hB5; B = 8'h66; #100;
A = 8'hB5; B = 8'h67; #100;
A = 8'hB5; B = 8'h68; #100;
A = 8'hB5; B = 8'h69; #100;
A = 8'hB5; B = 8'h6A; #100;
A = 8'hB5; B = 8'h6B; #100;
A = 8'hB5; B = 8'h6C; #100;
A = 8'hB5; B = 8'h6D; #100;
A = 8'hB5; B = 8'h6E; #100;
A = 8'hB5; B = 8'h6F; #100;
A = 8'hB5; B = 8'h70; #100;
A = 8'hB5; B = 8'h71; #100;
A = 8'hB5; B = 8'h72; #100;
A = 8'hB5; B = 8'h73; #100;
A = 8'hB5; B = 8'h74; #100;
A = 8'hB5; B = 8'h75; #100;
A = 8'hB5; B = 8'h76; #100;
A = 8'hB5; B = 8'h77; #100;
A = 8'hB5; B = 8'h78; #100;
A = 8'hB5; B = 8'h79; #100;
A = 8'hB5; B = 8'h7A; #100;
A = 8'hB5; B = 8'h7B; #100;
A = 8'hB5; B = 8'h7C; #100;
A = 8'hB5; B = 8'h7D; #100;
A = 8'hB5; B = 8'h7E; #100;
A = 8'hB5; B = 8'h7F; #100;
A = 8'hB5; B = 8'h80; #100;
A = 8'hB5; B = 8'h81; #100;
A = 8'hB5; B = 8'h82; #100;
A = 8'hB5; B = 8'h83; #100;
A = 8'hB5; B = 8'h84; #100;
A = 8'hB5; B = 8'h85; #100;
A = 8'hB5; B = 8'h86; #100;
A = 8'hB5; B = 8'h87; #100;
A = 8'hB5; B = 8'h88; #100;
A = 8'hB5; B = 8'h89; #100;
A = 8'hB5; B = 8'h8A; #100;
A = 8'hB5; B = 8'h8B; #100;
A = 8'hB5; B = 8'h8C; #100;
A = 8'hB5; B = 8'h8D; #100;
A = 8'hB5; B = 8'h8E; #100;
A = 8'hB5; B = 8'h8F; #100;
A = 8'hB5; B = 8'h90; #100;
A = 8'hB5; B = 8'h91; #100;
A = 8'hB5; B = 8'h92; #100;
A = 8'hB5; B = 8'h93; #100;
A = 8'hB5; B = 8'h94; #100;
A = 8'hB5; B = 8'h95; #100;
A = 8'hB5; B = 8'h96; #100;
A = 8'hB5; B = 8'h97; #100;
A = 8'hB5; B = 8'h98; #100;
A = 8'hB5; B = 8'h99; #100;
A = 8'hB5; B = 8'h9A; #100;
A = 8'hB5; B = 8'h9B; #100;
A = 8'hB5; B = 8'h9C; #100;
A = 8'hB5; B = 8'h9D; #100;
A = 8'hB5; B = 8'h9E; #100;
A = 8'hB5; B = 8'h9F; #100;
A = 8'hB5; B = 8'hA0; #100;
A = 8'hB5; B = 8'hA1; #100;
A = 8'hB5; B = 8'hA2; #100;
A = 8'hB5; B = 8'hA3; #100;
A = 8'hB5; B = 8'hA4; #100;
A = 8'hB5; B = 8'hA5; #100;
A = 8'hB5; B = 8'hA6; #100;
A = 8'hB5; B = 8'hA7; #100;
A = 8'hB5; B = 8'hA8; #100;
A = 8'hB5; B = 8'hA9; #100;
A = 8'hB5; B = 8'hAA; #100;
A = 8'hB5; B = 8'hAB; #100;
A = 8'hB5; B = 8'hAC; #100;
A = 8'hB5; B = 8'hAD; #100;
A = 8'hB5; B = 8'hAE; #100;
A = 8'hB5; B = 8'hAF; #100;
A = 8'hB5; B = 8'hB0; #100;
A = 8'hB5; B = 8'hB1; #100;
A = 8'hB5; B = 8'hB2; #100;
A = 8'hB5; B = 8'hB3; #100;
A = 8'hB5; B = 8'hB4; #100;
A = 8'hB5; B = 8'hB5; #100;
A = 8'hB5; B = 8'hB6; #100;
A = 8'hB5; B = 8'hB7; #100;
A = 8'hB5; B = 8'hB8; #100;
A = 8'hB5; B = 8'hB9; #100;
A = 8'hB5; B = 8'hBA; #100;
A = 8'hB5; B = 8'hBB; #100;
A = 8'hB5; B = 8'hBC; #100;
A = 8'hB5; B = 8'hBD; #100;
A = 8'hB5; B = 8'hBE; #100;
A = 8'hB5; B = 8'hBF; #100;
A = 8'hB5; B = 8'hC0; #100;
A = 8'hB5; B = 8'hC1; #100;
A = 8'hB5; B = 8'hC2; #100;
A = 8'hB5; B = 8'hC3; #100;
A = 8'hB5; B = 8'hC4; #100;
A = 8'hB5; B = 8'hC5; #100;
A = 8'hB5; B = 8'hC6; #100;
A = 8'hB5; B = 8'hC7; #100;
A = 8'hB5; B = 8'hC8; #100;
A = 8'hB5; B = 8'hC9; #100;
A = 8'hB5; B = 8'hCA; #100;
A = 8'hB5; B = 8'hCB; #100;
A = 8'hB5; B = 8'hCC; #100;
A = 8'hB5; B = 8'hCD; #100;
A = 8'hB5; B = 8'hCE; #100;
A = 8'hB5; B = 8'hCF; #100;
A = 8'hB5; B = 8'hD0; #100;
A = 8'hB5; B = 8'hD1; #100;
A = 8'hB5; B = 8'hD2; #100;
A = 8'hB5; B = 8'hD3; #100;
A = 8'hB5; B = 8'hD4; #100;
A = 8'hB5; B = 8'hD5; #100;
A = 8'hB5; B = 8'hD6; #100;
A = 8'hB5; B = 8'hD7; #100;
A = 8'hB5; B = 8'hD8; #100;
A = 8'hB5; B = 8'hD9; #100;
A = 8'hB5; B = 8'hDA; #100;
A = 8'hB5; B = 8'hDB; #100;
A = 8'hB5; B = 8'hDC; #100;
A = 8'hB5; B = 8'hDD; #100;
A = 8'hB5; B = 8'hDE; #100;
A = 8'hB5; B = 8'hDF; #100;
A = 8'hB5; B = 8'hE0; #100;
A = 8'hB5; B = 8'hE1; #100;
A = 8'hB5; B = 8'hE2; #100;
A = 8'hB5; B = 8'hE3; #100;
A = 8'hB5; B = 8'hE4; #100;
A = 8'hB5; B = 8'hE5; #100;
A = 8'hB5; B = 8'hE6; #100;
A = 8'hB5; B = 8'hE7; #100;
A = 8'hB5; B = 8'hE8; #100;
A = 8'hB5; B = 8'hE9; #100;
A = 8'hB5; B = 8'hEA; #100;
A = 8'hB5; B = 8'hEB; #100;
A = 8'hB5; B = 8'hEC; #100;
A = 8'hB5; B = 8'hED; #100;
A = 8'hB5; B = 8'hEE; #100;
A = 8'hB5; B = 8'hEF; #100;
A = 8'hB5; B = 8'hF0; #100;
A = 8'hB5; B = 8'hF1; #100;
A = 8'hB5; B = 8'hF2; #100;
A = 8'hB5; B = 8'hF3; #100;
A = 8'hB5; B = 8'hF4; #100;
A = 8'hB5; B = 8'hF5; #100;
A = 8'hB5; B = 8'hF6; #100;
A = 8'hB5; B = 8'hF7; #100;
A = 8'hB5; B = 8'hF8; #100;
A = 8'hB5; B = 8'hF9; #100;
A = 8'hB5; B = 8'hFA; #100;
A = 8'hB5; B = 8'hFB; #100;
A = 8'hB5; B = 8'hFC; #100;
A = 8'hB5; B = 8'hFD; #100;
A = 8'hB5; B = 8'hFE; #100;
A = 8'hB5; B = 8'hFF; #100;
A = 8'hB6; B = 8'h0; #100;
A = 8'hB6; B = 8'h1; #100;
A = 8'hB6; B = 8'h2; #100;
A = 8'hB6; B = 8'h3; #100;
A = 8'hB6; B = 8'h4; #100;
A = 8'hB6; B = 8'h5; #100;
A = 8'hB6; B = 8'h6; #100;
A = 8'hB6; B = 8'h7; #100;
A = 8'hB6; B = 8'h8; #100;
A = 8'hB6; B = 8'h9; #100;
A = 8'hB6; B = 8'hA; #100;
A = 8'hB6; B = 8'hB; #100;
A = 8'hB6; B = 8'hC; #100;
A = 8'hB6; B = 8'hD; #100;
A = 8'hB6; B = 8'hE; #100;
A = 8'hB6; B = 8'hF; #100;
A = 8'hB6; B = 8'h10; #100;
A = 8'hB6; B = 8'h11; #100;
A = 8'hB6; B = 8'h12; #100;
A = 8'hB6; B = 8'h13; #100;
A = 8'hB6; B = 8'h14; #100;
A = 8'hB6; B = 8'h15; #100;
A = 8'hB6; B = 8'h16; #100;
A = 8'hB6; B = 8'h17; #100;
A = 8'hB6; B = 8'h18; #100;
A = 8'hB6; B = 8'h19; #100;
A = 8'hB6; B = 8'h1A; #100;
A = 8'hB6; B = 8'h1B; #100;
A = 8'hB6; B = 8'h1C; #100;
A = 8'hB6; B = 8'h1D; #100;
A = 8'hB6; B = 8'h1E; #100;
A = 8'hB6; B = 8'h1F; #100;
A = 8'hB6; B = 8'h20; #100;
A = 8'hB6; B = 8'h21; #100;
A = 8'hB6; B = 8'h22; #100;
A = 8'hB6; B = 8'h23; #100;
A = 8'hB6; B = 8'h24; #100;
A = 8'hB6; B = 8'h25; #100;
A = 8'hB6; B = 8'h26; #100;
A = 8'hB6; B = 8'h27; #100;
A = 8'hB6; B = 8'h28; #100;
A = 8'hB6; B = 8'h29; #100;
A = 8'hB6; B = 8'h2A; #100;
A = 8'hB6; B = 8'h2B; #100;
A = 8'hB6; B = 8'h2C; #100;
A = 8'hB6; B = 8'h2D; #100;
A = 8'hB6; B = 8'h2E; #100;
A = 8'hB6; B = 8'h2F; #100;
A = 8'hB6; B = 8'h30; #100;
A = 8'hB6; B = 8'h31; #100;
A = 8'hB6; B = 8'h32; #100;
A = 8'hB6; B = 8'h33; #100;
A = 8'hB6; B = 8'h34; #100;
A = 8'hB6; B = 8'h35; #100;
A = 8'hB6; B = 8'h36; #100;
A = 8'hB6; B = 8'h37; #100;
A = 8'hB6; B = 8'h38; #100;
A = 8'hB6; B = 8'h39; #100;
A = 8'hB6; B = 8'h3A; #100;
A = 8'hB6; B = 8'h3B; #100;
A = 8'hB6; B = 8'h3C; #100;
A = 8'hB6; B = 8'h3D; #100;
A = 8'hB6; B = 8'h3E; #100;
A = 8'hB6; B = 8'h3F; #100;
A = 8'hB6; B = 8'h40; #100;
A = 8'hB6; B = 8'h41; #100;
A = 8'hB6; B = 8'h42; #100;
A = 8'hB6; B = 8'h43; #100;
A = 8'hB6; B = 8'h44; #100;
A = 8'hB6; B = 8'h45; #100;
A = 8'hB6; B = 8'h46; #100;
A = 8'hB6; B = 8'h47; #100;
A = 8'hB6; B = 8'h48; #100;
A = 8'hB6; B = 8'h49; #100;
A = 8'hB6; B = 8'h4A; #100;
A = 8'hB6; B = 8'h4B; #100;
A = 8'hB6; B = 8'h4C; #100;
A = 8'hB6; B = 8'h4D; #100;
A = 8'hB6; B = 8'h4E; #100;
A = 8'hB6; B = 8'h4F; #100;
A = 8'hB6; B = 8'h50; #100;
A = 8'hB6; B = 8'h51; #100;
A = 8'hB6; B = 8'h52; #100;
A = 8'hB6; B = 8'h53; #100;
A = 8'hB6; B = 8'h54; #100;
A = 8'hB6; B = 8'h55; #100;
A = 8'hB6; B = 8'h56; #100;
A = 8'hB6; B = 8'h57; #100;
A = 8'hB6; B = 8'h58; #100;
A = 8'hB6; B = 8'h59; #100;
A = 8'hB6; B = 8'h5A; #100;
A = 8'hB6; B = 8'h5B; #100;
A = 8'hB6; B = 8'h5C; #100;
A = 8'hB6; B = 8'h5D; #100;
A = 8'hB6; B = 8'h5E; #100;
A = 8'hB6; B = 8'h5F; #100;
A = 8'hB6; B = 8'h60; #100;
A = 8'hB6; B = 8'h61; #100;
A = 8'hB6; B = 8'h62; #100;
A = 8'hB6; B = 8'h63; #100;
A = 8'hB6; B = 8'h64; #100;
A = 8'hB6; B = 8'h65; #100;
A = 8'hB6; B = 8'h66; #100;
A = 8'hB6; B = 8'h67; #100;
A = 8'hB6; B = 8'h68; #100;
A = 8'hB6; B = 8'h69; #100;
A = 8'hB6; B = 8'h6A; #100;
A = 8'hB6; B = 8'h6B; #100;
A = 8'hB6; B = 8'h6C; #100;
A = 8'hB6; B = 8'h6D; #100;
A = 8'hB6; B = 8'h6E; #100;
A = 8'hB6; B = 8'h6F; #100;
A = 8'hB6; B = 8'h70; #100;
A = 8'hB6; B = 8'h71; #100;
A = 8'hB6; B = 8'h72; #100;
A = 8'hB6; B = 8'h73; #100;
A = 8'hB6; B = 8'h74; #100;
A = 8'hB6; B = 8'h75; #100;
A = 8'hB6; B = 8'h76; #100;
A = 8'hB6; B = 8'h77; #100;
A = 8'hB6; B = 8'h78; #100;
A = 8'hB6; B = 8'h79; #100;
A = 8'hB6; B = 8'h7A; #100;
A = 8'hB6; B = 8'h7B; #100;
A = 8'hB6; B = 8'h7C; #100;
A = 8'hB6; B = 8'h7D; #100;
A = 8'hB6; B = 8'h7E; #100;
A = 8'hB6; B = 8'h7F; #100;
A = 8'hB6; B = 8'h80; #100;
A = 8'hB6; B = 8'h81; #100;
A = 8'hB6; B = 8'h82; #100;
A = 8'hB6; B = 8'h83; #100;
A = 8'hB6; B = 8'h84; #100;
A = 8'hB6; B = 8'h85; #100;
A = 8'hB6; B = 8'h86; #100;
A = 8'hB6; B = 8'h87; #100;
A = 8'hB6; B = 8'h88; #100;
A = 8'hB6; B = 8'h89; #100;
A = 8'hB6; B = 8'h8A; #100;
A = 8'hB6; B = 8'h8B; #100;
A = 8'hB6; B = 8'h8C; #100;
A = 8'hB6; B = 8'h8D; #100;
A = 8'hB6; B = 8'h8E; #100;
A = 8'hB6; B = 8'h8F; #100;
A = 8'hB6; B = 8'h90; #100;
A = 8'hB6; B = 8'h91; #100;
A = 8'hB6; B = 8'h92; #100;
A = 8'hB6; B = 8'h93; #100;
A = 8'hB6; B = 8'h94; #100;
A = 8'hB6; B = 8'h95; #100;
A = 8'hB6; B = 8'h96; #100;
A = 8'hB6; B = 8'h97; #100;
A = 8'hB6; B = 8'h98; #100;
A = 8'hB6; B = 8'h99; #100;
A = 8'hB6; B = 8'h9A; #100;
A = 8'hB6; B = 8'h9B; #100;
A = 8'hB6; B = 8'h9C; #100;
A = 8'hB6; B = 8'h9D; #100;
A = 8'hB6; B = 8'h9E; #100;
A = 8'hB6; B = 8'h9F; #100;
A = 8'hB6; B = 8'hA0; #100;
A = 8'hB6; B = 8'hA1; #100;
A = 8'hB6; B = 8'hA2; #100;
A = 8'hB6; B = 8'hA3; #100;
A = 8'hB6; B = 8'hA4; #100;
A = 8'hB6; B = 8'hA5; #100;
A = 8'hB6; B = 8'hA6; #100;
A = 8'hB6; B = 8'hA7; #100;
A = 8'hB6; B = 8'hA8; #100;
A = 8'hB6; B = 8'hA9; #100;
A = 8'hB6; B = 8'hAA; #100;
A = 8'hB6; B = 8'hAB; #100;
A = 8'hB6; B = 8'hAC; #100;
A = 8'hB6; B = 8'hAD; #100;
A = 8'hB6; B = 8'hAE; #100;
A = 8'hB6; B = 8'hAF; #100;
A = 8'hB6; B = 8'hB0; #100;
A = 8'hB6; B = 8'hB1; #100;
A = 8'hB6; B = 8'hB2; #100;
A = 8'hB6; B = 8'hB3; #100;
A = 8'hB6; B = 8'hB4; #100;
A = 8'hB6; B = 8'hB5; #100;
A = 8'hB6; B = 8'hB6; #100;
A = 8'hB6; B = 8'hB7; #100;
A = 8'hB6; B = 8'hB8; #100;
A = 8'hB6; B = 8'hB9; #100;
A = 8'hB6; B = 8'hBA; #100;
A = 8'hB6; B = 8'hBB; #100;
A = 8'hB6; B = 8'hBC; #100;
A = 8'hB6; B = 8'hBD; #100;
A = 8'hB6; B = 8'hBE; #100;
A = 8'hB6; B = 8'hBF; #100;
A = 8'hB6; B = 8'hC0; #100;
A = 8'hB6; B = 8'hC1; #100;
A = 8'hB6; B = 8'hC2; #100;
A = 8'hB6; B = 8'hC3; #100;
A = 8'hB6; B = 8'hC4; #100;
A = 8'hB6; B = 8'hC5; #100;
A = 8'hB6; B = 8'hC6; #100;
A = 8'hB6; B = 8'hC7; #100;
A = 8'hB6; B = 8'hC8; #100;
A = 8'hB6; B = 8'hC9; #100;
A = 8'hB6; B = 8'hCA; #100;
A = 8'hB6; B = 8'hCB; #100;
A = 8'hB6; B = 8'hCC; #100;
A = 8'hB6; B = 8'hCD; #100;
A = 8'hB6; B = 8'hCE; #100;
A = 8'hB6; B = 8'hCF; #100;
A = 8'hB6; B = 8'hD0; #100;
A = 8'hB6; B = 8'hD1; #100;
A = 8'hB6; B = 8'hD2; #100;
A = 8'hB6; B = 8'hD3; #100;
A = 8'hB6; B = 8'hD4; #100;
A = 8'hB6; B = 8'hD5; #100;
A = 8'hB6; B = 8'hD6; #100;
A = 8'hB6; B = 8'hD7; #100;
A = 8'hB6; B = 8'hD8; #100;
A = 8'hB6; B = 8'hD9; #100;
A = 8'hB6; B = 8'hDA; #100;
A = 8'hB6; B = 8'hDB; #100;
A = 8'hB6; B = 8'hDC; #100;
A = 8'hB6; B = 8'hDD; #100;
A = 8'hB6; B = 8'hDE; #100;
A = 8'hB6; B = 8'hDF; #100;
A = 8'hB6; B = 8'hE0; #100;
A = 8'hB6; B = 8'hE1; #100;
A = 8'hB6; B = 8'hE2; #100;
A = 8'hB6; B = 8'hE3; #100;
A = 8'hB6; B = 8'hE4; #100;
A = 8'hB6; B = 8'hE5; #100;
A = 8'hB6; B = 8'hE6; #100;
A = 8'hB6; B = 8'hE7; #100;
A = 8'hB6; B = 8'hE8; #100;
A = 8'hB6; B = 8'hE9; #100;
A = 8'hB6; B = 8'hEA; #100;
A = 8'hB6; B = 8'hEB; #100;
A = 8'hB6; B = 8'hEC; #100;
A = 8'hB6; B = 8'hED; #100;
A = 8'hB6; B = 8'hEE; #100;
A = 8'hB6; B = 8'hEF; #100;
A = 8'hB6; B = 8'hF0; #100;
A = 8'hB6; B = 8'hF1; #100;
A = 8'hB6; B = 8'hF2; #100;
A = 8'hB6; B = 8'hF3; #100;
A = 8'hB6; B = 8'hF4; #100;
A = 8'hB6; B = 8'hF5; #100;
A = 8'hB6; B = 8'hF6; #100;
A = 8'hB6; B = 8'hF7; #100;
A = 8'hB6; B = 8'hF8; #100;
A = 8'hB6; B = 8'hF9; #100;
A = 8'hB6; B = 8'hFA; #100;
A = 8'hB6; B = 8'hFB; #100;
A = 8'hB6; B = 8'hFC; #100;
A = 8'hB6; B = 8'hFD; #100;
A = 8'hB6; B = 8'hFE; #100;
A = 8'hB6; B = 8'hFF; #100;
A = 8'hB7; B = 8'h0; #100;
A = 8'hB7; B = 8'h1; #100;
A = 8'hB7; B = 8'h2; #100;
A = 8'hB7; B = 8'h3; #100;
A = 8'hB7; B = 8'h4; #100;
A = 8'hB7; B = 8'h5; #100;
A = 8'hB7; B = 8'h6; #100;
A = 8'hB7; B = 8'h7; #100;
A = 8'hB7; B = 8'h8; #100;
A = 8'hB7; B = 8'h9; #100;
A = 8'hB7; B = 8'hA; #100;
A = 8'hB7; B = 8'hB; #100;
A = 8'hB7; B = 8'hC; #100;
A = 8'hB7; B = 8'hD; #100;
A = 8'hB7; B = 8'hE; #100;
A = 8'hB7; B = 8'hF; #100;
A = 8'hB7; B = 8'h10; #100;
A = 8'hB7; B = 8'h11; #100;
A = 8'hB7; B = 8'h12; #100;
A = 8'hB7; B = 8'h13; #100;
A = 8'hB7; B = 8'h14; #100;
A = 8'hB7; B = 8'h15; #100;
A = 8'hB7; B = 8'h16; #100;
A = 8'hB7; B = 8'h17; #100;
A = 8'hB7; B = 8'h18; #100;
A = 8'hB7; B = 8'h19; #100;
A = 8'hB7; B = 8'h1A; #100;
A = 8'hB7; B = 8'h1B; #100;
A = 8'hB7; B = 8'h1C; #100;
A = 8'hB7; B = 8'h1D; #100;
A = 8'hB7; B = 8'h1E; #100;
A = 8'hB7; B = 8'h1F; #100;
A = 8'hB7; B = 8'h20; #100;
A = 8'hB7; B = 8'h21; #100;
A = 8'hB7; B = 8'h22; #100;
A = 8'hB7; B = 8'h23; #100;
A = 8'hB7; B = 8'h24; #100;
A = 8'hB7; B = 8'h25; #100;
A = 8'hB7; B = 8'h26; #100;
A = 8'hB7; B = 8'h27; #100;
A = 8'hB7; B = 8'h28; #100;
A = 8'hB7; B = 8'h29; #100;
A = 8'hB7; B = 8'h2A; #100;
A = 8'hB7; B = 8'h2B; #100;
A = 8'hB7; B = 8'h2C; #100;
A = 8'hB7; B = 8'h2D; #100;
A = 8'hB7; B = 8'h2E; #100;
A = 8'hB7; B = 8'h2F; #100;
A = 8'hB7; B = 8'h30; #100;
A = 8'hB7; B = 8'h31; #100;
A = 8'hB7; B = 8'h32; #100;
A = 8'hB7; B = 8'h33; #100;
A = 8'hB7; B = 8'h34; #100;
A = 8'hB7; B = 8'h35; #100;
A = 8'hB7; B = 8'h36; #100;
A = 8'hB7; B = 8'h37; #100;
A = 8'hB7; B = 8'h38; #100;
A = 8'hB7; B = 8'h39; #100;
A = 8'hB7; B = 8'h3A; #100;
A = 8'hB7; B = 8'h3B; #100;
A = 8'hB7; B = 8'h3C; #100;
A = 8'hB7; B = 8'h3D; #100;
A = 8'hB7; B = 8'h3E; #100;
A = 8'hB7; B = 8'h3F; #100;
A = 8'hB7; B = 8'h40; #100;
A = 8'hB7; B = 8'h41; #100;
A = 8'hB7; B = 8'h42; #100;
A = 8'hB7; B = 8'h43; #100;
A = 8'hB7; B = 8'h44; #100;
A = 8'hB7; B = 8'h45; #100;
A = 8'hB7; B = 8'h46; #100;
A = 8'hB7; B = 8'h47; #100;
A = 8'hB7; B = 8'h48; #100;
A = 8'hB7; B = 8'h49; #100;
A = 8'hB7; B = 8'h4A; #100;
A = 8'hB7; B = 8'h4B; #100;
A = 8'hB7; B = 8'h4C; #100;
A = 8'hB7; B = 8'h4D; #100;
A = 8'hB7; B = 8'h4E; #100;
A = 8'hB7; B = 8'h4F; #100;
A = 8'hB7; B = 8'h50; #100;
A = 8'hB7; B = 8'h51; #100;
A = 8'hB7; B = 8'h52; #100;
A = 8'hB7; B = 8'h53; #100;
A = 8'hB7; B = 8'h54; #100;
A = 8'hB7; B = 8'h55; #100;
A = 8'hB7; B = 8'h56; #100;
A = 8'hB7; B = 8'h57; #100;
A = 8'hB7; B = 8'h58; #100;
A = 8'hB7; B = 8'h59; #100;
A = 8'hB7; B = 8'h5A; #100;
A = 8'hB7; B = 8'h5B; #100;
A = 8'hB7; B = 8'h5C; #100;
A = 8'hB7; B = 8'h5D; #100;
A = 8'hB7; B = 8'h5E; #100;
A = 8'hB7; B = 8'h5F; #100;
A = 8'hB7; B = 8'h60; #100;
A = 8'hB7; B = 8'h61; #100;
A = 8'hB7; B = 8'h62; #100;
A = 8'hB7; B = 8'h63; #100;
A = 8'hB7; B = 8'h64; #100;
A = 8'hB7; B = 8'h65; #100;
A = 8'hB7; B = 8'h66; #100;
A = 8'hB7; B = 8'h67; #100;
A = 8'hB7; B = 8'h68; #100;
A = 8'hB7; B = 8'h69; #100;
A = 8'hB7; B = 8'h6A; #100;
A = 8'hB7; B = 8'h6B; #100;
A = 8'hB7; B = 8'h6C; #100;
A = 8'hB7; B = 8'h6D; #100;
A = 8'hB7; B = 8'h6E; #100;
A = 8'hB7; B = 8'h6F; #100;
A = 8'hB7; B = 8'h70; #100;
A = 8'hB7; B = 8'h71; #100;
A = 8'hB7; B = 8'h72; #100;
A = 8'hB7; B = 8'h73; #100;
A = 8'hB7; B = 8'h74; #100;
A = 8'hB7; B = 8'h75; #100;
A = 8'hB7; B = 8'h76; #100;
A = 8'hB7; B = 8'h77; #100;
A = 8'hB7; B = 8'h78; #100;
A = 8'hB7; B = 8'h79; #100;
A = 8'hB7; B = 8'h7A; #100;
A = 8'hB7; B = 8'h7B; #100;
A = 8'hB7; B = 8'h7C; #100;
A = 8'hB7; B = 8'h7D; #100;
A = 8'hB7; B = 8'h7E; #100;
A = 8'hB7; B = 8'h7F; #100;
A = 8'hB7; B = 8'h80; #100;
A = 8'hB7; B = 8'h81; #100;
A = 8'hB7; B = 8'h82; #100;
A = 8'hB7; B = 8'h83; #100;
A = 8'hB7; B = 8'h84; #100;
A = 8'hB7; B = 8'h85; #100;
A = 8'hB7; B = 8'h86; #100;
A = 8'hB7; B = 8'h87; #100;
A = 8'hB7; B = 8'h88; #100;
A = 8'hB7; B = 8'h89; #100;
A = 8'hB7; B = 8'h8A; #100;
A = 8'hB7; B = 8'h8B; #100;
A = 8'hB7; B = 8'h8C; #100;
A = 8'hB7; B = 8'h8D; #100;
A = 8'hB7; B = 8'h8E; #100;
A = 8'hB7; B = 8'h8F; #100;
A = 8'hB7; B = 8'h90; #100;
A = 8'hB7; B = 8'h91; #100;
A = 8'hB7; B = 8'h92; #100;
A = 8'hB7; B = 8'h93; #100;
A = 8'hB7; B = 8'h94; #100;
A = 8'hB7; B = 8'h95; #100;
A = 8'hB7; B = 8'h96; #100;
A = 8'hB7; B = 8'h97; #100;
A = 8'hB7; B = 8'h98; #100;
A = 8'hB7; B = 8'h99; #100;
A = 8'hB7; B = 8'h9A; #100;
A = 8'hB7; B = 8'h9B; #100;
A = 8'hB7; B = 8'h9C; #100;
A = 8'hB7; B = 8'h9D; #100;
A = 8'hB7; B = 8'h9E; #100;
A = 8'hB7; B = 8'h9F; #100;
A = 8'hB7; B = 8'hA0; #100;
A = 8'hB7; B = 8'hA1; #100;
A = 8'hB7; B = 8'hA2; #100;
A = 8'hB7; B = 8'hA3; #100;
A = 8'hB7; B = 8'hA4; #100;
A = 8'hB7; B = 8'hA5; #100;
A = 8'hB7; B = 8'hA6; #100;
A = 8'hB7; B = 8'hA7; #100;
A = 8'hB7; B = 8'hA8; #100;
A = 8'hB7; B = 8'hA9; #100;
A = 8'hB7; B = 8'hAA; #100;
A = 8'hB7; B = 8'hAB; #100;
A = 8'hB7; B = 8'hAC; #100;
A = 8'hB7; B = 8'hAD; #100;
A = 8'hB7; B = 8'hAE; #100;
A = 8'hB7; B = 8'hAF; #100;
A = 8'hB7; B = 8'hB0; #100;
A = 8'hB7; B = 8'hB1; #100;
A = 8'hB7; B = 8'hB2; #100;
A = 8'hB7; B = 8'hB3; #100;
A = 8'hB7; B = 8'hB4; #100;
A = 8'hB7; B = 8'hB5; #100;
A = 8'hB7; B = 8'hB6; #100;
A = 8'hB7; B = 8'hB7; #100;
A = 8'hB7; B = 8'hB8; #100;
A = 8'hB7; B = 8'hB9; #100;
A = 8'hB7; B = 8'hBA; #100;
A = 8'hB7; B = 8'hBB; #100;
A = 8'hB7; B = 8'hBC; #100;
A = 8'hB7; B = 8'hBD; #100;
A = 8'hB7; B = 8'hBE; #100;
A = 8'hB7; B = 8'hBF; #100;
A = 8'hB7; B = 8'hC0; #100;
A = 8'hB7; B = 8'hC1; #100;
A = 8'hB7; B = 8'hC2; #100;
A = 8'hB7; B = 8'hC3; #100;
A = 8'hB7; B = 8'hC4; #100;
A = 8'hB7; B = 8'hC5; #100;
A = 8'hB7; B = 8'hC6; #100;
A = 8'hB7; B = 8'hC7; #100;
A = 8'hB7; B = 8'hC8; #100;
A = 8'hB7; B = 8'hC9; #100;
A = 8'hB7; B = 8'hCA; #100;
A = 8'hB7; B = 8'hCB; #100;
A = 8'hB7; B = 8'hCC; #100;
A = 8'hB7; B = 8'hCD; #100;
A = 8'hB7; B = 8'hCE; #100;
A = 8'hB7; B = 8'hCF; #100;
A = 8'hB7; B = 8'hD0; #100;
A = 8'hB7; B = 8'hD1; #100;
A = 8'hB7; B = 8'hD2; #100;
A = 8'hB7; B = 8'hD3; #100;
A = 8'hB7; B = 8'hD4; #100;
A = 8'hB7; B = 8'hD5; #100;
A = 8'hB7; B = 8'hD6; #100;
A = 8'hB7; B = 8'hD7; #100;
A = 8'hB7; B = 8'hD8; #100;
A = 8'hB7; B = 8'hD9; #100;
A = 8'hB7; B = 8'hDA; #100;
A = 8'hB7; B = 8'hDB; #100;
A = 8'hB7; B = 8'hDC; #100;
A = 8'hB7; B = 8'hDD; #100;
A = 8'hB7; B = 8'hDE; #100;
A = 8'hB7; B = 8'hDF; #100;
A = 8'hB7; B = 8'hE0; #100;
A = 8'hB7; B = 8'hE1; #100;
A = 8'hB7; B = 8'hE2; #100;
A = 8'hB7; B = 8'hE3; #100;
A = 8'hB7; B = 8'hE4; #100;
A = 8'hB7; B = 8'hE5; #100;
A = 8'hB7; B = 8'hE6; #100;
A = 8'hB7; B = 8'hE7; #100;
A = 8'hB7; B = 8'hE8; #100;
A = 8'hB7; B = 8'hE9; #100;
A = 8'hB7; B = 8'hEA; #100;
A = 8'hB7; B = 8'hEB; #100;
A = 8'hB7; B = 8'hEC; #100;
A = 8'hB7; B = 8'hED; #100;
A = 8'hB7; B = 8'hEE; #100;
A = 8'hB7; B = 8'hEF; #100;
A = 8'hB7; B = 8'hF0; #100;
A = 8'hB7; B = 8'hF1; #100;
A = 8'hB7; B = 8'hF2; #100;
A = 8'hB7; B = 8'hF3; #100;
A = 8'hB7; B = 8'hF4; #100;
A = 8'hB7; B = 8'hF5; #100;
A = 8'hB7; B = 8'hF6; #100;
A = 8'hB7; B = 8'hF7; #100;
A = 8'hB7; B = 8'hF8; #100;
A = 8'hB7; B = 8'hF9; #100;
A = 8'hB7; B = 8'hFA; #100;
A = 8'hB7; B = 8'hFB; #100;
A = 8'hB7; B = 8'hFC; #100;
A = 8'hB7; B = 8'hFD; #100;
A = 8'hB7; B = 8'hFE; #100;
A = 8'hB7; B = 8'hFF; #100;
A = 8'hB8; B = 8'h0; #100;
A = 8'hB8; B = 8'h1; #100;
A = 8'hB8; B = 8'h2; #100;
A = 8'hB8; B = 8'h3; #100;
A = 8'hB8; B = 8'h4; #100;
A = 8'hB8; B = 8'h5; #100;
A = 8'hB8; B = 8'h6; #100;
A = 8'hB8; B = 8'h7; #100;
A = 8'hB8; B = 8'h8; #100;
A = 8'hB8; B = 8'h9; #100;
A = 8'hB8; B = 8'hA; #100;
A = 8'hB8; B = 8'hB; #100;
A = 8'hB8; B = 8'hC; #100;
A = 8'hB8; B = 8'hD; #100;
A = 8'hB8; B = 8'hE; #100;
A = 8'hB8; B = 8'hF; #100;
A = 8'hB8; B = 8'h10; #100;
A = 8'hB8; B = 8'h11; #100;
A = 8'hB8; B = 8'h12; #100;
A = 8'hB8; B = 8'h13; #100;
A = 8'hB8; B = 8'h14; #100;
A = 8'hB8; B = 8'h15; #100;
A = 8'hB8; B = 8'h16; #100;
A = 8'hB8; B = 8'h17; #100;
A = 8'hB8; B = 8'h18; #100;
A = 8'hB8; B = 8'h19; #100;
A = 8'hB8; B = 8'h1A; #100;
A = 8'hB8; B = 8'h1B; #100;
A = 8'hB8; B = 8'h1C; #100;
A = 8'hB8; B = 8'h1D; #100;
A = 8'hB8; B = 8'h1E; #100;
A = 8'hB8; B = 8'h1F; #100;
A = 8'hB8; B = 8'h20; #100;
A = 8'hB8; B = 8'h21; #100;
A = 8'hB8; B = 8'h22; #100;
A = 8'hB8; B = 8'h23; #100;
A = 8'hB8; B = 8'h24; #100;
A = 8'hB8; B = 8'h25; #100;
A = 8'hB8; B = 8'h26; #100;
A = 8'hB8; B = 8'h27; #100;
A = 8'hB8; B = 8'h28; #100;
A = 8'hB8; B = 8'h29; #100;
A = 8'hB8; B = 8'h2A; #100;
A = 8'hB8; B = 8'h2B; #100;
A = 8'hB8; B = 8'h2C; #100;
A = 8'hB8; B = 8'h2D; #100;
A = 8'hB8; B = 8'h2E; #100;
A = 8'hB8; B = 8'h2F; #100;
A = 8'hB8; B = 8'h30; #100;
A = 8'hB8; B = 8'h31; #100;
A = 8'hB8; B = 8'h32; #100;
A = 8'hB8; B = 8'h33; #100;
A = 8'hB8; B = 8'h34; #100;
A = 8'hB8; B = 8'h35; #100;
A = 8'hB8; B = 8'h36; #100;
A = 8'hB8; B = 8'h37; #100;
A = 8'hB8; B = 8'h38; #100;
A = 8'hB8; B = 8'h39; #100;
A = 8'hB8; B = 8'h3A; #100;
A = 8'hB8; B = 8'h3B; #100;
A = 8'hB8; B = 8'h3C; #100;
A = 8'hB8; B = 8'h3D; #100;
A = 8'hB8; B = 8'h3E; #100;
A = 8'hB8; B = 8'h3F; #100;
A = 8'hB8; B = 8'h40; #100;
A = 8'hB8; B = 8'h41; #100;
A = 8'hB8; B = 8'h42; #100;
A = 8'hB8; B = 8'h43; #100;
A = 8'hB8; B = 8'h44; #100;
A = 8'hB8; B = 8'h45; #100;
A = 8'hB8; B = 8'h46; #100;
A = 8'hB8; B = 8'h47; #100;
A = 8'hB8; B = 8'h48; #100;
A = 8'hB8; B = 8'h49; #100;
A = 8'hB8; B = 8'h4A; #100;
A = 8'hB8; B = 8'h4B; #100;
A = 8'hB8; B = 8'h4C; #100;
A = 8'hB8; B = 8'h4D; #100;
A = 8'hB8; B = 8'h4E; #100;
A = 8'hB8; B = 8'h4F; #100;
A = 8'hB8; B = 8'h50; #100;
A = 8'hB8; B = 8'h51; #100;
A = 8'hB8; B = 8'h52; #100;
A = 8'hB8; B = 8'h53; #100;
A = 8'hB8; B = 8'h54; #100;
A = 8'hB8; B = 8'h55; #100;
A = 8'hB8; B = 8'h56; #100;
A = 8'hB8; B = 8'h57; #100;
A = 8'hB8; B = 8'h58; #100;
A = 8'hB8; B = 8'h59; #100;
A = 8'hB8; B = 8'h5A; #100;
A = 8'hB8; B = 8'h5B; #100;
A = 8'hB8; B = 8'h5C; #100;
A = 8'hB8; B = 8'h5D; #100;
A = 8'hB8; B = 8'h5E; #100;
A = 8'hB8; B = 8'h5F; #100;
A = 8'hB8; B = 8'h60; #100;
A = 8'hB8; B = 8'h61; #100;
A = 8'hB8; B = 8'h62; #100;
A = 8'hB8; B = 8'h63; #100;
A = 8'hB8; B = 8'h64; #100;
A = 8'hB8; B = 8'h65; #100;
A = 8'hB8; B = 8'h66; #100;
A = 8'hB8; B = 8'h67; #100;
A = 8'hB8; B = 8'h68; #100;
A = 8'hB8; B = 8'h69; #100;
A = 8'hB8; B = 8'h6A; #100;
A = 8'hB8; B = 8'h6B; #100;
A = 8'hB8; B = 8'h6C; #100;
A = 8'hB8; B = 8'h6D; #100;
A = 8'hB8; B = 8'h6E; #100;
A = 8'hB8; B = 8'h6F; #100;
A = 8'hB8; B = 8'h70; #100;
A = 8'hB8; B = 8'h71; #100;
A = 8'hB8; B = 8'h72; #100;
A = 8'hB8; B = 8'h73; #100;
A = 8'hB8; B = 8'h74; #100;
A = 8'hB8; B = 8'h75; #100;
A = 8'hB8; B = 8'h76; #100;
A = 8'hB8; B = 8'h77; #100;
A = 8'hB8; B = 8'h78; #100;
A = 8'hB8; B = 8'h79; #100;
A = 8'hB8; B = 8'h7A; #100;
A = 8'hB8; B = 8'h7B; #100;
A = 8'hB8; B = 8'h7C; #100;
A = 8'hB8; B = 8'h7D; #100;
A = 8'hB8; B = 8'h7E; #100;
A = 8'hB8; B = 8'h7F; #100;
A = 8'hB8; B = 8'h80; #100;
A = 8'hB8; B = 8'h81; #100;
A = 8'hB8; B = 8'h82; #100;
A = 8'hB8; B = 8'h83; #100;
A = 8'hB8; B = 8'h84; #100;
A = 8'hB8; B = 8'h85; #100;
A = 8'hB8; B = 8'h86; #100;
A = 8'hB8; B = 8'h87; #100;
A = 8'hB8; B = 8'h88; #100;
A = 8'hB8; B = 8'h89; #100;
A = 8'hB8; B = 8'h8A; #100;
A = 8'hB8; B = 8'h8B; #100;
A = 8'hB8; B = 8'h8C; #100;
A = 8'hB8; B = 8'h8D; #100;
A = 8'hB8; B = 8'h8E; #100;
A = 8'hB8; B = 8'h8F; #100;
A = 8'hB8; B = 8'h90; #100;
A = 8'hB8; B = 8'h91; #100;
A = 8'hB8; B = 8'h92; #100;
A = 8'hB8; B = 8'h93; #100;
A = 8'hB8; B = 8'h94; #100;
A = 8'hB8; B = 8'h95; #100;
A = 8'hB8; B = 8'h96; #100;
A = 8'hB8; B = 8'h97; #100;
A = 8'hB8; B = 8'h98; #100;
A = 8'hB8; B = 8'h99; #100;
A = 8'hB8; B = 8'h9A; #100;
A = 8'hB8; B = 8'h9B; #100;
A = 8'hB8; B = 8'h9C; #100;
A = 8'hB8; B = 8'h9D; #100;
A = 8'hB8; B = 8'h9E; #100;
A = 8'hB8; B = 8'h9F; #100;
A = 8'hB8; B = 8'hA0; #100;
A = 8'hB8; B = 8'hA1; #100;
A = 8'hB8; B = 8'hA2; #100;
A = 8'hB8; B = 8'hA3; #100;
A = 8'hB8; B = 8'hA4; #100;
A = 8'hB8; B = 8'hA5; #100;
A = 8'hB8; B = 8'hA6; #100;
A = 8'hB8; B = 8'hA7; #100;
A = 8'hB8; B = 8'hA8; #100;
A = 8'hB8; B = 8'hA9; #100;
A = 8'hB8; B = 8'hAA; #100;
A = 8'hB8; B = 8'hAB; #100;
A = 8'hB8; B = 8'hAC; #100;
A = 8'hB8; B = 8'hAD; #100;
A = 8'hB8; B = 8'hAE; #100;
A = 8'hB8; B = 8'hAF; #100;
A = 8'hB8; B = 8'hB0; #100;
A = 8'hB8; B = 8'hB1; #100;
A = 8'hB8; B = 8'hB2; #100;
A = 8'hB8; B = 8'hB3; #100;
A = 8'hB8; B = 8'hB4; #100;
A = 8'hB8; B = 8'hB5; #100;
A = 8'hB8; B = 8'hB6; #100;
A = 8'hB8; B = 8'hB7; #100;
A = 8'hB8; B = 8'hB8; #100;
A = 8'hB8; B = 8'hB9; #100;
A = 8'hB8; B = 8'hBA; #100;
A = 8'hB8; B = 8'hBB; #100;
A = 8'hB8; B = 8'hBC; #100;
A = 8'hB8; B = 8'hBD; #100;
A = 8'hB8; B = 8'hBE; #100;
A = 8'hB8; B = 8'hBF; #100;
A = 8'hB8; B = 8'hC0; #100;
A = 8'hB8; B = 8'hC1; #100;
A = 8'hB8; B = 8'hC2; #100;
A = 8'hB8; B = 8'hC3; #100;
A = 8'hB8; B = 8'hC4; #100;
A = 8'hB8; B = 8'hC5; #100;
A = 8'hB8; B = 8'hC6; #100;
A = 8'hB8; B = 8'hC7; #100;
A = 8'hB8; B = 8'hC8; #100;
A = 8'hB8; B = 8'hC9; #100;
A = 8'hB8; B = 8'hCA; #100;
A = 8'hB8; B = 8'hCB; #100;
A = 8'hB8; B = 8'hCC; #100;
A = 8'hB8; B = 8'hCD; #100;
A = 8'hB8; B = 8'hCE; #100;
A = 8'hB8; B = 8'hCF; #100;
A = 8'hB8; B = 8'hD0; #100;
A = 8'hB8; B = 8'hD1; #100;
A = 8'hB8; B = 8'hD2; #100;
A = 8'hB8; B = 8'hD3; #100;
A = 8'hB8; B = 8'hD4; #100;
A = 8'hB8; B = 8'hD5; #100;
A = 8'hB8; B = 8'hD6; #100;
A = 8'hB8; B = 8'hD7; #100;
A = 8'hB8; B = 8'hD8; #100;
A = 8'hB8; B = 8'hD9; #100;
A = 8'hB8; B = 8'hDA; #100;
A = 8'hB8; B = 8'hDB; #100;
A = 8'hB8; B = 8'hDC; #100;
A = 8'hB8; B = 8'hDD; #100;
A = 8'hB8; B = 8'hDE; #100;
A = 8'hB8; B = 8'hDF; #100;
A = 8'hB8; B = 8'hE0; #100;
A = 8'hB8; B = 8'hE1; #100;
A = 8'hB8; B = 8'hE2; #100;
A = 8'hB8; B = 8'hE3; #100;
A = 8'hB8; B = 8'hE4; #100;
A = 8'hB8; B = 8'hE5; #100;
A = 8'hB8; B = 8'hE6; #100;
A = 8'hB8; B = 8'hE7; #100;
A = 8'hB8; B = 8'hE8; #100;
A = 8'hB8; B = 8'hE9; #100;
A = 8'hB8; B = 8'hEA; #100;
A = 8'hB8; B = 8'hEB; #100;
A = 8'hB8; B = 8'hEC; #100;
A = 8'hB8; B = 8'hED; #100;
A = 8'hB8; B = 8'hEE; #100;
A = 8'hB8; B = 8'hEF; #100;
A = 8'hB8; B = 8'hF0; #100;
A = 8'hB8; B = 8'hF1; #100;
A = 8'hB8; B = 8'hF2; #100;
A = 8'hB8; B = 8'hF3; #100;
A = 8'hB8; B = 8'hF4; #100;
A = 8'hB8; B = 8'hF5; #100;
A = 8'hB8; B = 8'hF6; #100;
A = 8'hB8; B = 8'hF7; #100;
A = 8'hB8; B = 8'hF8; #100;
A = 8'hB8; B = 8'hF9; #100;
A = 8'hB8; B = 8'hFA; #100;
A = 8'hB8; B = 8'hFB; #100;
A = 8'hB8; B = 8'hFC; #100;
A = 8'hB8; B = 8'hFD; #100;
A = 8'hB8; B = 8'hFE; #100;
A = 8'hB8; B = 8'hFF; #100;
A = 8'hB9; B = 8'h0; #100;
A = 8'hB9; B = 8'h1; #100;
A = 8'hB9; B = 8'h2; #100;
A = 8'hB9; B = 8'h3; #100;
A = 8'hB9; B = 8'h4; #100;
A = 8'hB9; B = 8'h5; #100;
A = 8'hB9; B = 8'h6; #100;
A = 8'hB9; B = 8'h7; #100;
A = 8'hB9; B = 8'h8; #100;
A = 8'hB9; B = 8'h9; #100;
A = 8'hB9; B = 8'hA; #100;
A = 8'hB9; B = 8'hB; #100;
A = 8'hB9; B = 8'hC; #100;
A = 8'hB9; B = 8'hD; #100;
A = 8'hB9; B = 8'hE; #100;
A = 8'hB9; B = 8'hF; #100;
A = 8'hB9; B = 8'h10; #100;
A = 8'hB9; B = 8'h11; #100;
A = 8'hB9; B = 8'h12; #100;
A = 8'hB9; B = 8'h13; #100;
A = 8'hB9; B = 8'h14; #100;
A = 8'hB9; B = 8'h15; #100;
A = 8'hB9; B = 8'h16; #100;
A = 8'hB9; B = 8'h17; #100;
A = 8'hB9; B = 8'h18; #100;
A = 8'hB9; B = 8'h19; #100;
A = 8'hB9; B = 8'h1A; #100;
A = 8'hB9; B = 8'h1B; #100;
A = 8'hB9; B = 8'h1C; #100;
A = 8'hB9; B = 8'h1D; #100;
A = 8'hB9; B = 8'h1E; #100;
A = 8'hB9; B = 8'h1F; #100;
A = 8'hB9; B = 8'h20; #100;
A = 8'hB9; B = 8'h21; #100;
A = 8'hB9; B = 8'h22; #100;
A = 8'hB9; B = 8'h23; #100;
A = 8'hB9; B = 8'h24; #100;
A = 8'hB9; B = 8'h25; #100;
A = 8'hB9; B = 8'h26; #100;
A = 8'hB9; B = 8'h27; #100;
A = 8'hB9; B = 8'h28; #100;
A = 8'hB9; B = 8'h29; #100;
A = 8'hB9; B = 8'h2A; #100;
A = 8'hB9; B = 8'h2B; #100;
A = 8'hB9; B = 8'h2C; #100;
A = 8'hB9; B = 8'h2D; #100;
A = 8'hB9; B = 8'h2E; #100;
A = 8'hB9; B = 8'h2F; #100;
A = 8'hB9; B = 8'h30; #100;
A = 8'hB9; B = 8'h31; #100;
A = 8'hB9; B = 8'h32; #100;
A = 8'hB9; B = 8'h33; #100;
A = 8'hB9; B = 8'h34; #100;
A = 8'hB9; B = 8'h35; #100;
A = 8'hB9; B = 8'h36; #100;
A = 8'hB9; B = 8'h37; #100;
A = 8'hB9; B = 8'h38; #100;
A = 8'hB9; B = 8'h39; #100;
A = 8'hB9; B = 8'h3A; #100;
A = 8'hB9; B = 8'h3B; #100;
A = 8'hB9; B = 8'h3C; #100;
A = 8'hB9; B = 8'h3D; #100;
A = 8'hB9; B = 8'h3E; #100;
A = 8'hB9; B = 8'h3F; #100;
A = 8'hB9; B = 8'h40; #100;
A = 8'hB9; B = 8'h41; #100;
A = 8'hB9; B = 8'h42; #100;
A = 8'hB9; B = 8'h43; #100;
A = 8'hB9; B = 8'h44; #100;
A = 8'hB9; B = 8'h45; #100;
A = 8'hB9; B = 8'h46; #100;
A = 8'hB9; B = 8'h47; #100;
A = 8'hB9; B = 8'h48; #100;
A = 8'hB9; B = 8'h49; #100;
A = 8'hB9; B = 8'h4A; #100;
A = 8'hB9; B = 8'h4B; #100;
A = 8'hB9; B = 8'h4C; #100;
A = 8'hB9; B = 8'h4D; #100;
A = 8'hB9; B = 8'h4E; #100;
A = 8'hB9; B = 8'h4F; #100;
A = 8'hB9; B = 8'h50; #100;
A = 8'hB9; B = 8'h51; #100;
A = 8'hB9; B = 8'h52; #100;
A = 8'hB9; B = 8'h53; #100;
A = 8'hB9; B = 8'h54; #100;
A = 8'hB9; B = 8'h55; #100;
A = 8'hB9; B = 8'h56; #100;
A = 8'hB9; B = 8'h57; #100;
A = 8'hB9; B = 8'h58; #100;
A = 8'hB9; B = 8'h59; #100;
A = 8'hB9; B = 8'h5A; #100;
A = 8'hB9; B = 8'h5B; #100;
A = 8'hB9; B = 8'h5C; #100;
A = 8'hB9; B = 8'h5D; #100;
A = 8'hB9; B = 8'h5E; #100;
A = 8'hB9; B = 8'h5F; #100;
A = 8'hB9; B = 8'h60; #100;
A = 8'hB9; B = 8'h61; #100;
A = 8'hB9; B = 8'h62; #100;
A = 8'hB9; B = 8'h63; #100;
A = 8'hB9; B = 8'h64; #100;
A = 8'hB9; B = 8'h65; #100;
A = 8'hB9; B = 8'h66; #100;
A = 8'hB9; B = 8'h67; #100;
A = 8'hB9; B = 8'h68; #100;
A = 8'hB9; B = 8'h69; #100;
A = 8'hB9; B = 8'h6A; #100;
A = 8'hB9; B = 8'h6B; #100;
A = 8'hB9; B = 8'h6C; #100;
A = 8'hB9; B = 8'h6D; #100;
A = 8'hB9; B = 8'h6E; #100;
A = 8'hB9; B = 8'h6F; #100;
A = 8'hB9; B = 8'h70; #100;
A = 8'hB9; B = 8'h71; #100;
A = 8'hB9; B = 8'h72; #100;
A = 8'hB9; B = 8'h73; #100;
A = 8'hB9; B = 8'h74; #100;
A = 8'hB9; B = 8'h75; #100;
A = 8'hB9; B = 8'h76; #100;
A = 8'hB9; B = 8'h77; #100;
A = 8'hB9; B = 8'h78; #100;
A = 8'hB9; B = 8'h79; #100;
A = 8'hB9; B = 8'h7A; #100;
A = 8'hB9; B = 8'h7B; #100;
A = 8'hB9; B = 8'h7C; #100;
A = 8'hB9; B = 8'h7D; #100;
A = 8'hB9; B = 8'h7E; #100;
A = 8'hB9; B = 8'h7F; #100;
A = 8'hB9; B = 8'h80; #100;
A = 8'hB9; B = 8'h81; #100;
A = 8'hB9; B = 8'h82; #100;
A = 8'hB9; B = 8'h83; #100;
A = 8'hB9; B = 8'h84; #100;
A = 8'hB9; B = 8'h85; #100;
A = 8'hB9; B = 8'h86; #100;
A = 8'hB9; B = 8'h87; #100;
A = 8'hB9; B = 8'h88; #100;
A = 8'hB9; B = 8'h89; #100;
A = 8'hB9; B = 8'h8A; #100;
A = 8'hB9; B = 8'h8B; #100;
A = 8'hB9; B = 8'h8C; #100;
A = 8'hB9; B = 8'h8D; #100;
A = 8'hB9; B = 8'h8E; #100;
A = 8'hB9; B = 8'h8F; #100;
A = 8'hB9; B = 8'h90; #100;
A = 8'hB9; B = 8'h91; #100;
A = 8'hB9; B = 8'h92; #100;
A = 8'hB9; B = 8'h93; #100;
A = 8'hB9; B = 8'h94; #100;
A = 8'hB9; B = 8'h95; #100;
A = 8'hB9; B = 8'h96; #100;
A = 8'hB9; B = 8'h97; #100;
A = 8'hB9; B = 8'h98; #100;
A = 8'hB9; B = 8'h99; #100;
A = 8'hB9; B = 8'h9A; #100;
A = 8'hB9; B = 8'h9B; #100;
A = 8'hB9; B = 8'h9C; #100;
A = 8'hB9; B = 8'h9D; #100;
A = 8'hB9; B = 8'h9E; #100;
A = 8'hB9; B = 8'h9F; #100;
A = 8'hB9; B = 8'hA0; #100;
A = 8'hB9; B = 8'hA1; #100;
A = 8'hB9; B = 8'hA2; #100;
A = 8'hB9; B = 8'hA3; #100;
A = 8'hB9; B = 8'hA4; #100;
A = 8'hB9; B = 8'hA5; #100;
A = 8'hB9; B = 8'hA6; #100;
A = 8'hB9; B = 8'hA7; #100;
A = 8'hB9; B = 8'hA8; #100;
A = 8'hB9; B = 8'hA9; #100;
A = 8'hB9; B = 8'hAA; #100;
A = 8'hB9; B = 8'hAB; #100;
A = 8'hB9; B = 8'hAC; #100;
A = 8'hB9; B = 8'hAD; #100;
A = 8'hB9; B = 8'hAE; #100;
A = 8'hB9; B = 8'hAF; #100;
A = 8'hB9; B = 8'hB0; #100;
A = 8'hB9; B = 8'hB1; #100;
A = 8'hB9; B = 8'hB2; #100;
A = 8'hB9; B = 8'hB3; #100;
A = 8'hB9; B = 8'hB4; #100;
A = 8'hB9; B = 8'hB5; #100;
A = 8'hB9; B = 8'hB6; #100;
A = 8'hB9; B = 8'hB7; #100;
A = 8'hB9; B = 8'hB8; #100;
A = 8'hB9; B = 8'hB9; #100;
A = 8'hB9; B = 8'hBA; #100;
A = 8'hB9; B = 8'hBB; #100;
A = 8'hB9; B = 8'hBC; #100;
A = 8'hB9; B = 8'hBD; #100;
A = 8'hB9; B = 8'hBE; #100;
A = 8'hB9; B = 8'hBF; #100;
A = 8'hB9; B = 8'hC0; #100;
A = 8'hB9; B = 8'hC1; #100;
A = 8'hB9; B = 8'hC2; #100;
A = 8'hB9; B = 8'hC3; #100;
A = 8'hB9; B = 8'hC4; #100;
A = 8'hB9; B = 8'hC5; #100;
A = 8'hB9; B = 8'hC6; #100;
A = 8'hB9; B = 8'hC7; #100;
A = 8'hB9; B = 8'hC8; #100;
A = 8'hB9; B = 8'hC9; #100;
A = 8'hB9; B = 8'hCA; #100;
A = 8'hB9; B = 8'hCB; #100;
A = 8'hB9; B = 8'hCC; #100;
A = 8'hB9; B = 8'hCD; #100;
A = 8'hB9; B = 8'hCE; #100;
A = 8'hB9; B = 8'hCF; #100;
A = 8'hB9; B = 8'hD0; #100;
A = 8'hB9; B = 8'hD1; #100;
A = 8'hB9; B = 8'hD2; #100;
A = 8'hB9; B = 8'hD3; #100;
A = 8'hB9; B = 8'hD4; #100;
A = 8'hB9; B = 8'hD5; #100;
A = 8'hB9; B = 8'hD6; #100;
A = 8'hB9; B = 8'hD7; #100;
A = 8'hB9; B = 8'hD8; #100;
A = 8'hB9; B = 8'hD9; #100;
A = 8'hB9; B = 8'hDA; #100;
A = 8'hB9; B = 8'hDB; #100;
A = 8'hB9; B = 8'hDC; #100;
A = 8'hB9; B = 8'hDD; #100;
A = 8'hB9; B = 8'hDE; #100;
A = 8'hB9; B = 8'hDF; #100;
A = 8'hB9; B = 8'hE0; #100;
A = 8'hB9; B = 8'hE1; #100;
A = 8'hB9; B = 8'hE2; #100;
A = 8'hB9; B = 8'hE3; #100;
A = 8'hB9; B = 8'hE4; #100;
A = 8'hB9; B = 8'hE5; #100;
A = 8'hB9; B = 8'hE6; #100;
A = 8'hB9; B = 8'hE7; #100;
A = 8'hB9; B = 8'hE8; #100;
A = 8'hB9; B = 8'hE9; #100;
A = 8'hB9; B = 8'hEA; #100;
A = 8'hB9; B = 8'hEB; #100;
A = 8'hB9; B = 8'hEC; #100;
A = 8'hB9; B = 8'hED; #100;
A = 8'hB9; B = 8'hEE; #100;
A = 8'hB9; B = 8'hEF; #100;
A = 8'hB9; B = 8'hF0; #100;
A = 8'hB9; B = 8'hF1; #100;
A = 8'hB9; B = 8'hF2; #100;
A = 8'hB9; B = 8'hF3; #100;
A = 8'hB9; B = 8'hF4; #100;
A = 8'hB9; B = 8'hF5; #100;
A = 8'hB9; B = 8'hF6; #100;
A = 8'hB9; B = 8'hF7; #100;
A = 8'hB9; B = 8'hF8; #100;
A = 8'hB9; B = 8'hF9; #100;
A = 8'hB9; B = 8'hFA; #100;
A = 8'hB9; B = 8'hFB; #100;
A = 8'hB9; B = 8'hFC; #100;
A = 8'hB9; B = 8'hFD; #100;
A = 8'hB9; B = 8'hFE; #100;
A = 8'hB9; B = 8'hFF; #100;
A = 8'hBA; B = 8'h0; #100;
A = 8'hBA; B = 8'h1; #100;
A = 8'hBA; B = 8'h2; #100;
A = 8'hBA; B = 8'h3; #100;
A = 8'hBA; B = 8'h4; #100;
A = 8'hBA; B = 8'h5; #100;
A = 8'hBA; B = 8'h6; #100;
A = 8'hBA; B = 8'h7; #100;
A = 8'hBA; B = 8'h8; #100;
A = 8'hBA; B = 8'h9; #100;
A = 8'hBA; B = 8'hA; #100;
A = 8'hBA; B = 8'hB; #100;
A = 8'hBA; B = 8'hC; #100;
A = 8'hBA; B = 8'hD; #100;
A = 8'hBA; B = 8'hE; #100;
A = 8'hBA; B = 8'hF; #100;
A = 8'hBA; B = 8'h10; #100;
A = 8'hBA; B = 8'h11; #100;
A = 8'hBA; B = 8'h12; #100;
A = 8'hBA; B = 8'h13; #100;
A = 8'hBA; B = 8'h14; #100;
A = 8'hBA; B = 8'h15; #100;
A = 8'hBA; B = 8'h16; #100;
A = 8'hBA; B = 8'h17; #100;
A = 8'hBA; B = 8'h18; #100;
A = 8'hBA; B = 8'h19; #100;
A = 8'hBA; B = 8'h1A; #100;
A = 8'hBA; B = 8'h1B; #100;
A = 8'hBA; B = 8'h1C; #100;
A = 8'hBA; B = 8'h1D; #100;
A = 8'hBA; B = 8'h1E; #100;
A = 8'hBA; B = 8'h1F; #100;
A = 8'hBA; B = 8'h20; #100;
A = 8'hBA; B = 8'h21; #100;
A = 8'hBA; B = 8'h22; #100;
A = 8'hBA; B = 8'h23; #100;
A = 8'hBA; B = 8'h24; #100;
A = 8'hBA; B = 8'h25; #100;
A = 8'hBA; B = 8'h26; #100;
A = 8'hBA; B = 8'h27; #100;
A = 8'hBA; B = 8'h28; #100;
A = 8'hBA; B = 8'h29; #100;
A = 8'hBA; B = 8'h2A; #100;
A = 8'hBA; B = 8'h2B; #100;
A = 8'hBA; B = 8'h2C; #100;
A = 8'hBA; B = 8'h2D; #100;
A = 8'hBA; B = 8'h2E; #100;
A = 8'hBA; B = 8'h2F; #100;
A = 8'hBA; B = 8'h30; #100;
A = 8'hBA; B = 8'h31; #100;
A = 8'hBA; B = 8'h32; #100;
A = 8'hBA; B = 8'h33; #100;
A = 8'hBA; B = 8'h34; #100;
A = 8'hBA; B = 8'h35; #100;
A = 8'hBA; B = 8'h36; #100;
A = 8'hBA; B = 8'h37; #100;
A = 8'hBA; B = 8'h38; #100;
A = 8'hBA; B = 8'h39; #100;
A = 8'hBA; B = 8'h3A; #100;
A = 8'hBA; B = 8'h3B; #100;
A = 8'hBA; B = 8'h3C; #100;
A = 8'hBA; B = 8'h3D; #100;
A = 8'hBA; B = 8'h3E; #100;
A = 8'hBA; B = 8'h3F; #100;
A = 8'hBA; B = 8'h40; #100;
A = 8'hBA; B = 8'h41; #100;
A = 8'hBA; B = 8'h42; #100;
A = 8'hBA; B = 8'h43; #100;
A = 8'hBA; B = 8'h44; #100;
A = 8'hBA; B = 8'h45; #100;
A = 8'hBA; B = 8'h46; #100;
A = 8'hBA; B = 8'h47; #100;
A = 8'hBA; B = 8'h48; #100;
A = 8'hBA; B = 8'h49; #100;
A = 8'hBA; B = 8'h4A; #100;
A = 8'hBA; B = 8'h4B; #100;
A = 8'hBA; B = 8'h4C; #100;
A = 8'hBA; B = 8'h4D; #100;
A = 8'hBA; B = 8'h4E; #100;
A = 8'hBA; B = 8'h4F; #100;
A = 8'hBA; B = 8'h50; #100;
A = 8'hBA; B = 8'h51; #100;
A = 8'hBA; B = 8'h52; #100;
A = 8'hBA; B = 8'h53; #100;
A = 8'hBA; B = 8'h54; #100;
A = 8'hBA; B = 8'h55; #100;
A = 8'hBA; B = 8'h56; #100;
A = 8'hBA; B = 8'h57; #100;
A = 8'hBA; B = 8'h58; #100;
A = 8'hBA; B = 8'h59; #100;
A = 8'hBA; B = 8'h5A; #100;
A = 8'hBA; B = 8'h5B; #100;
A = 8'hBA; B = 8'h5C; #100;
A = 8'hBA; B = 8'h5D; #100;
A = 8'hBA; B = 8'h5E; #100;
A = 8'hBA; B = 8'h5F; #100;
A = 8'hBA; B = 8'h60; #100;
A = 8'hBA; B = 8'h61; #100;
A = 8'hBA; B = 8'h62; #100;
A = 8'hBA; B = 8'h63; #100;
A = 8'hBA; B = 8'h64; #100;
A = 8'hBA; B = 8'h65; #100;
A = 8'hBA; B = 8'h66; #100;
A = 8'hBA; B = 8'h67; #100;
A = 8'hBA; B = 8'h68; #100;
A = 8'hBA; B = 8'h69; #100;
A = 8'hBA; B = 8'h6A; #100;
A = 8'hBA; B = 8'h6B; #100;
A = 8'hBA; B = 8'h6C; #100;
A = 8'hBA; B = 8'h6D; #100;
A = 8'hBA; B = 8'h6E; #100;
A = 8'hBA; B = 8'h6F; #100;
A = 8'hBA; B = 8'h70; #100;
A = 8'hBA; B = 8'h71; #100;
A = 8'hBA; B = 8'h72; #100;
A = 8'hBA; B = 8'h73; #100;
A = 8'hBA; B = 8'h74; #100;
A = 8'hBA; B = 8'h75; #100;
A = 8'hBA; B = 8'h76; #100;
A = 8'hBA; B = 8'h77; #100;
A = 8'hBA; B = 8'h78; #100;
A = 8'hBA; B = 8'h79; #100;
A = 8'hBA; B = 8'h7A; #100;
A = 8'hBA; B = 8'h7B; #100;
A = 8'hBA; B = 8'h7C; #100;
A = 8'hBA; B = 8'h7D; #100;
A = 8'hBA; B = 8'h7E; #100;
A = 8'hBA; B = 8'h7F; #100;
A = 8'hBA; B = 8'h80; #100;
A = 8'hBA; B = 8'h81; #100;
A = 8'hBA; B = 8'h82; #100;
A = 8'hBA; B = 8'h83; #100;
A = 8'hBA; B = 8'h84; #100;
A = 8'hBA; B = 8'h85; #100;
A = 8'hBA; B = 8'h86; #100;
A = 8'hBA; B = 8'h87; #100;
A = 8'hBA; B = 8'h88; #100;
A = 8'hBA; B = 8'h89; #100;
A = 8'hBA; B = 8'h8A; #100;
A = 8'hBA; B = 8'h8B; #100;
A = 8'hBA; B = 8'h8C; #100;
A = 8'hBA; B = 8'h8D; #100;
A = 8'hBA; B = 8'h8E; #100;
A = 8'hBA; B = 8'h8F; #100;
A = 8'hBA; B = 8'h90; #100;
A = 8'hBA; B = 8'h91; #100;
A = 8'hBA; B = 8'h92; #100;
A = 8'hBA; B = 8'h93; #100;
A = 8'hBA; B = 8'h94; #100;
A = 8'hBA; B = 8'h95; #100;
A = 8'hBA; B = 8'h96; #100;
A = 8'hBA; B = 8'h97; #100;
A = 8'hBA; B = 8'h98; #100;
A = 8'hBA; B = 8'h99; #100;
A = 8'hBA; B = 8'h9A; #100;
A = 8'hBA; B = 8'h9B; #100;
A = 8'hBA; B = 8'h9C; #100;
A = 8'hBA; B = 8'h9D; #100;
A = 8'hBA; B = 8'h9E; #100;
A = 8'hBA; B = 8'h9F; #100;
A = 8'hBA; B = 8'hA0; #100;
A = 8'hBA; B = 8'hA1; #100;
A = 8'hBA; B = 8'hA2; #100;
A = 8'hBA; B = 8'hA3; #100;
A = 8'hBA; B = 8'hA4; #100;
A = 8'hBA; B = 8'hA5; #100;
A = 8'hBA; B = 8'hA6; #100;
A = 8'hBA; B = 8'hA7; #100;
A = 8'hBA; B = 8'hA8; #100;
A = 8'hBA; B = 8'hA9; #100;
A = 8'hBA; B = 8'hAA; #100;
A = 8'hBA; B = 8'hAB; #100;
A = 8'hBA; B = 8'hAC; #100;
A = 8'hBA; B = 8'hAD; #100;
A = 8'hBA; B = 8'hAE; #100;
A = 8'hBA; B = 8'hAF; #100;
A = 8'hBA; B = 8'hB0; #100;
A = 8'hBA; B = 8'hB1; #100;
A = 8'hBA; B = 8'hB2; #100;
A = 8'hBA; B = 8'hB3; #100;
A = 8'hBA; B = 8'hB4; #100;
A = 8'hBA; B = 8'hB5; #100;
A = 8'hBA; B = 8'hB6; #100;
A = 8'hBA; B = 8'hB7; #100;
A = 8'hBA; B = 8'hB8; #100;
A = 8'hBA; B = 8'hB9; #100;
A = 8'hBA; B = 8'hBA; #100;
A = 8'hBA; B = 8'hBB; #100;
A = 8'hBA; B = 8'hBC; #100;
A = 8'hBA; B = 8'hBD; #100;
A = 8'hBA; B = 8'hBE; #100;
A = 8'hBA; B = 8'hBF; #100;
A = 8'hBA; B = 8'hC0; #100;
A = 8'hBA; B = 8'hC1; #100;
A = 8'hBA; B = 8'hC2; #100;
A = 8'hBA; B = 8'hC3; #100;
A = 8'hBA; B = 8'hC4; #100;
A = 8'hBA; B = 8'hC5; #100;
A = 8'hBA; B = 8'hC6; #100;
A = 8'hBA; B = 8'hC7; #100;
A = 8'hBA; B = 8'hC8; #100;
A = 8'hBA; B = 8'hC9; #100;
A = 8'hBA; B = 8'hCA; #100;
A = 8'hBA; B = 8'hCB; #100;
A = 8'hBA; B = 8'hCC; #100;
A = 8'hBA; B = 8'hCD; #100;
A = 8'hBA; B = 8'hCE; #100;
A = 8'hBA; B = 8'hCF; #100;
A = 8'hBA; B = 8'hD0; #100;
A = 8'hBA; B = 8'hD1; #100;
A = 8'hBA; B = 8'hD2; #100;
A = 8'hBA; B = 8'hD3; #100;
A = 8'hBA; B = 8'hD4; #100;
A = 8'hBA; B = 8'hD5; #100;
A = 8'hBA; B = 8'hD6; #100;
A = 8'hBA; B = 8'hD7; #100;
A = 8'hBA; B = 8'hD8; #100;
A = 8'hBA; B = 8'hD9; #100;
A = 8'hBA; B = 8'hDA; #100;
A = 8'hBA; B = 8'hDB; #100;
A = 8'hBA; B = 8'hDC; #100;
A = 8'hBA; B = 8'hDD; #100;
A = 8'hBA; B = 8'hDE; #100;
A = 8'hBA; B = 8'hDF; #100;
A = 8'hBA; B = 8'hE0; #100;
A = 8'hBA; B = 8'hE1; #100;
A = 8'hBA; B = 8'hE2; #100;
A = 8'hBA; B = 8'hE3; #100;
A = 8'hBA; B = 8'hE4; #100;
A = 8'hBA; B = 8'hE5; #100;
A = 8'hBA; B = 8'hE6; #100;
A = 8'hBA; B = 8'hE7; #100;
A = 8'hBA; B = 8'hE8; #100;
A = 8'hBA; B = 8'hE9; #100;
A = 8'hBA; B = 8'hEA; #100;
A = 8'hBA; B = 8'hEB; #100;
A = 8'hBA; B = 8'hEC; #100;
A = 8'hBA; B = 8'hED; #100;
A = 8'hBA; B = 8'hEE; #100;
A = 8'hBA; B = 8'hEF; #100;
A = 8'hBA; B = 8'hF0; #100;
A = 8'hBA; B = 8'hF1; #100;
A = 8'hBA; B = 8'hF2; #100;
A = 8'hBA; B = 8'hF3; #100;
A = 8'hBA; B = 8'hF4; #100;
A = 8'hBA; B = 8'hF5; #100;
A = 8'hBA; B = 8'hF6; #100;
A = 8'hBA; B = 8'hF7; #100;
A = 8'hBA; B = 8'hF8; #100;
A = 8'hBA; B = 8'hF9; #100;
A = 8'hBA; B = 8'hFA; #100;
A = 8'hBA; B = 8'hFB; #100;
A = 8'hBA; B = 8'hFC; #100;
A = 8'hBA; B = 8'hFD; #100;
A = 8'hBA; B = 8'hFE; #100;
A = 8'hBA; B = 8'hFF; #100;
A = 8'hBB; B = 8'h0; #100;
A = 8'hBB; B = 8'h1; #100;
A = 8'hBB; B = 8'h2; #100;
A = 8'hBB; B = 8'h3; #100;
A = 8'hBB; B = 8'h4; #100;
A = 8'hBB; B = 8'h5; #100;
A = 8'hBB; B = 8'h6; #100;
A = 8'hBB; B = 8'h7; #100;
A = 8'hBB; B = 8'h8; #100;
A = 8'hBB; B = 8'h9; #100;
A = 8'hBB; B = 8'hA; #100;
A = 8'hBB; B = 8'hB; #100;
A = 8'hBB; B = 8'hC; #100;
A = 8'hBB; B = 8'hD; #100;
A = 8'hBB; B = 8'hE; #100;
A = 8'hBB; B = 8'hF; #100;
A = 8'hBB; B = 8'h10; #100;
A = 8'hBB; B = 8'h11; #100;
A = 8'hBB; B = 8'h12; #100;
A = 8'hBB; B = 8'h13; #100;
A = 8'hBB; B = 8'h14; #100;
A = 8'hBB; B = 8'h15; #100;
A = 8'hBB; B = 8'h16; #100;
A = 8'hBB; B = 8'h17; #100;
A = 8'hBB; B = 8'h18; #100;
A = 8'hBB; B = 8'h19; #100;
A = 8'hBB; B = 8'h1A; #100;
A = 8'hBB; B = 8'h1B; #100;
A = 8'hBB; B = 8'h1C; #100;
A = 8'hBB; B = 8'h1D; #100;
A = 8'hBB; B = 8'h1E; #100;
A = 8'hBB; B = 8'h1F; #100;
A = 8'hBB; B = 8'h20; #100;
A = 8'hBB; B = 8'h21; #100;
A = 8'hBB; B = 8'h22; #100;
A = 8'hBB; B = 8'h23; #100;
A = 8'hBB; B = 8'h24; #100;
A = 8'hBB; B = 8'h25; #100;
A = 8'hBB; B = 8'h26; #100;
A = 8'hBB; B = 8'h27; #100;
A = 8'hBB; B = 8'h28; #100;
A = 8'hBB; B = 8'h29; #100;
A = 8'hBB; B = 8'h2A; #100;
A = 8'hBB; B = 8'h2B; #100;
A = 8'hBB; B = 8'h2C; #100;
A = 8'hBB; B = 8'h2D; #100;
A = 8'hBB; B = 8'h2E; #100;
A = 8'hBB; B = 8'h2F; #100;
A = 8'hBB; B = 8'h30; #100;
A = 8'hBB; B = 8'h31; #100;
A = 8'hBB; B = 8'h32; #100;
A = 8'hBB; B = 8'h33; #100;
A = 8'hBB; B = 8'h34; #100;
A = 8'hBB; B = 8'h35; #100;
A = 8'hBB; B = 8'h36; #100;
A = 8'hBB; B = 8'h37; #100;
A = 8'hBB; B = 8'h38; #100;
A = 8'hBB; B = 8'h39; #100;
A = 8'hBB; B = 8'h3A; #100;
A = 8'hBB; B = 8'h3B; #100;
A = 8'hBB; B = 8'h3C; #100;
A = 8'hBB; B = 8'h3D; #100;
A = 8'hBB; B = 8'h3E; #100;
A = 8'hBB; B = 8'h3F; #100;
A = 8'hBB; B = 8'h40; #100;
A = 8'hBB; B = 8'h41; #100;
A = 8'hBB; B = 8'h42; #100;
A = 8'hBB; B = 8'h43; #100;
A = 8'hBB; B = 8'h44; #100;
A = 8'hBB; B = 8'h45; #100;
A = 8'hBB; B = 8'h46; #100;
A = 8'hBB; B = 8'h47; #100;
A = 8'hBB; B = 8'h48; #100;
A = 8'hBB; B = 8'h49; #100;
A = 8'hBB; B = 8'h4A; #100;
A = 8'hBB; B = 8'h4B; #100;
A = 8'hBB; B = 8'h4C; #100;
A = 8'hBB; B = 8'h4D; #100;
A = 8'hBB; B = 8'h4E; #100;
A = 8'hBB; B = 8'h4F; #100;
A = 8'hBB; B = 8'h50; #100;
A = 8'hBB; B = 8'h51; #100;
A = 8'hBB; B = 8'h52; #100;
A = 8'hBB; B = 8'h53; #100;
A = 8'hBB; B = 8'h54; #100;
A = 8'hBB; B = 8'h55; #100;
A = 8'hBB; B = 8'h56; #100;
A = 8'hBB; B = 8'h57; #100;
A = 8'hBB; B = 8'h58; #100;
A = 8'hBB; B = 8'h59; #100;
A = 8'hBB; B = 8'h5A; #100;
A = 8'hBB; B = 8'h5B; #100;
A = 8'hBB; B = 8'h5C; #100;
A = 8'hBB; B = 8'h5D; #100;
A = 8'hBB; B = 8'h5E; #100;
A = 8'hBB; B = 8'h5F; #100;
A = 8'hBB; B = 8'h60; #100;
A = 8'hBB; B = 8'h61; #100;
A = 8'hBB; B = 8'h62; #100;
A = 8'hBB; B = 8'h63; #100;
A = 8'hBB; B = 8'h64; #100;
A = 8'hBB; B = 8'h65; #100;
A = 8'hBB; B = 8'h66; #100;
A = 8'hBB; B = 8'h67; #100;
A = 8'hBB; B = 8'h68; #100;
A = 8'hBB; B = 8'h69; #100;
A = 8'hBB; B = 8'h6A; #100;
A = 8'hBB; B = 8'h6B; #100;
A = 8'hBB; B = 8'h6C; #100;
A = 8'hBB; B = 8'h6D; #100;
A = 8'hBB; B = 8'h6E; #100;
A = 8'hBB; B = 8'h6F; #100;
A = 8'hBB; B = 8'h70; #100;
A = 8'hBB; B = 8'h71; #100;
A = 8'hBB; B = 8'h72; #100;
A = 8'hBB; B = 8'h73; #100;
A = 8'hBB; B = 8'h74; #100;
A = 8'hBB; B = 8'h75; #100;
A = 8'hBB; B = 8'h76; #100;
A = 8'hBB; B = 8'h77; #100;
A = 8'hBB; B = 8'h78; #100;
A = 8'hBB; B = 8'h79; #100;
A = 8'hBB; B = 8'h7A; #100;
A = 8'hBB; B = 8'h7B; #100;
A = 8'hBB; B = 8'h7C; #100;
A = 8'hBB; B = 8'h7D; #100;
A = 8'hBB; B = 8'h7E; #100;
A = 8'hBB; B = 8'h7F; #100;
A = 8'hBB; B = 8'h80; #100;
A = 8'hBB; B = 8'h81; #100;
A = 8'hBB; B = 8'h82; #100;
A = 8'hBB; B = 8'h83; #100;
A = 8'hBB; B = 8'h84; #100;
A = 8'hBB; B = 8'h85; #100;
A = 8'hBB; B = 8'h86; #100;
A = 8'hBB; B = 8'h87; #100;
A = 8'hBB; B = 8'h88; #100;
A = 8'hBB; B = 8'h89; #100;
A = 8'hBB; B = 8'h8A; #100;
A = 8'hBB; B = 8'h8B; #100;
A = 8'hBB; B = 8'h8C; #100;
A = 8'hBB; B = 8'h8D; #100;
A = 8'hBB; B = 8'h8E; #100;
A = 8'hBB; B = 8'h8F; #100;
A = 8'hBB; B = 8'h90; #100;
A = 8'hBB; B = 8'h91; #100;
A = 8'hBB; B = 8'h92; #100;
A = 8'hBB; B = 8'h93; #100;
A = 8'hBB; B = 8'h94; #100;
A = 8'hBB; B = 8'h95; #100;
A = 8'hBB; B = 8'h96; #100;
A = 8'hBB; B = 8'h97; #100;
A = 8'hBB; B = 8'h98; #100;
A = 8'hBB; B = 8'h99; #100;
A = 8'hBB; B = 8'h9A; #100;
A = 8'hBB; B = 8'h9B; #100;
A = 8'hBB; B = 8'h9C; #100;
A = 8'hBB; B = 8'h9D; #100;
A = 8'hBB; B = 8'h9E; #100;
A = 8'hBB; B = 8'h9F; #100;
A = 8'hBB; B = 8'hA0; #100;
A = 8'hBB; B = 8'hA1; #100;
A = 8'hBB; B = 8'hA2; #100;
A = 8'hBB; B = 8'hA3; #100;
A = 8'hBB; B = 8'hA4; #100;
A = 8'hBB; B = 8'hA5; #100;
A = 8'hBB; B = 8'hA6; #100;
A = 8'hBB; B = 8'hA7; #100;
A = 8'hBB; B = 8'hA8; #100;
A = 8'hBB; B = 8'hA9; #100;
A = 8'hBB; B = 8'hAA; #100;
A = 8'hBB; B = 8'hAB; #100;
A = 8'hBB; B = 8'hAC; #100;
A = 8'hBB; B = 8'hAD; #100;
A = 8'hBB; B = 8'hAE; #100;
A = 8'hBB; B = 8'hAF; #100;
A = 8'hBB; B = 8'hB0; #100;
A = 8'hBB; B = 8'hB1; #100;
A = 8'hBB; B = 8'hB2; #100;
A = 8'hBB; B = 8'hB3; #100;
A = 8'hBB; B = 8'hB4; #100;
A = 8'hBB; B = 8'hB5; #100;
A = 8'hBB; B = 8'hB6; #100;
A = 8'hBB; B = 8'hB7; #100;
A = 8'hBB; B = 8'hB8; #100;
A = 8'hBB; B = 8'hB9; #100;
A = 8'hBB; B = 8'hBA; #100;
A = 8'hBB; B = 8'hBB; #100;
A = 8'hBB; B = 8'hBC; #100;
A = 8'hBB; B = 8'hBD; #100;
A = 8'hBB; B = 8'hBE; #100;
A = 8'hBB; B = 8'hBF; #100;
A = 8'hBB; B = 8'hC0; #100;
A = 8'hBB; B = 8'hC1; #100;
A = 8'hBB; B = 8'hC2; #100;
A = 8'hBB; B = 8'hC3; #100;
A = 8'hBB; B = 8'hC4; #100;
A = 8'hBB; B = 8'hC5; #100;
A = 8'hBB; B = 8'hC6; #100;
A = 8'hBB; B = 8'hC7; #100;
A = 8'hBB; B = 8'hC8; #100;
A = 8'hBB; B = 8'hC9; #100;
A = 8'hBB; B = 8'hCA; #100;
A = 8'hBB; B = 8'hCB; #100;
A = 8'hBB; B = 8'hCC; #100;
A = 8'hBB; B = 8'hCD; #100;
A = 8'hBB; B = 8'hCE; #100;
A = 8'hBB; B = 8'hCF; #100;
A = 8'hBB; B = 8'hD0; #100;
A = 8'hBB; B = 8'hD1; #100;
A = 8'hBB; B = 8'hD2; #100;
A = 8'hBB; B = 8'hD3; #100;
A = 8'hBB; B = 8'hD4; #100;
A = 8'hBB; B = 8'hD5; #100;
A = 8'hBB; B = 8'hD6; #100;
A = 8'hBB; B = 8'hD7; #100;
A = 8'hBB; B = 8'hD8; #100;
A = 8'hBB; B = 8'hD9; #100;
A = 8'hBB; B = 8'hDA; #100;
A = 8'hBB; B = 8'hDB; #100;
A = 8'hBB; B = 8'hDC; #100;
A = 8'hBB; B = 8'hDD; #100;
A = 8'hBB; B = 8'hDE; #100;
A = 8'hBB; B = 8'hDF; #100;
A = 8'hBB; B = 8'hE0; #100;
A = 8'hBB; B = 8'hE1; #100;
A = 8'hBB; B = 8'hE2; #100;
A = 8'hBB; B = 8'hE3; #100;
A = 8'hBB; B = 8'hE4; #100;
A = 8'hBB; B = 8'hE5; #100;
A = 8'hBB; B = 8'hE6; #100;
A = 8'hBB; B = 8'hE7; #100;
A = 8'hBB; B = 8'hE8; #100;
A = 8'hBB; B = 8'hE9; #100;
A = 8'hBB; B = 8'hEA; #100;
A = 8'hBB; B = 8'hEB; #100;
A = 8'hBB; B = 8'hEC; #100;
A = 8'hBB; B = 8'hED; #100;
A = 8'hBB; B = 8'hEE; #100;
A = 8'hBB; B = 8'hEF; #100;
A = 8'hBB; B = 8'hF0; #100;
A = 8'hBB; B = 8'hF1; #100;
A = 8'hBB; B = 8'hF2; #100;
A = 8'hBB; B = 8'hF3; #100;
A = 8'hBB; B = 8'hF4; #100;
A = 8'hBB; B = 8'hF5; #100;
A = 8'hBB; B = 8'hF6; #100;
A = 8'hBB; B = 8'hF7; #100;
A = 8'hBB; B = 8'hF8; #100;
A = 8'hBB; B = 8'hF9; #100;
A = 8'hBB; B = 8'hFA; #100;
A = 8'hBB; B = 8'hFB; #100;
A = 8'hBB; B = 8'hFC; #100;
A = 8'hBB; B = 8'hFD; #100;
A = 8'hBB; B = 8'hFE; #100;
A = 8'hBB; B = 8'hFF; #100;
A = 8'hBC; B = 8'h0; #100;
A = 8'hBC; B = 8'h1; #100;
A = 8'hBC; B = 8'h2; #100;
A = 8'hBC; B = 8'h3; #100;
A = 8'hBC; B = 8'h4; #100;
A = 8'hBC; B = 8'h5; #100;
A = 8'hBC; B = 8'h6; #100;
A = 8'hBC; B = 8'h7; #100;
A = 8'hBC; B = 8'h8; #100;
A = 8'hBC; B = 8'h9; #100;
A = 8'hBC; B = 8'hA; #100;
A = 8'hBC; B = 8'hB; #100;
A = 8'hBC; B = 8'hC; #100;
A = 8'hBC; B = 8'hD; #100;
A = 8'hBC; B = 8'hE; #100;
A = 8'hBC; B = 8'hF; #100;
A = 8'hBC; B = 8'h10; #100;
A = 8'hBC; B = 8'h11; #100;
A = 8'hBC; B = 8'h12; #100;
A = 8'hBC; B = 8'h13; #100;
A = 8'hBC; B = 8'h14; #100;
A = 8'hBC; B = 8'h15; #100;
A = 8'hBC; B = 8'h16; #100;
A = 8'hBC; B = 8'h17; #100;
A = 8'hBC; B = 8'h18; #100;
A = 8'hBC; B = 8'h19; #100;
A = 8'hBC; B = 8'h1A; #100;
A = 8'hBC; B = 8'h1B; #100;
A = 8'hBC; B = 8'h1C; #100;
A = 8'hBC; B = 8'h1D; #100;
A = 8'hBC; B = 8'h1E; #100;
A = 8'hBC; B = 8'h1F; #100;
A = 8'hBC; B = 8'h20; #100;
A = 8'hBC; B = 8'h21; #100;
A = 8'hBC; B = 8'h22; #100;
A = 8'hBC; B = 8'h23; #100;
A = 8'hBC; B = 8'h24; #100;
A = 8'hBC; B = 8'h25; #100;
A = 8'hBC; B = 8'h26; #100;
A = 8'hBC; B = 8'h27; #100;
A = 8'hBC; B = 8'h28; #100;
A = 8'hBC; B = 8'h29; #100;
A = 8'hBC; B = 8'h2A; #100;
A = 8'hBC; B = 8'h2B; #100;
A = 8'hBC; B = 8'h2C; #100;
A = 8'hBC; B = 8'h2D; #100;
A = 8'hBC; B = 8'h2E; #100;
A = 8'hBC; B = 8'h2F; #100;
A = 8'hBC; B = 8'h30; #100;
A = 8'hBC; B = 8'h31; #100;
A = 8'hBC; B = 8'h32; #100;
A = 8'hBC; B = 8'h33; #100;
A = 8'hBC; B = 8'h34; #100;
A = 8'hBC; B = 8'h35; #100;
A = 8'hBC; B = 8'h36; #100;
A = 8'hBC; B = 8'h37; #100;
A = 8'hBC; B = 8'h38; #100;
A = 8'hBC; B = 8'h39; #100;
A = 8'hBC; B = 8'h3A; #100;
A = 8'hBC; B = 8'h3B; #100;
A = 8'hBC; B = 8'h3C; #100;
A = 8'hBC; B = 8'h3D; #100;
A = 8'hBC; B = 8'h3E; #100;
A = 8'hBC; B = 8'h3F; #100;
A = 8'hBC; B = 8'h40; #100;
A = 8'hBC; B = 8'h41; #100;
A = 8'hBC; B = 8'h42; #100;
A = 8'hBC; B = 8'h43; #100;
A = 8'hBC; B = 8'h44; #100;
A = 8'hBC; B = 8'h45; #100;
A = 8'hBC; B = 8'h46; #100;
A = 8'hBC; B = 8'h47; #100;
A = 8'hBC; B = 8'h48; #100;
A = 8'hBC; B = 8'h49; #100;
A = 8'hBC; B = 8'h4A; #100;
A = 8'hBC; B = 8'h4B; #100;
A = 8'hBC; B = 8'h4C; #100;
A = 8'hBC; B = 8'h4D; #100;
A = 8'hBC; B = 8'h4E; #100;
A = 8'hBC; B = 8'h4F; #100;
A = 8'hBC; B = 8'h50; #100;
A = 8'hBC; B = 8'h51; #100;
A = 8'hBC; B = 8'h52; #100;
A = 8'hBC; B = 8'h53; #100;
A = 8'hBC; B = 8'h54; #100;
A = 8'hBC; B = 8'h55; #100;
A = 8'hBC; B = 8'h56; #100;
A = 8'hBC; B = 8'h57; #100;
A = 8'hBC; B = 8'h58; #100;
A = 8'hBC; B = 8'h59; #100;
A = 8'hBC; B = 8'h5A; #100;
A = 8'hBC; B = 8'h5B; #100;
A = 8'hBC; B = 8'h5C; #100;
A = 8'hBC; B = 8'h5D; #100;
A = 8'hBC; B = 8'h5E; #100;
A = 8'hBC; B = 8'h5F; #100;
A = 8'hBC; B = 8'h60; #100;
A = 8'hBC; B = 8'h61; #100;
A = 8'hBC; B = 8'h62; #100;
A = 8'hBC; B = 8'h63; #100;
A = 8'hBC; B = 8'h64; #100;
A = 8'hBC; B = 8'h65; #100;
A = 8'hBC; B = 8'h66; #100;
A = 8'hBC; B = 8'h67; #100;
A = 8'hBC; B = 8'h68; #100;
A = 8'hBC; B = 8'h69; #100;
A = 8'hBC; B = 8'h6A; #100;
A = 8'hBC; B = 8'h6B; #100;
A = 8'hBC; B = 8'h6C; #100;
A = 8'hBC; B = 8'h6D; #100;
A = 8'hBC; B = 8'h6E; #100;
A = 8'hBC; B = 8'h6F; #100;
A = 8'hBC; B = 8'h70; #100;
A = 8'hBC; B = 8'h71; #100;
A = 8'hBC; B = 8'h72; #100;
A = 8'hBC; B = 8'h73; #100;
A = 8'hBC; B = 8'h74; #100;
A = 8'hBC; B = 8'h75; #100;
A = 8'hBC; B = 8'h76; #100;
A = 8'hBC; B = 8'h77; #100;
A = 8'hBC; B = 8'h78; #100;
A = 8'hBC; B = 8'h79; #100;
A = 8'hBC; B = 8'h7A; #100;
A = 8'hBC; B = 8'h7B; #100;
A = 8'hBC; B = 8'h7C; #100;
A = 8'hBC; B = 8'h7D; #100;
A = 8'hBC; B = 8'h7E; #100;
A = 8'hBC; B = 8'h7F; #100;
A = 8'hBC; B = 8'h80; #100;
A = 8'hBC; B = 8'h81; #100;
A = 8'hBC; B = 8'h82; #100;
A = 8'hBC; B = 8'h83; #100;
A = 8'hBC; B = 8'h84; #100;
A = 8'hBC; B = 8'h85; #100;
A = 8'hBC; B = 8'h86; #100;
A = 8'hBC; B = 8'h87; #100;
A = 8'hBC; B = 8'h88; #100;
A = 8'hBC; B = 8'h89; #100;
A = 8'hBC; B = 8'h8A; #100;
A = 8'hBC; B = 8'h8B; #100;
A = 8'hBC; B = 8'h8C; #100;
A = 8'hBC; B = 8'h8D; #100;
A = 8'hBC; B = 8'h8E; #100;
A = 8'hBC; B = 8'h8F; #100;
A = 8'hBC; B = 8'h90; #100;
A = 8'hBC; B = 8'h91; #100;
A = 8'hBC; B = 8'h92; #100;
A = 8'hBC; B = 8'h93; #100;
A = 8'hBC; B = 8'h94; #100;
A = 8'hBC; B = 8'h95; #100;
A = 8'hBC; B = 8'h96; #100;
A = 8'hBC; B = 8'h97; #100;
A = 8'hBC; B = 8'h98; #100;
A = 8'hBC; B = 8'h99; #100;
A = 8'hBC; B = 8'h9A; #100;
A = 8'hBC; B = 8'h9B; #100;
A = 8'hBC; B = 8'h9C; #100;
A = 8'hBC; B = 8'h9D; #100;
A = 8'hBC; B = 8'h9E; #100;
A = 8'hBC; B = 8'h9F; #100;
A = 8'hBC; B = 8'hA0; #100;
A = 8'hBC; B = 8'hA1; #100;
A = 8'hBC; B = 8'hA2; #100;
A = 8'hBC; B = 8'hA3; #100;
A = 8'hBC; B = 8'hA4; #100;
A = 8'hBC; B = 8'hA5; #100;
A = 8'hBC; B = 8'hA6; #100;
A = 8'hBC; B = 8'hA7; #100;
A = 8'hBC; B = 8'hA8; #100;
A = 8'hBC; B = 8'hA9; #100;
A = 8'hBC; B = 8'hAA; #100;
A = 8'hBC; B = 8'hAB; #100;
A = 8'hBC; B = 8'hAC; #100;
A = 8'hBC; B = 8'hAD; #100;
A = 8'hBC; B = 8'hAE; #100;
A = 8'hBC; B = 8'hAF; #100;
A = 8'hBC; B = 8'hB0; #100;
A = 8'hBC; B = 8'hB1; #100;
A = 8'hBC; B = 8'hB2; #100;
A = 8'hBC; B = 8'hB3; #100;
A = 8'hBC; B = 8'hB4; #100;
A = 8'hBC; B = 8'hB5; #100;
A = 8'hBC; B = 8'hB6; #100;
A = 8'hBC; B = 8'hB7; #100;
A = 8'hBC; B = 8'hB8; #100;
A = 8'hBC; B = 8'hB9; #100;
A = 8'hBC; B = 8'hBA; #100;
A = 8'hBC; B = 8'hBB; #100;
A = 8'hBC; B = 8'hBC; #100;
A = 8'hBC; B = 8'hBD; #100;
A = 8'hBC; B = 8'hBE; #100;
A = 8'hBC; B = 8'hBF; #100;
A = 8'hBC; B = 8'hC0; #100;
A = 8'hBC; B = 8'hC1; #100;
A = 8'hBC; B = 8'hC2; #100;
A = 8'hBC; B = 8'hC3; #100;
A = 8'hBC; B = 8'hC4; #100;
A = 8'hBC; B = 8'hC5; #100;
A = 8'hBC; B = 8'hC6; #100;
A = 8'hBC; B = 8'hC7; #100;
A = 8'hBC; B = 8'hC8; #100;
A = 8'hBC; B = 8'hC9; #100;
A = 8'hBC; B = 8'hCA; #100;
A = 8'hBC; B = 8'hCB; #100;
A = 8'hBC; B = 8'hCC; #100;
A = 8'hBC; B = 8'hCD; #100;
A = 8'hBC; B = 8'hCE; #100;
A = 8'hBC; B = 8'hCF; #100;
A = 8'hBC; B = 8'hD0; #100;
A = 8'hBC; B = 8'hD1; #100;
A = 8'hBC; B = 8'hD2; #100;
A = 8'hBC; B = 8'hD3; #100;
A = 8'hBC; B = 8'hD4; #100;
A = 8'hBC; B = 8'hD5; #100;
A = 8'hBC; B = 8'hD6; #100;
A = 8'hBC; B = 8'hD7; #100;
A = 8'hBC; B = 8'hD8; #100;
A = 8'hBC; B = 8'hD9; #100;
A = 8'hBC; B = 8'hDA; #100;
A = 8'hBC; B = 8'hDB; #100;
A = 8'hBC; B = 8'hDC; #100;
A = 8'hBC; B = 8'hDD; #100;
A = 8'hBC; B = 8'hDE; #100;
A = 8'hBC; B = 8'hDF; #100;
A = 8'hBC; B = 8'hE0; #100;
A = 8'hBC; B = 8'hE1; #100;
A = 8'hBC; B = 8'hE2; #100;
A = 8'hBC; B = 8'hE3; #100;
A = 8'hBC; B = 8'hE4; #100;
A = 8'hBC; B = 8'hE5; #100;
A = 8'hBC; B = 8'hE6; #100;
A = 8'hBC; B = 8'hE7; #100;
A = 8'hBC; B = 8'hE8; #100;
A = 8'hBC; B = 8'hE9; #100;
A = 8'hBC; B = 8'hEA; #100;
A = 8'hBC; B = 8'hEB; #100;
A = 8'hBC; B = 8'hEC; #100;
A = 8'hBC; B = 8'hED; #100;
A = 8'hBC; B = 8'hEE; #100;
A = 8'hBC; B = 8'hEF; #100;
A = 8'hBC; B = 8'hF0; #100;
A = 8'hBC; B = 8'hF1; #100;
A = 8'hBC; B = 8'hF2; #100;
A = 8'hBC; B = 8'hF3; #100;
A = 8'hBC; B = 8'hF4; #100;
A = 8'hBC; B = 8'hF5; #100;
A = 8'hBC; B = 8'hF6; #100;
A = 8'hBC; B = 8'hF7; #100;
A = 8'hBC; B = 8'hF8; #100;
A = 8'hBC; B = 8'hF9; #100;
A = 8'hBC; B = 8'hFA; #100;
A = 8'hBC; B = 8'hFB; #100;
A = 8'hBC; B = 8'hFC; #100;
A = 8'hBC; B = 8'hFD; #100;
A = 8'hBC; B = 8'hFE; #100;
A = 8'hBC; B = 8'hFF; #100;
A = 8'hBD; B = 8'h0; #100;
A = 8'hBD; B = 8'h1; #100;
A = 8'hBD; B = 8'h2; #100;
A = 8'hBD; B = 8'h3; #100;
A = 8'hBD; B = 8'h4; #100;
A = 8'hBD; B = 8'h5; #100;
A = 8'hBD; B = 8'h6; #100;
A = 8'hBD; B = 8'h7; #100;
A = 8'hBD; B = 8'h8; #100;
A = 8'hBD; B = 8'h9; #100;
A = 8'hBD; B = 8'hA; #100;
A = 8'hBD; B = 8'hB; #100;
A = 8'hBD; B = 8'hC; #100;
A = 8'hBD; B = 8'hD; #100;
A = 8'hBD; B = 8'hE; #100;
A = 8'hBD; B = 8'hF; #100;
A = 8'hBD; B = 8'h10; #100;
A = 8'hBD; B = 8'h11; #100;
A = 8'hBD; B = 8'h12; #100;
A = 8'hBD; B = 8'h13; #100;
A = 8'hBD; B = 8'h14; #100;
A = 8'hBD; B = 8'h15; #100;
A = 8'hBD; B = 8'h16; #100;
A = 8'hBD; B = 8'h17; #100;
A = 8'hBD; B = 8'h18; #100;
A = 8'hBD; B = 8'h19; #100;
A = 8'hBD; B = 8'h1A; #100;
A = 8'hBD; B = 8'h1B; #100;
A = 8'hBD; B = 8'h1C; #100;
A = 8'hBD; B = 8'h1D; #100;
A = 8'hBD; B = 8'h1E; #100;
A = 8'hBD; B = 8'h1F; #100;
A = 8'hBD; B = 8'h20; #100;
A = 8'hBD; B = 8'h21; #100;
A = 8'hBD; B = 8'h22; #100;
A = 8'hBD; B = 8'h23; #100;
A = 8'hBD; B = 8'h24; #100;
A = 8'hBD; B = 8'h25; #100;
A = 8'hBD; B = 8'h26; #100;
A = 8'hBD; B = 8'h27; #100;
A = 8'hBD; B = 8'h28; #100;
A = 8'hBD; B = 8'h29; #100;
A = 8'hBD; B = 8'h2A; #100;
A = 8'hBD; B = 8'h2B; #100;
A = 8'hBD; B = 8'h2C; #100;
A = 8'hBD; B = 8'h2D; #100;
A = 8'hBD; B = 8'h2E; #100;
A = 8'hBD; B = 8'h2F; #100;
A = 8'hBD; B = 8'h30; #100;
A = 8'hBD; B = 8'h31; #100;
A = 8'hBD; B = 8'h32; #100;
A = 8'hBD; B = 8'h33; #100;
A = 8'hBD; B = 8'h34; #100;
A = 8'hBD; B = 8'h35; #100;
A = 8'hBD; B = 8'h36; #100;
A = 8'hBD; B = 8'h37; #100;
A = 8'hBD; B = 8'h38; #100;
A = 8'hBD; B = 8'h39; #100;
A = 8'hBD; B = 8'h3A; #100;
A = 8'hBD; B = 8'h3B; #100;
A = 8'hBD; B = 8'h3C; #100;
A = 8'hBD; B = 8'h3D; #100;
A = 8'hBD; B = 8'h3E; #100;
A = 8'hBD; B = 8'h3F; #100;
A = 8'hBD; B = 8'h40; #100;
A = 8'hBD; B = 8'h41; #100;
A = 8'hBD; B = 8'h42; #100;
A = 8'hBD; B = 8'h43; #100;
A = 8'hBD; B = 8'h44; #100;
A = 8'hBD; B = 8'h45; #100;
A = 8'hBD; B = 8'h46; #100;
A = 8'hBD; B = 8'h47; #100;
A = 8'hBD; B = 8'h48; #100;
A = 8'hBD; B = 8'h49; #100;
A = 8'hBD; B = 8'h4A; #100;
A = 8'hBD; B = 8'h4B; #100;
A = 8'hBD; B = 8'h4C; #100;
A = 8'hBD; B = 8'h4D; #100;
A = 8'hBD; B = 8'h4E; #100;
A = 8'hBD; B = 8'h4F; #100;
A = 8'hBD; B = 8'h50; #100;
A = 8'hBD; B = 8'h51; #100;
A = 8'hBD; B = 8'h52; #100;
A = 8'hBD; B = 8'h53; #100;
A = 8'hBD; B = 8'h54; #100;
A = 8'hBD; B = 8'h55; #100;
A = 8'hBD; B = 8'h56; #100;
A = 8'hBD; B = 8'h57; #100;
A = 8'hBD; B = 8'h58; #100;
A = 8'hBD; B = 8'h59; #100;
A = 8'hBD; B = 8'h5A; #100;
A = 8'hBD; B = 8'h5B; #100;
A = 8'hBD; B = 8'h5C; #100;
A = 8'hBD; B = 8'h5D; #100;
A = 8'hBD; B = 8'h5E; #100;
A = 8'hBD; B = 8'h5F; #100;
A = 8'hBD; B = 8'h60; #100;
A = 8'hBD; B = 8'h61; #100;
A = 8'hBD; B = 8'h62; #100;
A = 8'hBD; B = 8'h63; #100;
A = 8'hBD; B = 8'h64; #100;
A = 8'hBD; B = 8'h65; #100;
A = 8'hBD; B = 8'h66; #100;
A = 8'hBD; B = 8'h67; #100;
A = 8'hBD; B = 8'h68; #100;
A = 8'hBD; B = 8'h69; #100;
A = 8'hBD; B = 8'h6A; #100;
A = 8'hBD; B = 8'h6B; #100;
A = 8'hBD; B = 8'h6C; #100;
A = 8'hBD; B = 8'h6D; #100;
A = 8'hBD; B = 8'h6E; #100;
A = 8'hBD; B = 8'h6F; #100;
A = 8'hBD; B = 8'h70; #100;
A = 8'hBD; B = 8'h71; #100;
A = 8'hBD; B = 8'h72; #100;
A = 8'hBD; B = 8'h73; #100;
A = 8'hBD; B = 8'h74; #100;
A = 8'hBD; B = 8'h75; #100;
A = 8'hBD; B = 8'h76; #100;
A = 8'hBD; B = 8'h77; #100;
A = 8'hBD; B = 8'h78; #100;
A = 8'hBD; B = 8'h79; #100;
A = 8'hBD; B = 8'h7A; #100;
A = 8'hBD; B = 8'h7B; #100;
A = 8'hBD; B = 8'h7C; #100;
A = 8'hBD; B = 8'h7D; #100;
A = 8'hBD; B = 8'h7E; #100;
A = 8'hBD; B = 8'h7F; #100;
A = 8'hBD; B = 8'h80; #100;
A = 8'hBD; B = 8'h81; #100;
A = 8'hBD; B = 8'h82; #100;
A = 8'hBD; B = 8'h83; #100;
A = 8'hBD; B = 8'h84; #100;
A = 8'hBD; B = 8'h85; #100;
A = 8'hBD; B = 8'h86; #100;
A = 8'hBD; B = 8'h87; #100;
A = 8'hBD; B = 8'h88; #100;
A = 8'hBD; B = 8'h89; #100;
A = 8'hBD; B = 8'h8A; #100;
A = 8'hBD; B = 8'h8B; #100;
A = 8'hBD; B = 8'h8C; #100;
A = 8'hBD; B = 8'h8D; #100;
A = 8'hBD; B = 8'h8E; #100;
A = 8'hBD; B = 8'h8F; #100;
A = 8'hBD; B = 8'h90; #100;
A = 8'hBD; B = 8'h91; #100;
A = 8'hBD; B = 8'h92; #100;
A = 8'hBD; B = 8'h93; #100;
A = 8'hBD; B = 8'h94; #100;
A = 8'hBD; B = 8'h95; #100;
A = 8'hBD; B = 8'h96; #100;
A = 8'hBD; B = 8'h97; #100;
A = 8'hBD; B = 8'h98; #100;
A = 8'hBD; B = 8'h99; #100;
A = 8'hBD; B = 8'h9A; #100;
A = 8'hBD; B = 8'h9B; #100;
A = 8'hBD; B = 8'h9C; #100;
A = 8'hBD; B = 8'h9D; #100;
A = 8'hBD; B = 8'h9E; #100;
A = 8'hBD; B = 8'h9F; #100;
A = 8'hBD; B = 8'hA0; #100;
A = 8'hBD; B = 8'hA1; #100;
A = 8'hBD; B = 8'hA2; #100;
A = 8'hBD; B = 8'hA3; #100;
A = 8'hBD; B = 8'hA4; #100;
A = 8'hBD; B = 8'hA5; #100;
A = 8'hBD; B = 8'hA6; #100;
A = 8'hBD; B = 8'hA7; #100;
A = 8'hBD; B = 8'hA8; #100;
A = 8'hBD; B = 8'hA9; #100;
A = 8'hBD; B = 8'hAA; #100;
A = 8'hBD; B = 8'hAB; #100;
A = 8'hBD; B = 8'hAC; #100;
A = 8'hBD; B = 8'hAD; #100;
A = 8'hBD; B = 8'hAE; #100;
A = 8'hBD; B = 8'hAF; #100;
A = 8'hBD; B = 8'hB0; #100;
A = 8'hBD; B = 8'hB1; #100;
A = 8'hBD; B = 8'hB2; #100;
A = 8'hBD; B = 8'hB3; #100;
A = 8'hBD; B = 8'hB4; #100;
A = 8'hBD; B = 8'hB5; #100;
A = 8'hBD; B = 8'hB6; #100;
A = 8'hBD; B = 8'hB7; #100;
A = 8'hBD; B = 8'hB8; #100;
A = 8'hBD; B = 8'hB9; #100;
A = 8'hBD; B = 8'hBA; #100;
A = 8'hBD; B = 8'hBB; #100;
A = 8'hBD; B = 8'hBC; #100;
A = 8'hBD; B = 8'hBD; #100;
A = 8'hBD; B = 8'hBE; #100;
A = 8'hBD; B = 8'hBF; #100;
A = 8'hBD; B = 8'hC0; #100;
A = 8'hBD; B = 8'hC1; #100;
A = 8'hBD; B = 8'hC2; #100;
A = 8'hBD; B = 8'hC3; #100;
A = 8'hBD; B = 8'hC4; #100;
A = 8'hBD; B = 8'hC5; #100;
A = 8'hBD; B = 8'hC6; #100;
A = 8'hBD; B = 8'hC7; #100;
A = 8'hBD; B = 8'hC8; #100;
A = 8'hBD; B = 8'hC9; #100;
A = 8'hBD; B = 8'hCA; #100;
A = 8'hBD; B = 8'hCB; #100;
A = 8'hBD; B = 8'hCC; #100;
A = 8'hBD; B = 8'hCD; #100;
A = 8'hBD; B = 8'hCE; #100;
A = 8'hBD; B = 8'hCF; #100;
A = 8'hBD; B = 8'hD0; #100;
A = 8'hBD; B = 8'hD1; #100;
A = 8'hBD; B = 8'hD2; #100;
A = 8'hBD; B = 8'hD3; #100;
A = 8'hBD; B = 8'hD4; #100;
A = 8'hBD; B = 8'hD5; #100;
A = 8'hBD; B = 8'hD6; #100;
A = 8'hBD; B = 8'hD7; #100;
A = 8'hBD; B = 8'hD8; #100;
A = 8'hBD; B = 8'hD9; #100;
A = 8'hBD; B = 8'hDA; #100;
A = 8'hBD; B = 8'hDB; #100;
A = 8'hBD; B = 8'hDC; #100;
A = 8'hBD; B = 8'hDD; #100;
A = 8'hBD; B = 8'hDE; #100;
A = 8'hBD; B = 8'hDF; #100;
A = 8'hBD; B = 8'hE0; #100;
A = 8'hBD; B = 8'hE1; #100;
A = 8'hBD; B = 8'hE2; #100;
A = 8'hBD; B = 8'hE3; #100;
A = 8'hBD; B = 8'hE4; #100;
A = 8'hBD; B = 8'hE5; #100;
A = 8'hBD; B = 8'hE6; #100;
A = 8'hBD; B = 8'hE7; #100;
A = 8'hBD; B = 8'hE8; #100;
A = 8'hBD; B = 8'hE9; #100;
A = 8'hBD; B = 8'hEA; #100;
A = 8'hBD; B = 8'hEB; #100;
A = 8'hBD; B = 8'hEC; #100;
A = 8'hBD; B = 8'hED; #100;
A = 8'hBD; B = 8'hEE; #100;
A = 8'hBD; B = 8'hEF; #100;
A = 8'hBD; B = 8'hF0; #100;
A = 8'hBD; B = 8'hF1; #100;
A = 8'hBD; B = 8'hF2; #100;
A = 8'hBD; B = 8'hF3; #100;
A = 8'hBD; B = 8'hF4; #100;
A = 8'hBD; B = 8'hF5; #100;
A = 8'hBD; B = 8'hF6; #100;
A = 8'hBD; B = 8'hF7; #100;
A = 8'hBD; B = 8'hF8; #100;
A = 8'hBD; B = 8'hF9; #100;
A = 8'hBD; B = 8'hFA; #100;
A = 8'hBD; B = 8'hFB; #100;
A = 8'hBD; B = 8'hFC; #100;
A = 8'hBD; B = 8'hFD; #100;
A = 8'hBD; B = 8'hFE; #100;
A = 8'hBD; B = 8'hFF; #100;
A = 8'hBE; B = 8'h0; #100;
A = 8'hBE; B = 8'h1; #100;
A = 8'hBE; B = 8'h2; #100;
A = 8'hBE; B = 8'h3; #100;
A = 8'hBE; B = 8'h4; #100;
A = 8'hBE; B = 8'h5; #100;
A = 8'hBE; B = 8'h6; #100;
A = 8'hBE; B = 8'h7; #100;
A = 8'hBE; B = 8'h8; #100;
A = 8'hBE; B = 8'h9; #100;
A = 8'hBE; B = 8'hA; #100;
A = 8'hBE; B = 8'hB; #100;
A = 8'hBE; B = 8'hC; #100;
A = 8'hBE; B = 8'hD; #100;
A = 8'hBE; B = 8'hE; #100;
A = 8'hBE; B = 8'hF; #100;
A = 8'hBE; B = 8'h10; #100;
A = 8'hBE; B = 8'h11; #100;
A = 8'hBE; B = 8'h12; #100;
A = 8'hBE; B = 8'h13; #100;
A = 8'hBE; B = 8'h14; #100;
A = 8'hBE; B = 8'h15; #100;
A = 8'hBE; B = 8'h16; #100;
A = 8'hBE; B = 8'h17; #100;
A = 8'hBE; B = 8'h18; #100;
A = 8'hBE; B = 8'h19; #100;
A = 8'hBE; B = 8'h1A; #100;
A = 8'hBE; B = 8'h1B; #100;
A = 8'hBE; B = 8'h1C; #100;
A = 8'hBE; B = 8'h1D; #100;
A = 8'hBE; B = 8'h1E; #100;
A = 8'hBE; B = 8'h1F; #100;
A = 8'hBE; B = 8'h20; #100;
A = 8'hBE; B = 8'h21; #100;
A = 8'hBE; B = 8'h22; #100;
A = 8'hBE; B = 8'h23; #100;
A = 8'hBE; B = 8'h24; #100;
A = 8'hBE; B = 8'h25; #100;
A = 8'hBE; B = 8'h26; #100;
A = 8'hBE; B = 8'h27; #100;
A = 8'hBE; B = 8'h28; #100;
A = 8'hBE; B = 8'h29; #100;
A = 8'hBE; B = 8'h2A; #100;
A = 8'hBE; B = 8'h2B; #100;
A = 8'hBE; B = 8'h2C; #100;
A = 8'hBE; B = 8'h2D; #100;
A = 8'hBE; B = 8'h2E; #100;
A = 8'hBE; B = 8'h2F; #100;
A = 8'hBE; B = 8'h30; #100;
A = 8'hBE; B = 8'h31; #100;
A = 8'hBE; B = 8'h32; #100;
A = 8'hBE; B = 8'h33; #100;
A = 8'hBE; B = 8'h34; #100;
A = 8'hBE; B = 8'h35; #100;
A = 8'hBE; B = 8'h36; #100;
A = 8'hBE; B = 8'h37; #100;
A = 8'hBE; B = 8'h38; #100;
A = 8'hBE; B = 8'h39; #100;
A = 8'hBE; B = 8'h3A; #100;
A = 8'hBE; B = 8'h3B; #100;
A = 8'hBE; B = 8'h3C; #100;
A = 8'hBE; B = 8'h3D; #100;
A = 8'hBE; B = 8'h3E; #100;
A = 8'hBE; B = 8'h3F; #100;
A = 8'hBE; B = 8'h40; #100;
A = 8'hBE; B = 8'h41; #100;
A = 8'hBE; B = 8'h42; #100;
A = 8'hBE; B = 8'h43; #100;
A = 8'hBE; B = 8'h44; #100;
A = 8'hBE; B = 8'h45; #100;
A = 8'hBE; B = 8'h46; #100;
A = 8'hBE; B = 8'h47; #100;
A = 8'hBE; B = 8'h48; #100;
A = 8'hBE; B = 8'h49; #100;
A = 8'hBE; B = 8'h4A; #100;
A = 8'hBE; B = 8'h4B; #100;
A = 8'hBE; B = 8'h4C; #100;
A = 8'hBE; B = 8'h4D; #100;
A = 8'hBE; B = 8'h4E; #100;
A = 8'hBE; B = 8'h4F; #100;
A = 8'hBE; B = 8'h50; #100;
A = 8'hBE; B = 8'h51; #100;
A = 8'hBE; B = 8'h52; #100;
A = 8'hBE; B = 8'h53; #100;
A = 8'hBE; B = 8'h54; #100;
A = 8'hBE; B = 8'h55; #100;
A = 8'hBE; B = 8'h56; #100;
A = 8'hBE; B = 8'h57; #100;
A = 8'hBE; B = 8'h58; #100;
A = 8'hBE; B = 8'h59; #100;
A = 8'hBE; B = 8'h5A; #100;
A = 8'hBE; B = 8'h5B; #100;
A = 8'hBE; B = 8'h5C; #100;
A = 8'hBE; B = 8'h5D; #100;
A = 8'hBE; B = 8'h5E; #100;
A = 8'hBE; B = 8'h5F; #100;
A = 8'hBE; B = 8'h60; #100;
A = 8'hBE; B = 8'h61; #100;
A = 8'hBE; B = 8'h62; #100;
A = 8'hBE; B = 8'h63; #100;
A = 8'hBE; B = 8'h64; #100;
A = 8'hBE; B = 8'h65; #100;
A = 8'hBE; B = 8'h66; #100;
A = 8'hBE; B = 8'h67; #100;
A = 8'hBE; B = 8'h68; #100;
A = 8'hBE; B = 8'h69; #100;
A = 8'hBE; B = 8'h6A; #100;
A = 8'hBE; B = 8'h6B; #100;
A = 8'hBE; B = 8'h6C; #100;
A = 8'hBE; B = 8'h6D; #100;
A = 8'hBE; B = 8'h6E; #100;
A = 8'hBE; B = 8'h6F; #100;
A = 8'hBE; B = 8'h70; #100;
A = 8'hBE; B = 8'h71; #100;
A = 8'hBE; B = 8'h72; #100;
A = 8'hBE; B = 8'h73; #100;
A = 8'hBE; B = 8'h74; #100;
A = 8'hBE; B = 8'h75; #100;
A = 8'hBE; B = 8'h76; #100;
A = 8'hBE; B = 8'h77; #100;
A = 8'hBE; B = 8'h78; #100;
A = 8'hBE; B = 8'h79; #100;
A = 8'hBE; B = 8'h7A; #100;
A = 8'hBE; B = 8'h7B; #100;
A = 8'hBE; B = 8'h7C; #100;
A = 8'hBE; B = 8'h7D; #100;
A = 8'hBE; B = 8'h7E; #100;
A = 8'hBE; B = 8'h7F; #100;
A = 8'hBE; B = 8'h80; #100;
A = 8'hBE; B = 8'h81; #100;
A = 8'hBE; B = 8'h82; #100;
A = 8'hBE; B = 8'h83; #100;
A = 8'hBE; B = 8'h84; #100;
A = 8'hBE; B = 8'h85; #100;
A = 8'hBE; B = 8'h86; #100;
A = 8'hBE; B = 8'h87; #100;
A = 8'hBE; B = 8'h88; #100;
A = 8'hBE; B = 8'h89; #100;
A = 8'hBE; B = 8'h8A; #100;
A = 8'hBE; B = 8'h8B; #100;
A = 8'hBE; B = 8'h8C; #100;
A = 8'hBE; B = 8'h8D; #100;
A = 8'hBE; B = 8'h8E; #100;
A = 8'hBE; B = 8'h8F; #100;
A = 8'hBE; B = 8'h90; #100;
A = 8'hBE; B = 8'h91; #100;
A = 8'hBE; B = 8'h92; #100;
A = 8'hBE; B = 8'h93; #100;
A = 8'hBE; B = 8'h94; #100;
A = 8'hBE; B = 8'h95; #100;
A = 8'hBE; B = 8'h96; #100;
A = 8'hBE; B = 8'h97; #100;
A = 8'hBE; B = 8'h98; #100;
A = 8'hBE; B = 8'h99; #100;
A = 8'hBE; B = 8'h9A; #100;
A = 8'hBE; B = 8'h9B; #100;
A = 8'hBE; B = 8'h9C; #100;
A = 8'hBE; B = 8'h9D; #100;
A = 8'hBE; B = 8'h9E; #100;
A = 8'hBE; B = 8'h9F; #100;
A = 8'hBE; B = 8'hA0; #100;
A = 8'hBE; B = 8'hA1; #100;
A = 8'hBE; B = 8'hA2; #100;
A = 8'hBE; B = 8'hA3; #100;
A = 8'hBE; B = 8'hA4; #100;
A = 8'hBE; B = 8'hA5; #100;
A = 8'hBE; B = 8'hA6; #100;
A = 8'hBE; B = 8'hA7; #100;
A = 8'hBE; B = 8'hA8; #100;
A = 8'hBE; B = 8'hA9; #100;
A = 8'hBE; B = 8'hAA; #100;
A = 8'hBE; B = 8'hAB; #100;
A = 8'hBE; B = 8'hAC; #100;
A = 8'hBE; B = 8'hAD; #100;
A = 8'hBE; B = 8'hAE; #100;
A = 8'hBE; B = 8'hAF; #100;
A = 8'hBE; B = 8'hB0; #100;
A = 8'hBE; B = 8'hB1; #100;
A = 8'hBE; B = 8'hB2; #100;
A = 8'hBE; B = 8'hB3; #100;
A = 8'hBE; B = 8'hB4; #100;
A = 8'hBE; B = 8'hB5; #100;
A = 8'hBE; B = 8'hB6; #100;
A = 8'hBE; B = 8'hB7; #100;
A = 8'hBE; B = 8'hB8; #100;
A = 8'hBE; B = 8'hB9; #100;
A = 8'hBE; B = 8'hBA; #100;
A = 8'hBE; B = 8'hBB; #100;
A = 8'hBE; B = 8'hBC; #100;
A = 8'hBE; B = 8'hBD; #100;
A = 8'hBE; B = 8'hBE; #100;
A = 8'hBE; B = 8'hBF; #100;
A = 8'hBE; B = 8'hC0; #100;
A = 8'hBE; B = 8'hC1; #100;
A = 8'hBE; B = 8'hC2; #100;
A = 8'hBE; B = 8'hC3; #100;
A = 8'hBE; B = 8'hC4; #100;
A = 8'hBE; B = 8'hC5; #100;
A = 8'hBE; B = 8'hC6; #100;
A = 8'hBE; B = 8'hC7; #100;
A = 8'hBE; B = 8'hC8; #100;
A = 8'hBE; B = 8'hC9; #100;
A = 8'hBE; B = 8'hCA; #100;
A = 8'hBE; B = 8'hCB; #100;
A = 8'hBE; B = 8'hCC; #100;
A = 8'hBE; B = 8'hCD; #100;
A = 8'hBE; B = 8'hCE; #100;
A = 8'hBE; B = 8'hCF; #100;
A = 8'hBE; B = 8'hD0; #100;
A = 8'hBE; B = 8'hD1; #100;
A = 8'hBE; B = 8'hD2; #100;
A = 8'hBE; B = 8'hD3; #100;
A = 8'hBE; B = 8'hD4; #100;
A = 8'hBE; B = 8'hD5; #100;
A = 8'hBE; B = 8'hD6; #100;
A = 8'hBE; B = 8'hD7; #100;
A = 8'hBE; B = 8'hD8; #100;
A = 8'hBE; B = 8'hD9; #100;
A = 8'hBE; B = 8'hDA; #100;
A = 8'hBE; B = 8'hDB; #100;
A = 8'hBE; B = 8'hDC; #100;
A = 8'hBE; B = 8'hDD; #100;
A = 8'hBE; B = 8'hDE; #100;
A = 8'hBE; B = 8'hDF; #100;
A = 8'hBE; B = 8'hE0; #100;
A = 8'hBE; B = 8'hE1; #100;
A = 8'hBE; B = 8'hE2; #100;
A = 8'hBE; B = 8'hE3; #100;
A = 8'hBE; B = 8'hE4; #100;
A = 8'hBE; B = 8'hE5; #100;
A = 8'hBE; B = 8'hE6; #100;
A = 8'hBE; B = 8'hE7; #100;
A = 8'hBE; B = 8'hE8; #100;
A = 8'hBE; B = 8'hE9; #100;
A = 8'hBE; B = 8'hEA; #100;
A = 8'hBE; B = 8'hEB; #100;
A = 8'hBE; B = 8'hEC; #100;
A = 8'hBE; B = 8'hED; #100;
A = 8'hBE; B = 8'hEE; #100;
A = 8'hBE; B = 8'hEF; #100;
A = 8'hBE; B = 8'hF0; #100;
A = 8'hBE; B = 8'hF1; #100;
A = 8'hBE; B = 8'hF2; #100;
A = 8'hBE; B = 8'hF3; #100;
A = 8'hBE; B = 8'hF4; #100;
A = 8'hBE; B = 8'hF5; #100;
A = 8'hBE; B = 8'hF6; #100;
A = 8'hBE; B = 8'hF7; #100;
A = 8'hBE; B = 8'hF8; #100;
A = 8'hBE; B = 8'hF9; #100;
A = 8'hBE; B = 8'hFA; #100;
A = 8'hBE; B = 8'hFB; #100;
A = 8'hBE; B = 8'hFC; #100;
A = 8'hBE; B = 8'hFD; #100;
A = 8'hBE; B = 8'hFE; #100;
A = 8'hBE; B = 8'hFF; #100;
A = 8'hBF; B = 8'h0; #100;
A = 8'hBF; B = 8'h1; #100;
A = 8'hBF; B = 8'h2; #100;
A = 8'hBF; B = 8'h3; #100;
A = 8'hBF; B = 8'h4; #100;
A = 8'hBF; B = 8'h5; #100;
A = 8'hBF; B = 8'h6; #100;
A = 8'hBF; B = 8'h7; #100;
A = 8'hBF; B = 8'h8; #100;
A = 8'hBF; B = 8'h9; #100;
A = 8'hBF; B = 8'hA; #100;
A = 8'hBF; B = 8'hB; #100;
A = 8'hBF; B = 8'hC; #100;
A = 8'hBF; B = 8'hD; #100;
A = 8'hBF; B = 8'hE; #100;
A = 8'hBF; B = 8'hF; #100;
A = 8'hBF; B = 8'h10; #100;
A = 8'hBF; B = 8'h11; #100;
A = 8'hBF; B = 8'h12; #100;
A = 8'hBF; B = 8'h13; #100;
A = 8'hBF; B = 8'h14; #100;
A = 8'hBF; B = 8'h15; #100;
A = 8'hBF; B = 8'h16; #100;
A = 8'hBF; B = 8'h17; #100;
A = 8'hBF; B = 8'h18; #100;
A = 8'hBF; B = 8'h19; #100;
A = 8'hBF; B = 8'h1A; #100;
A = 8'hBF; B = 8'h1B; #100;
A = 8'hBF; B = 8'h1C; #100;
A = 8'hBF; B = 8'h1D; #100;
A = 8'hBF; B = 8'h1E; #100;
A = 8'hBF; B = 8'h1F; #100;
A = 8'hBF; B = 8'h20; #100;
A = 8'hBF; B = 8'h21; #100;
A = 8'hBF; B = 8'h22; #100;
A = 8'hBF; B = 8'h23; #100;
A = 8'hBF; B = 8'h24; #100;
A = 8'hBF; B = 8'h25; #100;
A = 8'hBF; B = 8'h26; #100;
A = 8'hBF; B = 8'h27; #100;
A = 8'hBF; B = 8'h28; #100;
A = 8'hBF; B = 8'h29; #100;
A = 8'hBF; B = 8'h2A; #100;
A = 8'hBF; B = 8'h2B; #100;
A = 8'hBF; B = 8'h2C; #100;
A = 8'hBF; B = 8'h2D; #100;
A = 8'hBF; B = 8'h2E; #100;
A = 8'hBF; B = 8'h2F; #100;
A = 8'hBF; B = 8'h30; #100;
A = 8'hBF; B = 8'h31; #100;
A = 8'hBF; B = 8'h32; #100;
A = 8'hBF; B = 8'h33; #100;
A = 8'hBF; B = 8'h34; #100;
A = 8'hBF; B = 8'h35; #100;
A = 8'hBF; B = 8'h36; #100;
A = 8'hBF; B = 8'h37; #100;
A = 8'hBF; B = 8'h38; #100;
A = 8'hBF; B = 8'h39; #100;
A = 8'hBF; B = 8'h3A; #100;
A = 8'hBF; B = 8'h3B; #100;
A = 8'hBF; B = 8'h3C; #100;
A = 8'hBF; B = 8'h3D; #100;
A = 8'hBF; B = 8'h3E; #100;
A = 8'hBF; B = 8'h3F; #100;
A = 8'hBF; B = 8'h40; #100;
A = 8'hBF; B = 8'h41; #100;
A = 8'hBF; B = 8'h42; #100;
A = 8'hBF; B = 8'h43; #100;
A = 8'hBF; B = 8'h44; #100;
A = 8'hBF; B = 8'h45; #100;
A = 8'hBF; B = 8'h46; #100;
A = 8'hBF; B = 8'h47; #100;
A = 8'hBF; B = 8'h48; #100;
A = 8'hBF; B = 8'h49; #100;
A = 8'hBF; B = 8'h4A; #100;
A = 8'hBF; B = 8'h4B; #100;
A = 8'hBF; B = 8'h4C; #100;
A = 8'hBF; B = 8'h4D; #100;
A = 8'hBF; B = 8'h4E; #100;
A = 8'hBF; B = 8'h4F; #100;
A = 8'hBF; B = 8'h50; #100;
A = 8'hBF; B = 8'h51; #100;
A = 8'hBF; B = 8'h52; #100;
A = 8'hBF; B = 8'h53; #100;
A = 8'hBF; B = 8'h54; #100;
A = 8'hBF; B = 8'h55; #100;
A = 8'hBF; B = 8'h56; #100;
A = 8'hBF; B = 8'h57; #100;
A = 8'hBF; B = 8'h58; #100;
A = 8'hBF; B = 8'h59; #100;
A = 8'hBF; B = 8'h5A; #100;
A = 8'hBF; B = 8'h5B; #100;
A = 8'hBF; B = 8'h5C; #100;
A = 8'hBF; B = 8'h5D; #100;
A = 8'hBF; B = 8'h5E; #100;
A = 8'hBF; B = 8'h5F; #100;
A = 8'hBF; B = 8'h60; #100;
A = 8'hBF; B = 8'h61; #100;
A = 8'hBF; B = 8'h62; #100;
A = 8'hBF; B = 8'h63; #100;
A = 8'hBF; B = 8'h64; #100;
A = 8'hBF; B = 8'h65; #100;
A = 8'hBF; B = 8'h66; #100;
A = 8'hBF; B = 8'h67; #100;
A = 8'hBF; B = 8'h68; #100;
A = 8'hBF; B = 8'h69; #100;
A = 8'hBF; B = 8'h6A; #100;
A = 8'hBF; B = 8'h6B; #100;
A = 8'hBF; B = 8'h6C; #100;
A = 8'hBF; B = 8'h6D; #100;
A = 8'hBF; B = 8'h6E; #100;
A = 8'hBF; B = 8'h6F; #100;
A = 8'hBF; B = 8'h70; #100;
A = 8'hBF; B = 8'h71; #100;
A = 8'hBF; B = 8'h72; #100;
A = 8'hBF; B = 8'h73; #100;
A = 8'hBF; B = 8'h74; #100;
A = 8'hBF; B = 8'h75; #100;
A = 8'hBF; B = 8'h76; #100;
A = 8'hBF; B = 8'h77; #100;
A = 8'hBF; B = 8'h78; #100;
A = 8'hBF; B = 8'h79; #100;
A = 8'hBF; B = 8'h7A; #100;
A = 8'hBF; B = 8'h7B; #100;
A = 8'hBF; B = 8'h7C; #100;
A = 8'hBF; B = 8'h7D; #100;
A = 8'hBF; B = 8'h7E; #100;
A = 8'hBF; B = 8'h7F; #100;
A = 8'hBF; B = 8'h80; #100;
A = 8'hBF; B = 8'h81; #100;
A = 8'hBF; B = 8'h82; #100;
A = 8'hBF; B = 8'h83; #100;
A = 8'hBF; B = 8'h84; #100;
A = 8'hBF; B = 8'h85; #100;
A = 8'hBF; B = 8'h86; #100;
A = 8'hBF; B = 8'h87; #100;
A = 8'hBF; B = 8'h88; #100;
A = 8'hBF; B = 8'h89; #100;
A = 8'hBF; B = 8'h8A; #100;
A = 8'hBF; B = 8'h8B; #100;
A = 8'hBF; B = 8'h8C; #100;
A = 8'hBF; B = 8'h8D; #100;
A = 8'hBF; B = 8'h8E; #100;
A = 8'hBF; B = 8'h8F; #100;
A = 8'hBF; B = 8'h90; #100;
A = 8'hBF; B = 8'h91; #100;
A = 8'hBF; B = 8'h92; #100;
A = 8'hBF; B = 8'h93; #100;
A = 8'hBF; B = 8'h94; #100;
A = 8'hBF; B = 8'h95; #100;
A = 8'hBF; B = 8'h96; #100;
A = 8'hBF; B = 8'h97; #100;
A = 8'hBF; B = 8'h98; #100;
A = 8'hBF; B = 8'h99; #100;
A = 8'hBF; B = 8'h9A; #100;
A = 8'hBF; B = 8'h9B; #100;
A = 8'hBF; B = 8'h9C; #100;
A = 8'hBF; B = 8'h9D; #100;
A = 8'hBF; B = 8'h9E; #100;
A = 8'hBF; B = 8'h9F; #100;
A = 8'hBF; B = 8'hA0; #100;
A = 8'hBF; B = 8'hA1; #100;
A = 8'hBF; B = 8'hA2; #100;
A = 8'hBF; B = 8'hA3; #100;
A = 8'hBF; B = 8'hA4; #100;
A = 8'hBF; B = 8'hA5; #100;
A = 8'hBF; B = 8'hA6; #100;
A = 8'hBF; B = 8'hA7; #100;
A = 8'hBF; B = 8'hA8; #100;
A = 8'hBF; B = 8'hA9; #100;
A = 8'hBF; B = 8'hAA; #100;
A = 8'hBF; B = 8'hAB; #100;
A = 8'hBF; B = 8'hAC; #100;
A = 8'hBF; B = 8'hAD; #100;
A = 8'hBF; B = 8'hAE; #100;
A = 8'hBF; B = 8'hAF; #100;
A = 8'hBF; B = 8'hB0; #100;
A = 8'hBF; B = 8'hB1; #100;
A = 8'hBF; B = 8'hB2; #100;
A = 8'hBF; B = 8'hB3; #100;
A = 8'hBF; B = 8'hB4; #100;
A = 8'hBF; B = 8'hB5; #100;
A = 8'hBF; B = 8'hB6; #100;
A = 8'hBF; B = 8'hB7; #100;
A = 8'hBF; B = 8'hB8; #100;
A = 8'hBF; B = 8'hB9; #100;
A = 8'hBF; B = 8'hBA; #100;
A = 8'hBF; B = 8'hBB; #100;
A = 8'hBF; B = 8'hBC; #100;
A = 8'hBF; B = 8'hBD; #100;
A = 8'hBF; B = 8'hBE; #100;
A = 8'hBF; B = 8'hBF; #100;
A = 8'hBF; B = 8'hC0; #100;
A = 8'hBF; B = 8'hC1; #100;
A = 8'hBF; B = 8'hC2; #100;
A = 8'hBF; B = 8'hC3; #100;
A = 8'hBF; B = 8'hC4; #100;
A = 8'hBF; B = 8'hC5; #100;
A = 8'hBF; B = 8'hC6; #100;
A = 8'hBF; B = 8'hC7; #100;
A = 8'hBF; B = 8'hC8; #100;
A = 8'hBF; B = 8'hC9; #100;
A = 8'hBF; B = 8'hCA; #100;
A = 8'hBF; B = 8'hCB; #100;
A = 8'hBF; B = 8'hCC; #100;
A = 8'hBF; B = 8'hCD; #100;
A = 8'hBF; B = 8'hCE; #100;
A = 8'hBF; B = 8'hCF; #100;
A = 8'hBF; B = 8'hD0; #100;
A = 8'hBF; B = 8'hD1; #100;
A = 8'hBF; B = 8'hD2; #100;
A = 8'hBF; B = 8'hD3; #100;
A = 8'hBF; B = 8'hD4; #100;
A = 8'hBF; B = 8'hD5; #100;
A = 8'hBF; B = 8'hD6; #100;
A = 8'hBF; B = 8'hD7; #100;
A = 8'hBF; B = 8'hD8; #100;
A = 8'hBF; B = 8'hD9; #100;
A = 8'hBF; B = 8'hDA; #100;
A = 8'hBF; B = 8'hDB; #100;
A = 8'hBF; B = 8'hDC; #100;
A = 8'hBF; B = 8'hDD; #100;
A = 8'hBF; B = 8'hDE; #100;
A = 8'hBF; B = 8'hDF; #100;
A = 8'hBF; B = 8'hE0; #100;
A = 8'hBF; B = 8'hE1; #100;
A = 8'hBF; B = 8'hE2; #100;
A = 8'hBF; B = 8'hE3; #100;
A = 8'hBF; B = 8'hE4; #100;
A = 8'hBF; B = 8'hE5; #100;
A = 8'hBF; B = 8'hE6; #100;
A = 8'hBF; B = 8'hE7; #100;
A = 8'hBF; B = 8'hE8; #100;
A = 8'hBF; B = 8'hE9; #100;
A = 8'hBF; B = 8'hEA; #100;
A = 8'hBF; B = 8'hEB; #100;
A = 8'hBF; B = 8'hEC; #100;
A = 8'hBF; B = 8'hED; #100;
A = 8'hBF; B = 8'hEE; #100;
A = 8'hBF; B = 8'hEF; #100;
A = 8'hBF; B = 8'hF0; #100;
A = 8'hBF; B = 8'hF1; #100;
A = 8'hBF; B = 8'hF2; #100;
A = 8'hBF; B = 8'hF3; #100;
A = 8'hBF; B = 8'hF4; #100;
A = 8'hBF; B = 8'hF5; #100;
A = 8'hBF; B = 8'hF6; #100;
A = 8'hBF; B = 8'hF7; #100;
A = 8'hBF; B = 8'hF8; #100;
A = 8'hBF; B = 8'hF9; #100;
A = 8'hBF; B = 8'hFA; #100;
A = 8'hBF; B = 8'hFB; #100;
A = 8'hBF; B = 8'hFC; #100;
A = 8'hBF; B = 8'hFD; #100;
A = 8'hBF; B = 8'hFE; #100;
A = 8'hBF; B = 8'hFF; #100;
A = 8'hC0; B = 8'h0; #100;
A = 8'hC0; B = 8'h1; #100;
A = 8'hC0; B = 8'h2; #100;
A = 8'hC0; B = 8'h3; #100;
A = 8'hC0; B = 8'h4; #100;
A = 8'hC0; B = 8'h5; #100;
A = 8'hC0; B = 8'h6; #100;
A = 8'hC0; B = 8'h7; #100;
A = 8'hC0; B = 8'h8; #100;
A = 8'hC0; B = 8'h9; #100;
A = 8'hC0; B = 8'hA; #100;
A = 8'hC0; B = 8'hB; #100;
A = 8'hC0; B = 8'hC; #100;
A = 8'hC0; B = 8'hD; #100;
A = 8'hC0; B = 8'hE; #100;
A = 8'hC0; B = 8'hF; #100;
A = 8'hC0; B = 8'h10; #100;
A = 8'hC0; B = 8'h11; #100;
A = 8'hC0; B = 8'h12; #100;
A = 8'hC0; B = 8'h13; #100;
A = 8'hC0; B = 8'h14; #100;
A = 8'hC0; B = 8'h15; #100;
A = 8'hC0; B = 8'h16; #100;
A = 8'hC0; B = 8'h17; #100;
A = 8'hC0; B = 8'h18; #100;
A = 8'hC0; B = 8'h19; #100;
A = 8'hC0; B = 8'h1A; #100;
A = 8'hC0; B = 8'h1B; #100;
A = 8'hC0; B = 8'h1C; #100;
A = 8'hC0; B = 8'h1D; #100;
A = 8'hC0; B = 8'h1E; #100;
A = 8'hC0; B = 8'h1F; #100;
A = 8'hC0; B = 8'h20; #100;
A = 8'hC0; B = 8'h21; #100;
A = 8'hC0; B = 8'h22; #100;
A = 8'hC0; B = 8'h23; #100;
A = 8'hC0; B = 8'h24; #100;
A = 8'hC0; B = 8'h25; #100;
A = 8'hC0; B = 8'h26; #100;
A = 8'hC0; B = 8'h27; #100;
A = 8'hC0; B = 8'h28; #100;
A = 8'hC0; B = 8'h29; #100;
A = 8'hC0; B = 8'h2A; #100;
A = 8'hC0; B = 8'h2B; #100;
A = 8'hC0; B = 8'h2C; #100;
A = 8'hC0; B = 8'h2D; #100;
A = 8'hC0; B = 8'h2E; #100;
A = 8'hC0; B = 8'h2F; #100;
A = 8'hC0; B = 8'h30; #100;
A = 8'hC0; B = 8'h31; #100;
A = 8'hC0; B = 8'h32; #100;
A = 8'hC0; B = 8'h33; #100;
A = 8'hC0; B = 8'h34; #100;
A = 8'hC0; B = 8'h35; #100;
A = 8'hC0; B = 8'h36; #100;
A = 8'hC0; B = 8'h37; #100;
A = 8'hC0; B = 8'h38; #100;
A = 8'hC0; B = 8'h39; #100;
A = 8'hC0; B = 8'h3A; #100;
A = 8'hC0; B = 8'h3B; #100;
A = 8'hC0; B = 8'h3C; #100;
A = 8'hC0; B = 8'h3D; #100;
A = 8'hC0; B = 8'h3E; #100;
A = 8'hC0; B = 8'h3F; #100;
A = 8'hC0; B = 8'h40; #100;
A = 8'hC0; B = 8'h41; #100;
A = 8'hC0; B = 8'h42; #100;
A = 8'hC0; B = 8'h43; #100;
A = 8'hC0; B = 8'h44; #100;
A = 8'hC0; B = 8'h45; #100;
A = 8'hC0; B = 8'h46; #100;
A = 8'hC0; B = 8'h47; #100;
A = 8'hC0; B = 8'h48; #100;
A = 8'hC0; B = 8'h49; #100;
A = 8'hC0; B = 8'h4A; #100;
A = 8'hC0; B = 8'h4B; #100;
A = 8'hC0; B = 8'h4C; #100;
A = 8'hC0; B = 8'h4D; #100;
A = 8'hC0; B = 8'h4E; #100;
A = 8'hC0; B = 8'h4F; #100;
A = 8'hC0; B = 8'h50; #100;
A = 8'hC0; B = 8'h51; #100;
A = 8'hC0; B = 8'h52; #100;
A = 8'hC0; B = 8'h53; #100;
A = 8'hC0; B = 8'h54; #100;
A = 8'hC0; B = 8'h55; #100;
A = 8'hC0; B = 8'h56; #100;
A = 8'hC0; B = 8'h57; #100;
A = 8'hC0; B = 8'h58; #100;
A = 8'hC0; B = 8'h59; #100;
A = 8'hC0; B = 8'h5A; #100;
A = 8'hC0; B = 8'h5B; #100;
A = 8'hC0; B = 8'h5C; #100;
A = 8'hC0; B = 8'h5D; #100;
A = 8'hC0; B = 8'h5E; #100;
A = 8'hC0; B = 8'h5F; #100;
A = 8'hC0; B = 8'h60; #100;
A = 8'hC0; B = 8'h61; #100;
A = 8'hC0; B = 8'h62; #100;
A = 8'hC0; B = 8'h63; #100;
A = 8'hC0; B = 8'h64; #100;
A = 8'hC0; B = 8'h65; #100;
A = 8'hC0; B = 8'h66; #100;
A = 8'hC0; B = 8'h67; #100;
A = 8'hC0; B = 8'h68; #100;
A = 8'hC0; B = 8'h69; #100;
A = 8'hC0; B = 8'h6A; #100;
A = 8'hC0; B = 8'h6B; #100;
A = 8'hC0; B = 8'h6C; #100;
A = 8'hC0; B = 8'h6D; #100;
A = 8'hC0; B = 8'h6E; #100;
A = 8'hC0; B = 8'h6F; #100;
A = 8'hC0; B = 8'h70; #100;
A = 8'hC0; B = 8'h71; #100;
A = 8'hC0; B = 8'h72; #100;
A = 8'hC0; B = 8'h73; #100;
A = 8'hC0; B = 8'h74; #100;
A = 8'hC0; B = 8'h75; #100;
A = 8'hC0; B = 8'h76; #100;
A = 8'hC0; B = 8'h77; #100;
A = 8'hC0; B = 8'h78; #100;
A = 8'hC0; B = 8'h79; #100;
A = 8'hC0; B = 8'h7A; #100;
A = 8'hC0; B = 8'h7B; #100;
A = 8'hC0; B = 8'h7C; #100;
A = 8'hC0; B = 8'h7D; #100;
A = 8'hC0; B = 8'h7E; #100;
A = 8'hC0; B = 8'h7F; #100;
A = 8'hC0; B = 8'h80; #100;
A = 8'hC0; B = 8'h81; #100;
A = 8'hC0; B = 8'h82; #100;
A = 8'hC0; B = 8'h83; #100;
A = 8'hC0; B = 8'h84; #100;
A = 8'hC0; B = 8'h85; #100;
A = 8'hC0; B = 8'h86; #100;
A = 8'hC0; B = 8'h87; #100;
A = 8'hC0; B = 8'h88; #100;
A = 8'hC0; B = 8'h89; #100;
A = 8'hC0; B = 8'h8A; #100;
A = 8'hC0; B = 8'h8B; #100;
A = 8'hC0; B = 8'h8C; #100;
A = 8'hC0; B = 8'h8D; #100;
A = 8'hC0; B = 8'h8E; #100;
A = 8'hC0; B = 8'h8F; #100;
A = 8'hC0; B = 8'h90; #100;
A = 8'hC0; B = 8'h91; #100;
A = 8'hC0; B = 8'h92; #100;
A = 8'hC0; B = 8'h93; #100;
A = 8'hC0; B = 8'h94; #100;
A = 8'hC0; B = 8'h95; #100;
A = 8'hC0; B = 8'h96; #100;
A = 8'hC0; B = 8'h97; #100;
A = 8'hC0; B = 8'h98; #100;
A = 8'hC0; B = 8'h99; #100;
A = 8'hC0; B = 8'h9A; #100;
A = 8'hC0; B = 8'h9B; #100;
A = 8'hC0; B = 8'h9C; #100;
A = 8'hC0; B = 8'h9D; #100;
A = 8'hC0; B = 8'h9E; #100;
A = 8'hC0; B = 8'h9F; #100;
A = 8'hC0; B = 8'hA0; #100;
A = 8'hC0; B = 8'hA1; #100;
A = 8'hC0; B = 8'hA2; #100;
A = 8'hC0; B = 8'hA3; #100;
A = 8'hC0; B = 8'hA4; #100;
A = 8'hC0; B = 8'hA5; #100;
A = 8'hC0; B = 8'hA6; #100;
A = 8'hC0; B = 8'hA7; #100;
A = 8'hC0; B = 8'hA8; #100;
A = 8'hC0; B = 8'hA9; #100;
A = 8'hC0; B = 8'hAA; #100;
A = 8'hC0; B = 8'hAB; #100;
A = 8'hC0; B = 8'hAC; #100;
A = 8'hC0; B = 8'hAD; #100;
A = 8'hC0; B = 8'hAE; #100;
A = 8'hC0; B = 8'hAF; #100;
A = 8'hC0; B = 8'hB0; #100;
A = 8'hC0; B = 8'hB1; #100;
A = 8'hC0; B = 8'hB2; #100;
A = 8'hC0; B = 8'hB3; #100;
A = 8'hC0; B = 8'hB4; #100;
A = 8'hC0; B = 8'hB5; #100;
A = 8'hC0; B = 8'hB6; #100;
A = 8'hC0; B = 8'hB7; #100;
A = 8'hC0; B = 8'hB8; #100;
A = 8'hC0; B = 8'hB9; #100;
A = 8'hC0; B = 8'hBA; #100;
A = 8'hC0; B = 8'hBB; #100;
A = 8'hC0; B = 8'hBC; #100;
A = 8'hC0; B = 8'hBD; #100;
A = 8'hC0; B = 8'hBE; #100;
A = 8'hC0; B = 8'hBF; #100;
A = 8'hC0; B = 8'hC0; #100;
A = 8'hC0; B = 8'hC1; #100;
A = 8'hC0; B = 8'hC2; #100;
A = 8'hC0; B = 8'hC3; #100;
A = 8'hC0; B = 8'hC4; #100;
A = 8'hC0; B = 8'hC5; #100;
A = 8'hC0; B = 8'hC6; #100;
A = 8'hC0; B = 8'hC7; #100;
A = 8'hC0; B = 8'hC8; #100;
A = 8'hC0; B = 8'hC9; #100;
A = 8'hC0; B = 8'hCA; #100;
A = 8'hC0; B = 8'hCB; #100;
A = 8'hC0; B = 8'hCC; #100;
A = 8'hC0; B = 8'hCD; #100;
A = 8'hC0; B = 8'hCE; #100;
A = 8'hC0; B = 8'hCF; #100;
A = 8'hC0; B = 8'hD0; #100;
A = 8'hC0; B = 8'hD1; #100;
A = 8'hC0; B = 8'hD2; #100;
A = 8'hC0; B = 8'hD3; #100;
A = 8'hC0; B = 8'hD4; #100;
A = 8'hC0; B = 8'hD5; #100;
A = 8'hC0; B = 8'hD6; #100;
A = 8'hC0; B = 8'hD7; #100;
A = 8'hC0; B = 8'hD8; #100;
A = 8'hC0; B = 8'hD9; #100;
A = 8'hC0; B = 8'hDA; #100;
A = 8'hC0; B = 8'hDB; #100;
A = 8'hC0; B = 8'hDC; #100;
A = 8'hC0; B = 8'hDD; #100;
A = 8'hC0; B = 8'hDE; #100;
A = 8'hC0; B = 8'hDF; #100;
A = 8'hC0; B = 8'hE0; #100;
A = 8'hC0; B = 8'hE1; #100;
A = 8'hC0; B = 8'hE2; #100;
A = 8'hC0; B = 8'hE3; #100;
A = 8'hC0; B = 8'hE4; #100;
A = 8'hC0; B = 8'hE5; #100;
A = 8'hC0; B = 8'hE6; #100;
A = 8'hC0; B = 8'hE7; #100;
A = 8'hC0; B = 8'hE8; #100;
A = 8'hC0; B = 8'hE9; #100;
A = 8'hC0; B = 8'hEA; #100;
A = 8'hC0; B = 8'hEB; #100;
A = 8'hC0; B = 8'hEC; #100;
A = 8'hC0; B = 8'hED; #100;
A = 8'hC0; B = 8'hEE; #100;
A = 8'hC0; B = 8'hEF; #100;
A = 8'hC0; B = 8'hF0; #100;
A = 8'hC0; B = 8'hF1; #100;
A = 8'hC0; B = 8'hF2; #100;
A = 8'hC0; B = 8'hF3; #100;
A = 8'hC0; B = 8'hF4; #100;
A = 8'hC0; B = 8'hF5; #100;
A = 8'hC0; B = 8'hF6; #100;
A = 8'hC0; B = 8'hF7; #100;
A = 8'hC0; B = 8'hF8; #100;
A = 8'hC0; B = 8'hF9; #100;
A = 8'hC0; B = 8'hFA; #100;
A = 8'hC0; B = 8'hFB; #100;
A = 8'hC0; B = 8'hFC; #100;
A = 8'hC0; B = 8'hFD; #100;
A = 8'hC0; B = 8'hFE; #100;
A = 8'hC0; B = 8'hFF; #100;
A = 8'hC1; B = 8'h0; #100;
A = 8'hC1; B = 8'h1; #100;
A = 8'hC1; B = 8'h2; #100;
A = 8'hC1; B = 8'h3; #100;
A = 8'hC1; B = 8'h4; #100;
A = 8'hC1; B = 8'h5; #100;
A = 8'hC1; B = 8'h6; #100;
A = 8'hC1; B = 8'h7; #100;
A = 8'hC1; B = 8'h8; #100;
A = 8'hC1; B = 8'h9; #100;
A = 8'hC1; B = 8'hA; #100;
A = 8'hC1; B = 8'hB; #100;
A = 8'hC1; B = 8'hC; #100;
A = 8'hC1; B = 8'hD; #100;
A = 8'hC1; B = 8'hE; #100;
A = 8'hC1; B = 8'hF; #100;
A = 8'hC1; B = 8'h10; #100;
A = 8'hC1; B = 8'h11; #100;
A = 8'hC1; B = 8'h12; #100;
A = 8'hC1; B = 8'h13; #100;
A = 8'hC1; B = 8'h14; #100;
A = 8'hC1; B = 8'h15; #100;
A = 8'hC1; B = 8'h16; #100;
A = 8'hC1; B = 8'h17; #100;
A = 8'hC1; B = 8'h18; #100;
A = 8'hC1; B = 8'h19; #100;
A = 8'hC1; B = 8'h1A; #100;
A = 8'hC1; B = 8'h1B; #100;
A = 8'hC1; B = 8'h1C; #100;
A = 8'hC1; B = 8'h1D; #100;
A = 8'hC1; B = 8'h1E; #100;
A = 8'hC1; B = 8'h1F; #100;
A = 8'hC1; B = 8'h20; #100;
A = 8'hC1; B = 8'h21; #100;
A = 8'hC1; B = 8'h22; #100;
A = 8'hC1; B = 8'h23; #100;
A = 8'hC1; B = 8'h24; #100;
A = 8'hC1; B = 8'h25; #100;
A = 8'hC1; B = 8'h26; #100;
A = 8'hC1; B = 8'h27; #100;
A = 8'hC1; B = 8'h28; #100;
A = 8'hC1; B = 8'h29; #100;
A = 8'hC1; B = 8'h2A; #100;
A = 8'hC1; B = 8'h2B; #100;
A = 8'hC1; B = 8'h2C; #100;
A = 8'hC1; B = 8'h2D; #100;
A = 8'hC1; B = 8'h2E; #100;
A = 8'hC1; B = 8'h2F; #100;
A = 8'hC1; B = 8'h30; #100;
A = 8'hC1; B = 8'h31; #100;
A = 8'hC1; B = 8'h32; #100;
A = 8'hC1; B = 8'h33; #100;
A = 8'hC1; B = 8'h34; #100;
A = 8'hC1; B = 8'h35; #100;
A = 8'hC1; B = 8'h36; #100;
A = 8'hC1; B = 8'h37; #100;
A = 8'hC1; B = 8'h38; #100;
A = 8'hC1; B = 8'h39; #100;
A = 8'hC1; B = 8'h3A; #100;
A = 8'hC1; B = 8'h3B; #100;
A = 8'hC1; B = 8'h3C; #100;
A = 8'hC1; B = 8'h3D; #100;
A = 8'hC1; B = 8'h3E; #100;
A = 8'hC1; B = 8'h3F; #100;
A = 8'hC1; B = 8'h40; #100;
A = 8'hC1; B = 8'h41; #100;
A = 8'hC1; B = 8'h42; #100;
A = 8'hC1; B = 8'h43; #100;
A = 8'hC1; B = 8'h44; #100;
A = 8'hC1; B = 8'h45; #100;
A = 8'hC1; B = 8'h46; #100;
A = 8'hC1; B = 8'h47; #100;
A = 8'hC1; B = 8'h48; #100;
A = 8'hC1; B = 8'h49; #100;
A = 8'hC1; B = 8'h4A; #100;
A = 8'hC1; B = 8'h4B; #100;
A = 8'hC1; B = 8'h4C; #100;
A = 8'hC1; B = 8'h4D; #100;
A = 8'hC1; B = 8'h4E; #100;
A = 8'hC1; B = 8'h4F; #100;
A = 8'hC1; B = 8'h50; #100;
A = 8'hC1; B = 8'h51; #100;
A = 8'hC1; B = 8'h52; #100;
A = 8'hC1; B = 8'h53; #100;
A = 8'hC1; B = 8'h54; #100;
A = 8'hC1; B = 8'h55; #100;
A = 8'hC1; B = 8'h56; #100;
A = 8'hC1; B = 8'h57; #100;
A = 8'hC1; B = 8'h58; #100;
A = 8'hC1; B = 8'h59; #100;
A = 8'hC1; B = 8'h5A; #100;
A = 8'hC1; B = 8'h5B; #100;
A = 8'hC1; B = 8'h5C; #100;
A = 8'hC1; B = 8'h5D; #100;
A = 8'hC1; B = 8'h5E; #100;
A = 8'hC1; B = 8'h5F; #100;
A = 8'hC1; B = 8'h60; #100;
A = 8'hC1; B = 8'h61; #100;
A = 8'hC1; B = 8'h62; #100;
A = 8'hC1; B = 8'h63; #100;
A = 8'hC1; B = 8'h64; #100;
A = 8'hC1; B = 8'h65; #100;
A = 8'hC1; B = 8'h66; #100;
A = 8'hC1; B = 8'h67; #100;
A = 8'hC1; B = 8'h68; #100;
A = 8'hC1; B = 8'h69; #100;
A = 8'hC1; B = 8'h6A; #100;
A = 8'hC1; B = 8'h6B; #100;
A = 8'hC1; B = 8'h6C; #100;
A = 8'hC1; B = 8'h6D; #100;
A = 8'hC1; B = 8'h6E; #100;
A = 8'hC1; B = 8'h6F; #100;
A = 8'hC1; B = 8'h70; #100;
A = 8'hC1; B = 8'h71; #100;
A = 8'hC1; B = 8'h72; #100;
A = 8'hC1; B = 8'h73; #100;
A = 8'hC1; B = 8'h74; #100;
A = 8'hC1; B = 8'h75; #100;
A = 8'hC1; B = 8'h76; #100;
A = 8'hC1; B = 8'h77; #100;
A = 8'hC1; B = 8'h78; #100;
A = 8'hC1; B = 8'h79; #100;
A = 8'hC1; B = 8'h7A; #100;
A = 8'hC1; B = 8'h7B; #100;
A = 8'hC1; B = 8'h7C; #100;
A = 8'hC1; B = 8'h7D; #100;
A = 8'hC1; B = 8'h7E; #100;
A = 8'hC1; B = 8'h7F; #100;
A = 8'hC1; B = 8'h80; #100;
A = 8'hC1; B = 8'h81; #100;
A = 8'hC1; B = 8'h82; #100;
A = 8'hC1; B = 8'h83; #100;
A = 8'hC1; B = 8'h84; #100;
A = 8'hC1; B = 8'h85; #100;
A = 8'hC1; B = 8'h86; #100;
A = 8'hC1; B = 8'h87; #100;
A = 8'hC1; B = 8'h88; #100;
A = 8'hC1; B = 8'h89; #100;
A = 8'hC1; B = 8'h8A; #100;
A = 8'hC1; B = 8'h8B; #100;
A = 8'hC1; B = 8'h8C; #100;
A = 8'hC1; B = 8'h8D; #100;
A = 8'hC1; B = 8'h8E; #100;
A = 8'hC1; B = 8'h8F; #100;
A = 8'hC1; B = 8'h90; #100;
A = 8'hC1; B = 8'h91; #100;
A = 8'hC1; B = 8'h92; #100;
A = 8'hC1; B = 8'h93; #100;
A = 8'hC1; B = 8'h94; #100;
A = 8'hC1; B = 8'h95; #100;
A = 8'hC1; B = 8'h96; #100;
A = 8'hC1; B = 8'h97; #100;
A = 8'hC1; B = 8'h98; #100;
A = 8'hC1; B = 8'h99; #100;
A = 8'hC1; B = 8'h9A; #100;
A = 8'hC1; B = 8'h9B; #100;
A = 8'hC1; B = 8'h9C; #100;
A = 8'hC1; B = 8'h9D; #100;
A = 8'hC1; B = 8'h9E; #100;
A = 8'hC1; B = 8'h9F; #100;
A = 8'hC1; B = 8'hA0; #100;
A = 8'hC1; B = 8'hA1; #100;
A = 8'hC1; B = 8'hA2; #100;
A = 8'hC1; B = 8'hA3; #100;
A = 8'hC1; B = 8'hA4; #100;
A = 8'hC1; B = 8'hA5; #100;
A = 8'hC1; B = 8'hA6; #100;
A = 8'hC1; B = 8'hA7; #100;
A = 8'hC1; B = 8'hA8; #100;
A = 8'hC1; B = 8'hA9; #100;
A = 8'hC1; B = 8'hAA; #100;
A = 8'hC1; B = 8'hAB; #100;
A = 8'hC1; B = 8'hAC; #100;
A = 8'hC1; B = 8'hAD; #100;
A = 8'hC1; B = 8'hAE; #100;
A = 8'hC1; B = 8'hAF; #100;
A = 8'hC1; B = 8'hB0; #100;
A = 8'hC1; B = 8'hB1; #100;
A = 8'hC1; B = 8'hB2; #100;
A = 8'hC1; B = 8'hB3; #100;
A = 8'hC1; B = 8'hB4; #100;
A = 8'hC1; B = 8'hB5; #100;
A = 8'hC1; B = 8'hB6; #100;
A = 8'hC1; B = 8'hB7; #100;
A = 8'hC1; B = 8'hB8; #100;
A = 8'hC1; B = 8'hB9; #100;
A = 8'hC1; B = 8'hBA; #100;
A = 8'hC1; B = 8'hBB; #100;
A = 8'hC1; B = 8'hBC; #100;
A = 8'hC1; B = 8'hBD; #100;
A = 8'hC1; B = 8'hBE; #100;
A = 8'hC1; B = 8'hBF; #100;
A = 8'hC1; B = 8'hC0; #100;
A = 8'hC1; B = 8'hC1; #100;
A = 8'hC1; B = 8'hC2; #100;
A = 8'hC1; B = 8'hC3; #100;
A = 8'hC1; B = 8'hC4; #100;
A = 8'hC1; B = 8'hC5; #100;
A = 8'hC1; B = 8'hC6; #100;
A = 8'hC1; B = 8'hC7; #100;
A = 8'hC1; B = 8'hC8; #100;
A = 8'hC1; B = 8'hC9; #100;
A = 8'hC1; B = 8'hCA; #100;
A = 8'hC1; B = 8'hCB; #100;
A = 8'hC1; B = 8'hCC; #100;
A = 8'hC1; B = 8'hCD; #100;
A = 8'hC1; B = 8'hCE; #100;
A = 8'hC1; B = 8'hCF; #100;
A = 8'hC1; B = 8'hD0; #100;
A = 8'hC1; B = 8'hD1; #100;
A = 8'hC1; B = 8'hD2; #100;
A = 8'hC1; B = 8'hD3; #100;
A = 8'hC1; B = 8'hD4; #100;
A = 8'hC1; B = 8'hD5; #100;
A = 8'hC1; B = 8'hD6; #100;
A = 8'hC1; B = 8'hD7; #100;
A = 8'hC1; B = 8'hD8; #100;
A = 8'hC1; B = 8'hD9; #100;
A = 8'hC1; B = 8'hDA; #100;
A = 8'hC1; B = 8'hDB; #100;
A = 8'hC1; B = 8'hDC; #100;
A = 8'hC1; B = 8'hDD; #100;
A = 8'hC1; B = 8'hDE; #100;
A = 8'hC1; B = 8'hDF; #100;
A = 8'hC1; B = 8'hE0; #100;
A = 8'hC1; B = 8'hE1; #100;
A = 8'hC1; B = 8'hE2; #100;
A = 8'hC1; B = 8'hE3; #100;
A = 8'hC1; B = 8'hE4; #100;
A = 8'hC1; B = 8'hE5; #100;
A = 8'hC1; B = 8'hE6; #100;
A = 8'hC1; B = 8'hE7; #100;
A = 8'hC1; B = 8'hE8; #100;
A = 8'hC1; B = 8'hE9; #100;
A = 8'hC1; B = 8'hEA; #100;
A = 8'hC1; B = 8'hEB; #100;
A = 8'hC1; B = 8'hEC; #100;
A = 8'hC1; B = 8'hED; #100;
A = 8'hC1; B = 8'hEE; #100;
A = 8'hC1; B = 8'hEF; #100;
A = 8'hC1; B = 8'hF0; #100;
A = 8'hC1; B = 8'hF1; #100;
A = 8'hC1; B = 8'hF2; #100;
A = 8'hC1; B = 8'hF3; #100;
A = 8'hC1; B = 8'hF4; #100;
A = 8'hC1; B = 8'hF5; #100;
A = 8'hC1; B = 8'hF6; #100;
A = 8'hC1; B = 8'hF7; #100;
A = 8'hC1; B = 8'hF8; #100;
A = 8'hC1; B = 8'hF9; #100;
A = 8'hC1; B = 8'hFA; #100;
A = 8'hC1; B = 8'hFB; #100;
A = 8'hC1; B = 8'hFC; #100;
A = 8'hC1; B = 8'hFD; #100;
A = 8'hC1; B = 8'hFE; #100;
A = 8'hC1; B = 8'hFF; #100;
A = 8'hC2; B = 8'h0; #100;
A = 8'hC2; B = 8'h1; #100;
A = 8'hC2; B = 8'h2; #100;
A = 8'hC2; B = 8'h3; #100;
A = 8'hC2; B = 8'h4; #100;
A = 8'hC2; B = 8'h5; #100;
A = 8'hC2; B = 8'h6; #100;
A = 8'hC2; B = 8'h7; #100;
A = 8'hC2; B = 8'h8; #100;
A = 8'hC2; B = 8'h9; #100;
A = 8'hC2; B = 8'hA; #100;
A = 8'hC2; B = 8'hB; #100;
A = 8'hC2; B = 8'hC; #100;
A = 8'hC2; B = 8'hD; #100;
A = 8'hC2; B = 8'hE; #100;
A = 8'hC2; B = 8'hF; #100;
A = 8'hC2; B = 8'h10; #100;
A = 8'hC2; B = 8'h11; #100;
A = 8'hC2; B = 8'h12; #100;
A = 8'hC2; B = 8'h13; #100;
A = 8'hC2; B = 8'h14; #100;
A = 8'hC2; B = 8'h15; #100;
A = 8'hC2; B = 8'h16; #100;
A = 8'hC2; B = 8'h17; #100;
A = 8'hC2; B = 8'h18; #100;
A = 8'hC2; B = 8'h19; #100;
A = 8'hC2; B = 8'h1A; #100;
A = 8'hC2; B = 8'h1B; #100;
A = 8'hC2; B = 8'h1C; #100;
A = 8'hC2; B = 8'h1D; #100;
A = 8'hC2; B = 8'h1E; #100;
A = 8'hC2; B = 8'h1F; #100;
A = 8'hC2; B = 8'h20; #100;
A = 8'hC2; B = 8'h21; #100;
A = 8'hC2; B = 8'h22; #100;
A = 8'hC2; B = 8'h23; #100;
A = 8'hC2; B = 8'h24; #100;
A = 8'hC2; B = 8'h25; #100;
A = 8'hC2; B = 8'h26; #100;
A = 8'hC2; B = 8'h27; #100;
A = 8'hC2; B = 8'h28; #100;
A = 8'hC2; B = 8'h29; #100;
A = 8'hC2; B = 8'h2A; #100;
A = 8'hC2; B = 8'h2B; #100;
A = 8'hC2; B = 8'h2C; #100;
A = 8'hC2; B = 8'h2D; #100;
A = 8'hC2; B = 8'h2E; #100;
A = 8'hC2; B = 8'h2F; #100;
A = 8'hC2; B = 8'h30; #100;
A = 8'hC2; B = 8'h31; #100;
A = 8'hC2; B = 8'h32; #100;
A = 8'hC2; B = 8'h33; #100;
A = 8'hC2; B = 8'h34; #100;
A = 8'hC2; B = 8'h35; #100;
A = 8'hC2; B = 8'h36; #100;
A = 8'hC2; B = 8'h37; #100;
A = 8'hC2; B = 8'h38; #100;
A = 8'hC2; B = 8'h39; #100;
A = 8'hC2; B = 8'h3A; #100;
A = 8'hC2; B = 8'h3B; #100;
A = 8'hC2; B = 8'h3C; #100;
A = 8'hC2; B = 8'h3D; #100;
A = 8'hC2; B = 8'h3E; #100;
A = 8'hC2; B = 8'h3F; #100;
A = 8'hC2; B = 8'h40; #100;
A = 8'hC2; B = 8'h41; #100;
A = 8'hC2; B = 8'h42; #100;
A = 8'hC2; B = 8'h43; #100;
A = 8'hC2; B = 8'h44; #100;
A = 8'hC2; B = 8'h45; #100;
A = 8'hC2; B = 8'h46; #100;
A = 8'hC2; B = 8'h47; #100;
A = 8'hC2; B = 8'h48; #100;
A = 8'hC2; B = 8'h49; #100;
A = 8'hC2; B = 8'h4A; #100;
A = 8'hC2; B = 8'h4B; #100;
A = 8'hC2; B = 8'h4C; #100;
A = 8'hC2; B = 8'h4D; #100;
A = 8'hC2; B = 8'h4E; #100;
A = 8'hC2; B = 8'h4F; #100;
A = 8'hC2; B = 8'h50; #100;
A = 8'hC2; B = 8'h51; #100;
A = 8'hC2; B = 8'h52; #100;
A = 8'hC2; B = 8'h53; #100;
A = 8'hC2; B = 8'h54; #100;
A = 8'hC2; B = 8'h55; #100;
A = 8'hC2; B = 8'h56; #100;
A = 8'hC2; B = 8'h57; #100;
A = 8'hC2; B = 8'h58; #100;
A = 8'hC2; B = 8'h59; #100;
A = 8'hC2; B = 8'h5A; #100;
A = 8'hC2; B = 8'h5B; #100;
A = 8'hC2; B = 8'h5C; #100;
A = 8'hC2; B = 8'h5D; #100;
A = 8'hC2; B = 8'h5E; #100;
A = 8'hC2; B = 8'h5F; #100;
A = 8'hC2; B = 8'h60; #100;
A = 8'hC2; B = 8'h61; #100;
A = 8'hC2; B = 8'h62; #100;
A = 8'hC2; B = 8'h63; #100;
A = 8'hC2; B = 8'h64; #100;
A = 8'hC2; B = 8'h65; #100;
A = 8'hC2; B = 8'h66; #100;
A = 8'hC2; B = 8'h67; #100;
A = 8'hC2; B = 8'h68; #100;
A = 8'hC2; B = 8'h69; #100;
A = 8'hC2; B = 8'h6A; #100;
A = 8'hC2; B = 8'h6B; #100;
A = 8'hC2; B = 8'h6C; #100;
A = 8'hC2; B = 8'h6D; #100;
A = 8'hC2; B = 8'h6E; #100;
A = 8'hC2; B = 8'h6F; #100;
A = 8'hC2; B = 8'h70; #100;
A = 8'hC2; B = 8'h71; #100;
A = 8'hC2; B = 8'h72; #100;
A = 8'hC2; B = 8'h73; #100;
A = 8'hC2; B = 8'h74; #100;
A = 8'hC2; B = 8'h75; #100;
A = 8'hC2; B = 8'h76; #100;
A = 8'hC2; B = 8'h77; #100;
A = 8'hC2; B = 8'h78; #100;
A = 8'hC2; B = 8'h79; #100;
A = 8'hC2; B = 8'h7A; #100;
A = 8'hC2; B = 8'h7B; #100;
A = 8'hC2; B = 8'h7C; #100;
A = 8'hC2; B = 8'h7D; #100;
A = 8'hC2; B = 8'h7E; #100;
A = 8'hC2; B = 8'h7F; #100;
A = 8'hC2; B = 8'h80; #100;
A = 8'hC2; B = 8'h81; #100;
A = 8'hC2; B = 8'h82; #100;
A = 8'hC2; B = 8'h83; #100;
A = 8'hC2; B = 8'h84; #100;
A = 8'hC2; B = 8'h85; #100;
A = 8'hC2; B = 8'h86; #100;
A = 8'hC2; B = 8'h87; #100;
A = 8'hC2; B = 8'h88; #100;
A = 8'hC2; B = 8'h89; #100;
A = 8'hC2; B = 8'h8A; #100;
A = 8'hC2; B = 8'h8B; #100;
A = 8'hC2; B = 8'h8C; #100;
A = 8'hC2; B = 8'h8D; #100;
A = 8'hC2; B = 8'h8E; #100;
A = 8'hC2; B = 8'h8F; #100;
A = 8'hC2; B = 8'h90; #100;
A = 8'hC2; B = 8'h91; #100;
A = 8'hC2; B = 8'h92; #100;
A = 8'hC2; B = 8'h93; #100;
A = 8'hC2; B = 8'h94; #100;
A = 8'hC2; B = 8'h95; #100;
A = 8'hC2; B = 8'h96; #100;
A = 8'hC2; B = 8'h97; #100;
A = 8'hC2; B = 8'h98; #100;
A = 8'hC2; B = 8'h99; #100;
A = 8'hC2; B = 8'h9A; #100;
A = 8'hC2; B = 8'h9B; #100;
A = 8'hC2; B = 8'h9C; #100;
A = 8'hC2; B = 8'h9D; #100;
A = 8'hC2; B = 8'h9E; #100;
A = 8'hC2; B = 8'h9F; #100;
A = 8'hC2; B = 8'hA0; #100;
A = 8'hC2; B = 8'hA1; #100;
A = 8'hC2; B = 8'hA2; #100;
A = 8'hC2; B = 8'hA3; #100;
A = 8'hC2; B = 8'hA4; #100;
A = 8'hC2; B = 8'hA5; #100;
A = 8'hC2; B = 8'hA6; #100;
A = 8'hC2; B = 8'hA7; #100;
A = 8'hC2; B = 8'hA8; #100;
A = 8'hC2; B = 8'hA9; #100;
A = 8'hC2; B = 8'hAA; #100;
A = 8'hC2; B = 8'hAB; #100;
A = 8'hC2; B = 8'hAC; #100;
A = 8'hC2; B = 8'hAD; #100;
A = 8'hC2; B = 8'hAE; #100;
A = 8'hC2; B = 8'hAF; #100;
A = 8'hC2; B = 8'hB0; #100;
A = 8'hC2; B = 8'hB1; #100;
A = 8'hC2; B = 8'hB2; #100;
A = 8'hC2; B = 8'hB3; #100;
A = 8'hC2; B = 8'hB4; #100;
A = 8'hC2; B = 8'hB5; #100;
A = 8'hC2; B = 8'hB6; #100;
A = 8'hC2; B = 8'hB7; #100;
A = 8'hC2; B = 8'hB8; #100;
A = 8'hC2; B = 8'hB9; #100;
A = 8'hC2; B = 8'hBA; #100;
A = 8'hC2; B = 8'hBB; #100;
A = 8'hC2; B = 8'hBC; #100;
A = 8'hC2; B = 8'hBD; #100;
A = 8'hC2; B = 8'hBE; #100;
A = 8'hC2; B = 8'hBF; #100;
A = 8'hC2; B = 8'hC0; #100;
A = 8'hC2; B = 8'hC1; #100;
A = 8'hC2; B = 8'hC2; #100;
A = 8'hC2; B = 8'hC3; #100;
A = 8'hC2; B = 8'hC4; #100;
A = 8'hC2; B = 8'hC5; #100;
A = 8'hC2; B = 8'hC6; #100;
A = 8'hC2; B = 8'hC7; #100;
A = 8'hC2; B = 8'hC8; #100;
A = 8'hC2; B = 8'hC9; #100;
A = 8'hC2; B = 8'hCA; #100;
A = 8'hC2; B = 8'hCB; #100;
A = 8'hC2; B = 8'hCC; #100;
A = 8'hC2; B = 8'hCD; #100;
A = 8'hC2; B = 8'hCE; #100;
A = 8'hC2; B = 8'hCF; #100;
A = 8'hC2; B = 8'hD0; #100;
A = 8'hC2; B = 8'hD1; #100;
A = 8'hC2; B = 8'hD2; #100;
A = 8'hC2; B = 8'hD3; #100;
A = 8'hC2; B = 8'hD4; #100;
A = 8'hC2; B = 8'hD5; #100;
A = 8'hC2; B = 8'hD6; #100;
A = 8'hC2; B = 8'hD7; #100;
A = 8'hC2; B = 8'hD8; #100;
A = 8'hC2; B = 8'hD9; #100;
A = 8'hC2; B = 8'hDA; #100;
A = 8'hC2; B = 8'hDB; #100;
A = 8'hC2; B = 8'hDC; #100;
A = 8'hC2; B = 8'hDD; #100;
A = 8'hC2; B = 8'hDE; #100;
A = 8'hC2; B = 8'hDF; #100;
A = 8'hC2; B = 8'hE0; #100;
A = 8'hC2; B = 8'hE1; #100;
A = 8'hC2; B = 8'hE2; #100;
A = 8'hC2; B = 8'hE3; #100;
A = 8'hC2; B = 8'hE4; #100;
A = 8'hC2; B = 8'hE5; #100;
A = 8'hC2; B = 8'hE6; #100;
A = 8'hC2; B = 8'hE7; #100;
A = 8'hC2; B = 8'hE8; #100;
A = 8'hC2; B = 8'hE9; #100;
A = 8'hC2; B = 8'hEA; #100;
A = 8'hC2; B = 8'hEB; #100;
A = 8'hC2; B = 8'hEC; #100;
A = 8'hC2; B = 8'hED; #100;
A = 8'hC2; B = 8'hEE; #100;
A = 8'hC2; B = 8'hEF; #100;
A = 8'hC2; B = 8'hF0; #100;
A = 8'hC2; B = 8'hF1; #100;
A = 8'hC2; B = 8'hF2; #100;
A = 8'hC2; B = 8'hF3; #100;
A = 8'hC2; B = 8'hF4; #100;
A = 8'hC2; B = 8'hF5; #100;
A = 8'hC2; B = 8'hF6; #100;
A = 8'hC2; B = 8'hF7; #100;
A = 8'hC2; B = 8'hF8; #100;
A = 8'hC2; B = 8'hF9; #100;
A = 8'hC2; B = 8'hFA; #100;
A = 8'hC2; B = 8'hFB; #100;
A = 8'hC2; B = 8'hFC; #100;
A = 8'hC2; B = 8'hFD; #100;
A = 8'hC2; B = 8'hFE; #100;
A = 8'hC2; B = 8'hFF; #100;
A = 8'hC3; B = 8'h0; #100;
A = 8'hC3; B = 8'h1; #100;
A = 8'hC3; B = 8'h2; #100;
A = 8'hC3; B = 8'h3; #100;
A = 8'hC3; B = 8'h4; #100;
A = 8'hC3; B = 8'h5; #100;
A = 8'hC3; B = 8'h6; #100;
A = 8'hC3; B = 8'h7; #100;
A = 8'hC3; B = 8'h8; #100;
A = 8'hC3; B = 8'h9; #100;
A = 8'hC3; B = 8'hA; #100;
A = 8'hC3; B = 8'hB; #100;
A = 8'hC3; B = 8'hC; #100;
A = 8'hC3; B = 8'hD; #100;
A = 8'hC3; B = 8'hE; #100;
A = 8'hC3; B = 8'hF; #100;
A = 8'hC3; B = 8'h10; #100;
A = 8'hC3; B = 8'h11; #100;
A = 8'hC3; B = 8'h12; #100;
A = 8'hC3; B = 8'h13; #100;
A = 8'hC3; B = 8'h14; #100;
A = 8'hC3; B = 8'h15; #100;
A = 8'hC3; B = 8'h16; #100;
A = 8'hC3; B = 8'h17; #100;
A = 8'hC3; B = 8'h18; #100;
A = 8'hC3; B = 8'h19; #100;
A = 8'hC3; B = 8'h1A; #100;
A = 8'hC3; B = 8'h1B; #100;
A = 8'hC3; B = 8'h1C; #100;
A = 8'hC3; B = 8'h1D; #100;
A = 8'hC3; B = 8'h1E; #100;
A = 8'hC3; B = 8'h1F; #100;
A = 8'hC3; B = 8'h20; #100;
A = 8'hC3; B = 8'h21; #100;
A = 8'hC3; B = 8'h22; #100;
A = 8'hC3; B = 8'h23; #100;
A = 8'hC3; B = 8'h24; #100;
A = 8'hC3; B = 8'h25; #100;
A = 8'hC3; B = 8'h26; #100;
A = 8'hC3; B = 8'h27; #100;
A = 8'hC3; B = 8'h28; #100;
A = 8'hC3; B = 8'h29; #100;
A = 8'hC3; B = 8'h2A; #100;
A = 8'hC3; B = 8'h2B; #100;
A = 8'hC3; B = 8'h2C; #100;
A = 8'hC3; B = 8'h2D; #100;
A = 8'hC3; B = 8'h2E; #100;
A = 8'hC3; B = 8'h2F; #100;
A = 8'hC3; B = 8'h30; #100;
A = 8'hC3; B = 8'h31; #100;
A = 8'hC3; B = 8'h32; #100;
A = 8'hC3; B = 8'h33; #100;
A = 8'hC3; B = 8'h34; #100;
A = 8'hC3; B = 8'h35; #100;
A = 8'hC3; B = 8'h36; #100;
A = 8'hC3; B = 8'h37; #100;
A = 8'hC3; B = 8'h38; #100;
A = 8'hC3; B = 8'h39; #100;
A = 8'hC3; B = 8'h3A; #100;
A = 8'hC3; B = 8'h3B; #100;
A = 8'hC3; B = 8'h3C; #100;
A = 8'hC3; B = 8'h3D; #100;
A = 8'hC3; B = 8'h3E; #100;
A = 8'hC3; B = 8'h3F; #100;
A = 8'hC3; B = 8'h40; #100;
A = 8'hC3; B = 8'h41; #100;
A = 8'hC3; B = 8'h42; #100;
A = 8'hC3; B = 8'h43; #100;
A = 8'hC3; B = 8'h44; #100;
A = 8'hC3; B = 8'h45; #100;
A = 8'hC3; B = 8'h46; #100;
A = 8'hC3; B = 8'h47; #100;
A = 8'hC3; B = 8'h48; #100;
A = 8'hC3; B = 8'h49; #100;
A = 8'hC3; B = 8'h4A; #100;
A = 8'hC3; B = 8'h4B; #100;
A = 8'hC3; B = 8'h4C; #100;
A = 8'hC3; B = 8'h4D; #100;
A = 8'hC3; B = 8'h4E; #100;
A = 8'hC3; B = 8'h4F; #100;
A = 8'hC3; B = 8'h50; #100;
A = 8'hC3; B = 8'h51; #100;
A = 8'hC3; B = 8'h52; #100;
A = 8'hC3; B = 8'h53; #100;
A = 8'hC3; B = 8'h54; #100;
A = 8'hC3; B = 8'h55; #100;
A = 8'hC3; B = 8'h56; #100;
A = 8'hC3; B = 8'h57; #100;
A = 8'hC3; B = 8'h58; #100;
A = 8'hC3; B = 8'h59; #100;
A = 8'hC3; B = 8'h5A; #100;
A = 8'hC3; B = 8'h5B; #100;
A = 8'hC3; B = 8'h5C; #100;
A = 8'hC3; B = 8'h5D; #100;
A = 8'hC3; B = 8'h5E; #100;
A = 8'hC3; B = 8'h5F; #100;
A = 8'hC3; B = 8'h60; #100;
A = 8'hC3; B = 8'h61; #100;
A = 8'hC3; B = 8'h62; #100;
A = 8'hC3; B = 8'h63; #100;
A = 8'hC3; B = 8'h64; #100;
A = 8'hC3; B = 8'h65; #100;
A = 8'hC3; B = 8'h66; #100;
A = 8'hC3; B = 8'h67; #100;
A = 8'hC3; B = 8'h68; #100;
A = 8'hC3; B = 8'h69; #100;
A = 8'hC3; B = 8'h6A; #100;
A = 8'hC3; B = 8'h6B; #100;
A = 8'hC3; B = 8'h6C; #100;
A = 8'hC3; B = 8'h6D; #100;
A = 8'hC3; B = 8'h6E; #100;
A = 8'hC3; B = 8'h6F; #100;
A = 8'hC3; B = 8'h70; #100;
A = 8'hC3; B = 8'h71; #100;
A = 8'hC3; B = 8'h72; #100;
A = 8'hC3; B = 8'h73; #100;
A = 8'hC3; B = 8'h74; #100;
A = 8'hC3; B = 8'h75; #100;
A = 8'hC3; B = 8'h76; #100;
A = 8'hC3; B = 8'h77; #100;
A = 8'hC3; B = 8'h78; #100;
A = 8'hC3; B = 8'h79; #100;
A = 8'hC3; B = 8'h7A; #100;
A = 8'hC3; B = 8'h7B; #100;
A = 8'hC3; B = 8'h7C; #100;
A = 8'hC3; B = 8'h7D; #100;
A = 8'hC3; B = 8'h7E; #100;
A = 8'hC3; B = 8'h7F; #100;
A = 8'hC3; B = 8'h80; #100;
A = 8'hC3; B = 8'h81; #100;
A = 8'hC3; B = 8'h82; #100;
A = 8'hC3; B = 8'h83; #100;
A = 8'hC3; B = 8'h84; #100;
A = 8'hC3; B = 8'h85; #100;
A = 8'hC3; B = 8'h86; #100;
A = 8'hC3; B = 8'h87; #100;
A = 8'hC3; B = 8'h88; #100;
A = 8'hC3; B = 8'h89; #100;
A = 8'hC3; B = 8'h8A; #100;
A = 8'hC3; B = 8'h8B; #100;
A = 8'hC3; B = 8'h8C; #100;
A = 8'hC3; B = 8'h8D; #100;
A = 8'hC3; B = 8'h8E; #100;
A = 8'hC3; B = 8'h8F; #100;
A = 8'hC3; B = 8'h90; #100;
A = 8'hC3; B = 8'h91; #100;
A = 8'hC3; B = 8'h92; #100;
A = 8'hC3; B = 8'h93; #100;
A = 8'hC3; B = 8'h94; #100;
A = 8'hC3; B = 8'h95; #100;
A = 8'hC3; B = 8'h96; #100;
A = 8'hC3; B = 8'h97; #100;
A = 8'hC3; B = 8'h98; #100;
A = 8'hC3; B = 8'h99; #100;
A = 8'hC3; B = 8'h9A; #100;
A = 8'hC3; B = 8'h9B; #100;
A = 8'hC3; B = 8'h9C; #100;
A = 8'hC3; B = 8'h9D; #100;
A = 8'hC3; B = 8'h9E; #100;
A = 8'hC3; B = 8'h9F; #100;
A = 8'hC3; B = 8'hA0; #100;
A = 8'hC3; B = 8'hA1; #100;
A = 8'hC3; B = 8'hA2; #100;
A = 8'hC3; B = 8'hA3; #100;
A = 8'hC3; B = 8'hA4; #100;
A = 8'hC3; B = 8'hA5; #100;
A = 8'hC3; B = 8'hA6; #100;
A = 8'hC3; B = 8'hA7; #100;
A = 8'hC3; B = 8'hA8; #100;
A = 8'hC3; B = 8'hA9; #100;
A = 8'hC3; B = 8'hAA; #100;
A = 8'hC3; B = 8'hAB; #100;
A = 8'hC3; B = 8'hAC; #100;
A = 8'hC3; B = 8'hAD; #100;
A = 8'hC3; B = 8'hAE; #100;
A = 8'hC3; B = 8'hAF; #100;
A = 8'hC3; B = 8'hB0; #100;
A = 8'hC3; B = 8'hB1; #100;
A = 8'hC3; B = 8'hB2; #100;
A = 8'hC3; B = 8'hB3; #100;
A = 8'hC3; B = 8'hB4; #100;
A = 8'hC3; B = 8'hB5; #100;
A = 8'hC3; B = 8'hB6; #100;
A = 8'hC3; B = 8'hB7; #100;
A = 8'hC3; B = 8'hB8; #100;
A = 8'hC3; B = 8'hB9; #100;
A = 8'hC3; B = 8'hBA; #100;
A = 8'hC3; B = 8'hBB; #100;
A = 8'hC3; B = 8'hBC; #100;
A = 8'hC3; B = 8'hBD; #100;
A = 8'hC3; B = 8'hBE; #100;
A = 8'hC3; B = 8'hBF; #100;
A = 8'hC3; B = 8'hC0; #100;
A = 8'hC3; B = 8'hC1; #100;
A = 8'hC3; B = 8'hC2; #100;
A = 8'hC3; B = 8'hC3; #100;
A = 8'hC3; B = 8'hC4; #100;
A = 8'hC3; B = 8'hC5; #100;
A = 8'hC3; B = 8'hC6; #100;
A = 8'hC3; B = 8'hC7; #100;
A = 8'hC3; B = 8'hC8; #100;
A = 8'hC3; B = 8'hC9; #100;
A = 8'hC3; B = 8'hCA; #100;
A = 8'hC3; B = 8'hCB; #100;
A = 8'hC3; B = 8'hCC; #100;
A = 8'hC3; B = 8'hCD; #100;
A = 8'hC3; B = 8'hCE; #100;
A = 8'hC3; B = 8'hCF; #100;
A = 8'hC3; B = 8'hD0; #100;
A = 8'hC3; B = 8'hD1; #100;
A = 8'hC3; B = 8'hD2; #100;
A = 8'hC3; B = 8'hD3; #100;
A = 8'hC3; B = 8'hD4; #100;
A = 8'hC3; B = 8'hD5; #100;
A = 8'hC3; B = 8'hD6; #100;
A = 8'hC3; B = 8'hD7; #100;
A = 8'hC3; B = 8'hD8; #100;
A = 8'hC3; B = 8'hD9; #100;
A = 8'hC3; B = 8'hDA; #100;
A = 8'hC3; B = 8'hDB; #100;
A = 8'hC3; B = 8'hDC; #100;
A = 8'hC3; B = 8'hDD; #100;
A = 8'hC3; B = 8'hDE; #100;
A = 8'hC3; B = 8'hDF; #100;
A = 8'hC3; B = 8'hE0; #100;
A = 8'hC3; B = 8'hE1; #100;
A = 8'hC3; B = 8'hE2; #100;
A = 8'hC3; B = 8'hE3; #100;
A = 8'hC3; B = 8'hE4; #100;
A = 8'hC3; B = 8'hE5; #100;
A = 8'hC3; B = 8'hE6; #100;
A = 8'hC3; B = 8'hE7; #100;
A = 8'hC3; B = 8'hE8; #100;
A = 8'hC3; B = 8'hE9; #100;
A = 8'hC3; B = 8'hEA; #100;
A = 8'hC3; B = 8'hEB; #100;
A = 8'hC3; B = 8'hEC; #100;
A = 8'hC3; B = 8'hED; #100;
A = 8'hC3; B = 8'hEE; #100;
A = 8'hC3; B = 8'hEF; #100;
A = 8'hC3; B = 8'hF0; #100;
A = 8'hC3; B = 8'hF1; #100;
A = 8'hC3; B = 8'hF2; #100;
A = 8'hC3; B = 8'hF3; #100;
A = 8'hC3; B = 8'hF4; #100;
A = 8'hC3; B = 8'hF5; #100;
A = 8'hC3; B = 8'hF6; #100;
A = 8'hC3; B = 8'hF7; #100;
A = 8'hC3; B = 8'hF8; #100;
A = 8'hC3; B = 8'hF9; #100;
A = 8'hC3; B = 8'hFA; #100;
A = 8'hC3; B = 8'hFB; #100;
A = 8'hC3; B = 8'hFC; #100;
A = 8'hC3; B = 8'hFD; #100;
A = 8'hC3; B = 8'hFE; #100;
A = 8'hC3; B = 8'hFF; #100;
A = 8'hC4; B = 8'h0; #100;
A = 8'hC4; B = 8'h1; #100;
A = 8'hC4; B = 8'h2; #100;
A = 8'hC4; B = 8'h3; #100;
A = 8'hC4; B = 8'h4; #100;
A = 8'hC4; B = 8'h5; #100;
A = 8'hC4; B = 8'h6; #100;
A = 8'hC4; B = 8'h7; #100;
A = 8'hC4; B = 8'h8; #100;
A = 8'hC4; B = 8'h9; #100;
A = 8'hC4; B = 8'hA; #100;
A = 8'hC4; B = 8'hB; #100;
A = 8'hC4; B = 8'hC; #100;
A = 8'hC4; B = 8'hD; #100;
A = 8'hC4; B = 8'hE; #100;
A = 8'hC4; B = 8'hF; #100;
A = 8'hC4; B = 8'h10; #100;
A = 8'hC4; B = 8'h11; #100;
A = 8'hC4; B = 8'h12; #100;
A = 8'hC4; B = 8'h13; #100;
A = 8'hC4; B = 8'h14; #100;
A = 8'hC4; B = 8'h15; #100;
A = 8'hC4; B = 8'h16; #100;
A = 8'hC4; B = 8'h17; #100;
A = 8'hC4; B = 8'h18; #100;
A = 8'hC4; B = 8'h19; #100;
A = 8'hC4; B = 8'h1A; #100;
A = 8'hC4; B = 8'h1B; #100;
A = 8'hC4; B = 8'h1C; #100;
A = 8'hC4; B = 8'h1D; #100;
A = 8'hC4; B = 8'h1E; #100;
A = 8'hC4; B = 8'h1F; #100;
A = 8'hC4; B = 8'h20; #100;
A = 8'hC4; B = 8'h21; #100;
A = 8'hC4; B = 8'h22; #100;
A = 8'hC4; B = 8'h23; #100;
A = 8'hC4; B = 8'h24; #100;
A = 8'hC4; B = 8'h25; #100;
A = 8'hC4; B = 8'h26; #100;
A = 8'hC4; B = 8'h27; #100;
A = 8'hC4; B = 8'h28; #100;
A = 8'hC4; B = 8'h29; #100;
A = 8'hC4; B = 8'h2A; #100;
A = 8'hC4; B = 8'h2B; #100;
A = 8'hC4; B = 8'h2C; #100;
A = 8'hC4; B = 8'h2D; #100;
A = 8'hC4; B = 8'h2E; #100;
A = 8'hC4; B = 8'h2F; #100;
A = 8'hC4; B = 8'h30; #100;
A = 8'hC4; B = 8'h31; #100;
A = 8'hC4; B = 8'h32; #100;
A = 8'hC4; B = 8'h33; #100;
A = 8'hC4; B = 8'h34; #100;
A = 8'hC4; B = 8'h35; #100;
A = 8'hC4; B = 8'h36; #100;
A = 8'hC4; B = 8'h37; #100;
A = 8'hC4; B = 8'h38; #100;
A = 8'hC4; B = 8'h39; #100;
A = 8'hC4; B = 8'h3A; #100;
A = 8'hC4; B = 8'h3B; #100;
A = 8'hC4; B = 8'h3C; #100;
A = 8'hC4; B = 8'h3D; #100;
A = 8'hC4; B = 8'h3E; #100;
A = 8'hC4; B = 8'h3F; #100;
A = 8'hC4; B = 8'h40; #100;
A = 8'hC4; B = 8'h41; #100;
A = 8'hC4; B = 8'h42; #100;
A = 8'hC4; B = 8'h43; #100;
A = 8'hC4; B = 8'h44; #100;
A = 8'hC4; B = 8'h45; #100;
A = 8'hC4; B = 8'h46; #100;
A = 8'hC4; B = 8'h47; #100;
A = 8'hC4; B = 8'h48; #100;
A = 8'hC4; B = 8'h49; #100;
A = 8'hC4; B = 8'h4A; #100;
A = 8'hC4; B = 8'h4B; #100;
A = 8'hC4; B = 8'h4C; #100;
A = 8'hC4; B = 8'h4D; #100;
A = 8'hC4; B = 8'h4E; #100;
A = 8'hC4; B = 8'h4F; #100;
A = 8'hC4; B = 8'h50; #100;
A = 8'hC4; B = 8'h51; #100;
A = 8'hC4; B = 8'h52; #100;
A = 8'hC4; B = 8'h53; #100;
A = 8'hC4; B = 8'h54; #100;
A = 8'hC4; B = 8'h55; #100;
A = 8'hC4; B = 8'h56; #100;
A = 8'hC4; B = 8'h57; #100;
A = 8'hC4; B = 8'h58; #100;
A = 8'hC4; B = 8'h59; #100;
A = 8'hC4; B = 8'h5A; #100;
A = 8'hC4; B = 8'h5B; #100;
A = 8'hC4; B = 8'h5C; #100;
A = 8'hC4; B = 8'h5D; #100;
A = 8'hC4; B = 8'h5E; #100;
A = 8'hC4; B = 8'h5F; #100;
A = 8'hC4; B = 8'h60; #100;
A = 8'hC4; B = 8'h61; #100;
A = 8'hC4; B = 8'h62; #100;
A = 8'hC4; B = 8'h63; #100;
A = 8'hC4; B = 8'h64; #100;
A = 8'hC4; B = 8'h65; #100;
A = 8'hC4; B = 8'h66; #100;
A = 8'hC4; B = 8'h67; #100;
A = 8'hC4; B = 8'h68; #100;
A = 8'hC4; B = 8'h69; #100;
A = 8'hC4; B = 8'h6A; #100;
A = 8'hC4; B = 8'h6B; #100;
A = 8'hC4; B = 8'h6C; #100;
A = 8'hC4; B = 8'h6D; #100;
A = 8'hC4; B = 8'h6E; #100;
A = 8'hC4; B = 8'h6F; #100;
A = 8'hC4; B = 8'h70; #100;
A = 8'hC4; B = 8'h71; #100;
A = 8'hC4; B = 8'h72; #100;
A = 8'hC4; B = 8'h73; #100;
A = 8'hC4; B = 8'h74; #100;
A = 8'hC4; B = 8'h75; #100;
A = 8'hC4; B = 8'h76; #100;
A = 8'hC4; B = 8'h77; #100;
A = 8'hC4; B = 8'h78; #100;
A = 8'hC4; B = 8'h79; #100;
A = 8'hC4; B = 8'h7A; #100;
A = 8'hC4; B = 8'h7B; #100;
A = 8'hC4; B = 8'h7C; #100;
A = 8'hC4; B = 8'h7D; #100;
A = 8'hC4; B = 8'h7E; #100;
A = 8'hC4; B = 8'h7F; #100;
A = 8'hC4; B = 8'h80; #100;
A = 8'hC4; B = 8'h81; #100;
A = 8'hC4; B = 8'h82; #100;
A = 8'hC4; B = 8'h83; #100;
A = 8'hC4; B = 8'h84; #100;
A = 8'hC4; B = 8'h85; #100;
A = 8'hC4; B = 8'h86; #100;
A = 8'hC4; B = 8'h87; #100;
A = 8'hC4; B = 8'h88; #100;
A = 8'hC4; B = 8'h89; #100;
A = 8'hC4; B = 8'h8A; #100;
A = 8'hC4; B = 8'h8B; #100;
A = 8'hC4; B = 8'h8C; #100;
A = 8'hC4; B = 8'h8D; #100;
A = 8'hC4; B = 8'h8E; #100;
A = 8'hC4; B = 8'h8F; #100;
A = 8'hC4; B = 8'h90; #100;
A = 8'hC4; B = 8'h91; #100;
A = 8'hC4; B = 8'h92; #100;
A = 8'hC4; B = 8'h93; #100;
A = 8'hC4; B = 8'h94; #100;
A = 8'hC4; B = 8'h95; #100;
A = 8'hC4; B = 8'h96; #100;
A = 8'hC4; B = 8'h97; #100;
A = 8'hC4; B = 8'h98; #100;
A = 8'hC4; B = 8'h99; #100;
A = 8'hC4; B = 8'h9A; #100;
A = 8'hC4; B = 8'h9B; #100;
A = 8'hC4; B = 8'h9C; #100;
A = 8'hC4; B = 8'h9D; #100;
A = 8'hC4; B = 8'h9E; #100;
A = 8'hC4; B = 8'h9F; #100;
A = 8'hC4; B = 8'hA0; #100;
A = 8'hC4; B = 8'hA1; #100;
A = 8'hC4; B = 8'hA2; #100;
A = 8'hC4; B = 8'hA3; #100;
A = 8'hC4; B = 8'hA4; #100;
A = 8'hC4; B = 8'hA5; #100;
A = 8'hC4; B = 8'hA6; #100;
A = 8'hC4; B = 8'hA7; #100;
A = 8'hC4; B = 8'hA8; #100;
A = 8'hC4; B = 8'hA9; #100;
A = 8'hC4; B = 8'hAA; #100;
A = 8'hC4; B = 8'hAB; #100;
A = 8'hC4; B = 8'hAC; #100;
A = 8'hC4; B = 8'hAD; #100;
A = 8'hC4; B = 8'hAE; #100;
A = 8'hC4; B = 8'hAF; #100;
A = 8'hC4; B = 8'hB0; #100;
A = 8'hC4; B = 8'hB1; #100;
A = 8'hC4; B = 8'hB2; #100;
A = 8'hC4; B = 8'hB3; #100;
A = 8'hC4; B = 8'hB4; #100;
A = 8'hC4; B = 8'hB5; #100;
A = 8'hC4; B = 8'hB6; #100;
A = 8'hC4; B = 8'hB7; #100;
A = 8'hC4; B = 8'hB8; #100;
A = 8'hC4; B = 8'hB9; #100;
A = 8'hC4; B = 8'hBA; #100;
A = 8'hC4; B = 8'hBB; #100;
A = 8'hC4; B = 8'hBC; #100;
A = 8'hC4; B = 8'hBD; #100;
A = 8'hC4; B = 8'hBE; #100;
A = 8'hC4; B = 8'hBF; #100;
A = 8'hC4; B = 8'hC0; #100;
A = 8'hC4; B = 8'hC1; #100;
A = 8'hC4; B = 8'hC2; #100;
A = 8'hC4; B = 8'hC3; #100;
A = 8'hC4; B = 8'hC4; #100;
A = 8'hC4; B = 8'hC5; #100;
A = 8'hC4; B = 8'hC6; #100;
A = 8'hC4; B = 8'hC7; #100;
A = 8'hC4; B = 8'hC8; #100;
A = 8'hC4; B = 8'hC9; #100;
A = 8'hC4; B = 8'hCA; #100;
A = 8'hC4; B = 8'hCB; #100;
A = 8'hC4; B = 8'hCC; #100;
A = 8'hC4; B = 8'hCD; #100;
A = 8'hC4; B = 8'hCE; #100;
A = 8'hC4; B = 8'hCF; #100;
A = 8'hC4; B = 8'hD0; #100;
A = 8'hC4; B = 8'hD1; #100;
A = 8'hC4; B = 8'hD2; #100;
A = 8'hC4; B = 8'hD3; #100;
A = 8'hC4; B = 8'hD4; #100;
A = 8'hC4; B = 8'hD5; #100;
A = 8'hC4; B = 8'hD6; #100;
A = 8'hC4; B = 8'hD7; #100;
A = 8'hC4; B = 8'hD8; #100;
A = 8'hC4; B = 8'hD9; #100;
A = 8'hC4; B = 8'hDA; #100;
A = 8'hC4; B = 8'hDB; #100;
A = 8'hC4; B = 8'hDC; #100;
A = 8'hC4; B = 8'hDD; #100;
A = 8'hC4; B = 8'hDE; #100;
A = 8'hC4; B = 8'hDF; #100;
A = 8'hC4; B = 8'hE0; #100;
A = 8'hC4; B = 8'hE1; #100;
A = 8'hC4; B = 8'hE2; #100;
A = 8'hC4; B = 8'hE3; #100;
A = 8'hC4; B = 8'hE4; #100;
A = 8'hC4; B = 8'hE5; #100;
A = 8'hC4; B = 8'hE6; #100;
A = 8'hC4; B = 8'hE7; #100;
A = 8'hC4; B = 8'hE8; #100;
A = 8'hC4; B = 8'hE9; #100;
A = 8'hC4; B = 8'hEA; #100;
A = 8'hC4; B = 8'hEB; #100;
A = 8'hC4; B = 8'hEC; #100;
A = 8'hC4; B = 8'hED; #100;
A = 8'hC4; B = 8'hEE; #100;
A = 8'hC4; B = 8'hEF; #100;
A = 8'hC4; B = 8'hF0; #100;
A = 8'hC4; B = 8'hF1; #100;
A = 8'hC4; B = 8'hF2; #100;
A = 8'hC4; B = 8'hF3; #100;
A = 8'hC4; B = 8'hF4; #100;
A = 8'hC4; B = 8'hF5; #100;
A = 8'hC4; B = 8'hF6; #100;
A = 8'hC4; B = 8'hF7; #100;
A = 8'hC4; B = 8'hF8; #100;
A = 8'hC4; B = 8'hF9; #100;
A = 8'hC4; B = 8'hFA; #100;
A = 8'hC4; B = 8'hFB; #100;
A = 8'hC4; B = 8'hFC; #100;
A = 8'hC4; B = 8'hFD; #100;
A = 8'hC4; B = 8'hFE; #100;
A = 8'hC4; B = 8'hFF; #100;
A = 8'hC5; B = 8'h0; #100;
A = 8'hC5; B = 8'h1; #100;
A = 8'hC5; B = 8'h2; #100;
A = 8'hC5; B = 8'h3; #100;
A = 8'hC5; B = 8'h4; #100;
A = 8'hC5; B = 8'h5; #100;
A = 8'hC5; B = 8'h6; #100;
A = 8'hC5; B = 8'h7; #100;
A = 8'hC5; B = 8'h8; #100;
A = 8'hC5; B = 8'h9; #100;
A = 8'hC5; B = 8'hA; #100;
A = 8'hC5; B = 8'hB; #100;
A = 8'hC5; B = 8'hC; #100;
A = 8'hC5; B = 8'hD; #100;
A = 8'hC5; B = 8'hE; #100;
A = 8'hC5; B = 8'hF; #100;
A = 8'hC5; B = 8'h10; #100;
A = 8'hC5; B = 8'h11; #100;
A = 8'hC5; B = 8'h12; #100;
A = 8'hC5; B = 8'h13; #100;
A = 8'hC5; B = 8'h14; #100;
A = 8'hC5; B = 8'h15; #100;
A = 8'hC5; B = 8'h16; #100;
A = 8'hC5; B = 8'h17; #100;
A = 8'hC5; B = 8'h18; #100;
A = 8'hC5; B = 8'h19; #100;
A = 8'hC5; B = 8'h1A; #100;
A = 8'hC5; B = 8'h1B; #100;
A = 8'hC5; B = 8'h1C; #100;
A = 8'hC5; B = 8'h1D; #100;
A = 8'hC5; B = 8'h1E; #100;
A = 8'hC5; B = 8'h1F; #100;
A = 8'hC5; B = 8'h20; #100;
A = 8'hC5; B = 8'h21; #100;
A = 8'hC5; B = 8'h22; #100;
A = 8'hC5; B = 8'h23; #100;
A = 8'hC5; B = 8'h24; #100;
A = 8'hC5; B = 8'h25; #100;
A = 8'hC5; B = 8'h26; #100;
A = 8'hC5; B = 8'h27; #100;
A = 8'hC5; B = 8'h28; #100;
A = 8'hC5; B = 8'h29; #100;
A = 8'hC5; B = 8'h2A; #100;
A = 8'hC5; B = 8'h2B; #100;
A = 8'hC5; B = 8'h2C; #100;
A = 8'hC5; B = 8'h2D; #100;
A = 8'hC5; B = 8'h2E; #100;
A = 8'hC5; B = 8'h2F; #100;
A = 8'hC5; B = 8'h30; #100;
A = 8'hC5; B = 8'h31; #100;
A = 8'hC5; B = 8'h32; #100;
A = 8'hC5; B = 8'h33; #100;
A = 8'hC5; B = 8'h34; #100;
A = 8'hC5; B = 8'h35; #100;
A = 8'hC5; B = 8'h36; #100;
A = 8'hC5; B = 8'h37; #100;
A = 8'hC5; B = 8'h38; #100;
A = 8'hC5; B = 8'h39; #100;
A = 8'hC5; B = 8'h3A; #100;
A = 8'hC5; B = 8'h3B; #100;
A = 8'hC5; B = 8'h3C; #100;
A = 8'hC5; B = 8'h3D; #100;
A = 8'hC5; B = 8'h3E; #100;
A = 8'hC5; B = 8'h3F; #100;
A = 8'hC5; B = 8'h40; #100;
A = 8'hC5; B = 8'h41; #100;
A = 8'hC5; B = 8'h42; #100;
A = 8'hC5; B = 8'h43; #100;
A = 8'hC5; B = 8'h44; #100;
A = 8'hC5; B = 8'h45; #100;
A = 8'hC5; B = 8'h46; #100;
A = 8'hC5; B = 8'h47; #100;
A = 8'hC5; B = 8'h48; #100;
A = 8'hC5; B = 8'h49; #100;
A = 8'hC5; B = 8'h4A; #100;
A = 8'hC5; B = 8'h4B; #100;
A = 8'hC5; B = 8'h4C; #100;
A = 8'hC5; B = 8'h4D; #100;
A = 8'hC5; B = 8'h4E; #100;
A = 8'hC5; B = 8'h4F; #100;
A = 8'hC5; B = 8'h50; #100;
A = 8'hC5; B = 8'h51; #100;
A = 8'hC5; B = 8'h52; #100;
A = 8'hC5; B = 8'h53; #100;
A = 8'hC5; B = 8'h54; #100;
A = 8'hC5; B = 8'h55; #100;
A = 8'hC5; B = 8'h56; #100;
A = 8'hC5; B = 8'h57; #100;
A = 8'hC5; B = 8'h58; #100;
A = 8'hC5; B = 8'h59; #100;
A = 8'hC5; B = 8'h5A; #100;
A = 8'hC5; B = 8'h5B; #100;
A = 8'hC5; B = 8'h5C; #100;
A = 8'hC5; B = 8'h5D; #100;
A = 8'hC5; B = 8'h5E; #100;
A = 8'hC5; B = 8'h5F; #100;
A = 8'hC5; B = 8'h60; #100;
A = 8'hC5; B = 8'h61; #100;
A = 8'hC5; B = 8'h62; #100;
A = 8'hC5; B = 8'h63; #100;
A = 8'hC5; B = 8'h64; #100;
A = 8'hC5; B = 8'h65; #100;
A = 8'hC5; B = 8'h66; #100;
A = 8'hC5; B = 8'h67; #100;
A = 8'hC5; B = 8'h68; #100;
A = 8'hC5; B = 8'h69; #100;
A = 8'hC5; B = 8'h6A; #100;
A = 8'hC5; B = 8'h6B; #100;
A = 8'hC5; B = 8'h6C; #100;
A = 8'hC5; B = 8'h6D; #100;
A = 8'hC5; B = 8'h6E; #100;
A = 8'hC5; B = 8'h6F; #100;
A = 8'hC5; B = 8'h70; #100;
A = 8'hC5; B = 8'h71; #100;
A = 8'hC5; B = 8'h72; #100;
A = 8'hC5; B = 8'h73; #100;
A = 8'hC5; B = 8'h74; #100;
A = 8'hC5; B = 8'h75; #100;
A = 8'hC5; B = 8'h76; #100;
A = 8'hC5; B = 8'h77; #100;
A = 8'hC5; B = 8'h78; #100;
A = 8'hC5; B = 8'h79; #100;
A = 8'hC5; B = 8'h7A; #100;
A = 8'hC5; B = 8'h7B; #100;
A = 8'hC5; B = 8'h7C; #100;
A = 8'hC5; B = 8'h7D; #100;
A = 8'hC5; B = 8'h7E; #100;
A = 8'hC5; B = 8'h7F; #100;
A = 8'hC5; B = 8'h80; #100;
A = 8'hC5; B = 8'h81; #100;
A = 8'hC5; B = 8'h82; #100;
A = 8'hC5; B = 8'h83; #100;
A = 8'hC5; B = 8'h84; #100;
A = 8'hC5; B = 8'h85; #100;
A = 8'hC5; B = 8'h86; #100;
A = 8'hC5; B = 8'h87; #100;
A = 8'hC5; B = 8'h88; #100;
A = 8'hC5; B = 8'h89; #100;
A = 8'hC5; B = 8'h8A; #100;
A = 8'hC5; B = 8'h8B; #100;
A = 8'hC5; B = 8'h8C; #100;
A = 8'hC5; B = 8'h8D; #100;
A = 8'hC5; B = 8'h8E; #100;
A = 8'hC5; B = 8'h8F; #100;
A = 8'hC5; B = 8'h90; #100;
A = 8'hC5; B = 8'h91; #100;
A = 8'hC5; B = 8'h92; #100;
A = 8'hC5; B = 8'h93; #100;
A = 8'hC5; B = 8'h94; #100;
A = 8'hC5; B = 8'h95; #100;
A = 8'hC5; B = 8'h96; #100;
A = 8'hC5; B = 8'h97; #100;
A = 8'hC5; B = 8'h98; #100;
A = 8'hC5; B = 8'h99; #100;
A = 8'hC5; B = 8'h9A; #100;
A = 8'hC5; B = 8'h9B; #100;
A = 8'hC5; B = 8'h9C; #100;
A = 8'hC5; B = 8'h9D; #100;
A = 8'hC5; B = 8'h9E; #100;
A = 8'hC5; B = 8'h9F; #100;
A = 8'hC5; B = 8'hA0; #100;
A = 8'hC5; B = 8'hA1; #100;
A = 8'hC5; B = 8'hA2; #100;
A = 8'hC5; B = 8'hA3; #100;
A = 8'hC5; B = 8'hA4; #100;
A = 8'hC5; B = 8'hA5; #100;
A = 8'hC5; B = 8'hA6; #100;
A = 8'hC5; B = 8'hA7; #100;
A = 8'hC5; B = 8'hA8; #100;
A = 8'hC5; B = 8'hA9; #100;
A = 8'hC5; B = 8'hAA; #100;
A = 8'hC5; B = 8'hAB; #100;
A = 8'hC5; B = 8'hAC; #100;
A = 8'hC5; B = 8'hAD; #100;
A = 8'hC5; B = 8'hAE; #100;
A = 8'hC5; B = 8'hAF; #100;
A = 8'hC5; B = 8'hB0; #100;
A = 8'hC5; B = 8'hB1; #100;
A = 8'hC5; B = 8'hB2; #100;
A = 8'hC5; B = 8'hB3; #100;
A = 8'hC5; B = 8'hB4; #100;
A = 8'hC5; B = 8'hB5; #100;
A = 8'hC5; B = 8'hB6; #100;
A = 8'hC5; B = 8'hB7; #100;
A = 8'hC5; B = 8'hB8; #100;
A = 8'hC5; B = 8'hB9; #100;
A = 8'hC5; B = 8'hBA; #100;
A = 8'hC5; B = 8'hBB; #100;
A = 8'hC5; B = 8'hBC; #100;
A = 8'hC5; B = 8'hBD; #100;
A = 8'hC5; B = 8'hBE; #100;
A = 8'hC5; B = 8'hBF; #100;
A = 8'hC5; B = 8'hC0; #100;
A = 8'hC5; B = 8'hC1; #100;
A = 8'hC5; B = 8'hC2; #100;
A = 8'hC5; B = 8'hC3; #100;
A = 8'hC5; B = 8'hC4; #100;
A = 8'hC5; B = 8'hC5; #100;
A = 8'hC5; B = 8'hC6; #100;
A = 8'hC5; B = 8'hC7; #100;
A = 8'hC5; B = 8'hC8; #100;
A = 8'hC5; B = 8'hC9; #100;
A = 8'hC5; B = 8'hCA; #100;
A = 8'hC5; B = 8'hCB; #100;
A = 8'hC5; B = 8'hCC; #100;
A = 8'hC5; B = 8'hCD; #100;
A = 8'hC5; B = 8'hCE; #100;
A = 8'hC5; B = 8'hCF; #100;
A = 8'hC5; B = 8'hD0; #100;
A = 8'hC5; B = 8'hD1; #100;
A = 8'hC5; B = 8'hD2; #100;
A = 8'hC5; B = 8'hD3; #100;
A = 8'hC5; B = 8'hD4; #100;
A = 8'hC5; B = 8'hD5; #100;
A = 8'hC5; B = 8'hD6; #100;
A = 8'hC5; B = 8'hD7; #100;
A = 8'hC5; B = 8'hD8; #100;
A = 8'hC5; B = 8'hD9; #100;
A = 8'hC5; B = 8'hDA; #100;
A = 8'hC5; B = 8'hDB; #100;
A = 8'hC5; B = 8'hDC; #100;
A = 8'hC5; B = 8'hDD; #100;
A = 8'hC5; B = 8'hDE; #100;
A = 8'hC5; B = 8'hDF; #100;
A = 8'hC5; B = 8'hE0; #100;
A = 8'hC5; B = 8'hE1; #100;
A = 8'hC5; B = 8'hE2; #100;
A = 8'hC5; B = 8'hE3; #100;
A = 8'hC5; B = 8'hE4; #100;
A = 8'hC5; B = 8'hE5; #100;
A = 8'hC5; B = 8'hE6; #100;
A = 8'hC5; B = 8'hE7; #100;
A = 8'hC5; B = 8'hE8; #100;
A = 8'hC5; B = 8'hE9; #100;
A = 8'hC5; B = 8'hEA; #100;
A = 8'hC5; B = 8'hEB; #100;
A = 8'hC5; B = 8'hEC; #100;
A = 8'hC5; B = 8'hED; #100;
A = 8'hC5; B = 8'hEE; #100;
A = 8'hC5; B = 8'hEF; #100;
A = 8'hC5; B = 8'hF0; #100;
A = 8'hC5; B = 8'hF1; #100;
A = 8'hC5; B = 8'hF2; #100;
A = 8'hC5; B = 8'hF3; #100;
A = 8'hC5; B = 8'hF4; #100;
A = 8'hC5; B = 8'hF5; #100;
A = 8'hC5; B = 8'hF6; #100;
A = 8'hC5; B = 8'hF7; #100;
A = 8'hC5; B = 8'hF8; #100;
A = 8'hC5; B = 8'hF9; #100;
A = 8'hC5; B = 8'hFA; #100;
A = 8'hC5; B = 8'hFB; #100;
A = 8'hC5; B = 8'hFC; #100;
A = 8'hC5; B = 8'hFD; #100;
A = 8'hC5; B = 8'hFE; #100;
A = 8'hC5; B = 8'hFF; #100;
A = 8'hC6; B = 8'h0; #100;
A = 8'hC6; B = 8'h1; #100;
A = 8'hC6; B = 8'h2; #100;
A = 8'hC6; B = 8'h3; #100;
A = 8'hC6; B = 8'h4; #100;
A = 8'hC6; B = 8'h5; #100;
A = 8'hC6; B = 8'h6; #100;
A = 8'hC6; B = 8'h7; #100;
A = 8'hC6; B = 8'h8; #100;
A = 8'hC6; B = 8'h9; #100;
A = 8'hC6; B = 8'hA; #100;
A = 8'hC6; B = 8'hB; #100;
A = 8'hC6; B = 8'hC; #100;
A = 8'hC6; B = 8'hD; #100;
A = 8'hC6; B = 8'hE; #100;
A = 8'hC6; B = 8'hF; #100;
A = 8'hC6; B = 8'h10; #100;
A = 8'hC6; B = 8'h11; #100;
A = 8'hC6; B = 8'h12; #100;
A = 8'hC6; B = 8'h13; #100;
A = 8'hC6; B = 8'h14; #100;
A = 8'hC6; B = 8'h15; #100;
A = 8'hC6; B = 8'h16; #100;
A = 8'hC6; B = 8'h17; #100;
A = 8'hC6; B = 8'h18; #100;
A = 8'hC6; B = 8'h19; #100;
A = 8'hC6; B = 8'h1A; #100;
A = 8'hC6; B = 8'h1B; #100;
A = 8'hC6; B = 8'h1C; #100;
A = 8'hC6; B = 8'h1D; #100;
A = 8'hC6; B = 8'h1E; #100;
A = 8'hC6; B = 8'h1F; #100;
A = 8'hC6; B = 8'h20; #100;
A = 8'hC6; B = 8'h21; #100;
A = 8'hC6; B = 8'h22; #100;
A = 8'hC6; B = 8'h23; #100;
A = 8'hC6; B = 8'h24; #100;
A = 8'hC6; B = 8'h25; #100;
A = 8'hC6; B = 8'h26; #100;
A = 8'hC6; B = 8'h27; #100;
A = 8'hC6; B = 8'h28; #100;
A = 8'hC6; B = 8'h29; #100;
A = 8'hC6; B = 8'h2A; #100;
A = 8'hC6; B = 8'h2B; #100;
A = 8'hC6; B = 8'h2C; #100;
A = 8'hC6; B = 8'h2D; #100;
A = 8'hC6; B = 8'h2E; #100;
A = 8'hC6; B = 8'h2F; #100;
A = 8'hC6; B = 8'h30; #100;
A = 8'hC6; B = 8'h31; #100;
A = 8'hC6; B = 8'h32; #100;
A = 8'hC6; B = 8'h33; #100;
A = 8'hC6; B = 8'h34; #100;
A = 8'hC6; B = 8'h35; #100;
A = 8'hC6; B = 8'h36; #100;
A = 8'hC6; B = 8'h37; #100;
A = 8'hC6; B = 8'h38; #100;
A = 8'hC6; B = 8'h39; #100;
A = 8'hC6; B = 8'h3A; #100;
A = 8'hC6; B = 8'h3B; #100;
A = 8'hC6; B = 8'h3C; #100;
A = 8'hC6; B = 8'h3D; #100;
A = 8'hC6; B = 8'h3E; #100;
A = 8'hC6; B = 8'h3F; #100;
A = 8'hC6; B = 8'h40; #100;
A = 8'hC6; B = 8'h41; #100;
A = 8'hC6; B = 8'h42; #100;
A = 8'hC6; B = 8'h43; #100;
A = 8'hC6; B = 8'h44; #100;
A = 8'hC6; B = 8'h45; #100;
A = 8'hC6; B = 8'h46; #100;
A = 8'hC6; B = 8'h47; #100;
A = 8'hC6; B = 8'h48; #100;
A = 8'hC6; B = 8'h49; #100;
A = 8'hC6; B = 8'h4A; #100;
A = 8'hC6; B = 8'h4B; #100;
A = 8'hC6; B = 8'h4C; #100;
A = 8'hC6; B = 8'h4D; #100;
A = 8'hC6; B = 8'h4E; #100;
A = 8'hC6; B = 8'h4F; #100;
A = 8'hC6; B = 8'h50; #100;
A = 8'hC6; B = 8'h51; #100;
A = 8'hC6; B = 8'h52; #100;
A = 8'hC6; B = 8'h53; #100;
A = 8'hC6; B = 8'h54; #100;
A = 8'hC6; B = 8'h55; #100;
A = 8'hC6; B = 8'h56; #100;
A = 8'hC6; B = 8'h57; #100;
A = 8'hC6; B = 8'h58; #100;
A = 8'hC6; B = 8'h59; #100;
A = 8'hC6; B = 8'h5A; #100;
A = 8'hC6; B = 8'h5B; #100;
A = 8'hC6; B = 8'h5C; #100;
A = 8'hC6; B = 8'h5D; #100;
A = 8'hC6; B = 8'h5E; #100;
A = 8'hC6; B = 8'h5F; #100;
A = 8'hC6; B = 8'h60; #100;
A = 8'hC6; B = 8'h61; #100;
A = 8'hC6; B = 8'h62; #100;
A = 8'hC6; B = 8'h63; #100;
A = 8'hC6; B = 8'h64; #100;
A = 8'hC6; B = 8'h65; #100;
A = 8'hC6; B = 8'h66; #100;
A = 8'hC6; B = 8'h67; #100;
A = 8'hC6; B = 8'h68; #100;
A = 8'hC6; B = 8'h69; #100;
A = 8'hC6; B = 8'h6A; #100;
A = 8'hC6; B = 8'h6B; #100;
A = 8'hC6; B = 8'h6C; #100;
A = 8'hC6; B = 8'h6D; #100;
A = 8'hC6; B = 8'h6E; #100;
A = 8'hC6; B = 8'h6F; #100;
A = 8'hC6; B = 8'h70; #100;
A = 8'hC6; B = 8'h71; #100;
A = 8'hC6; B = 8'h72; #100;
A = 8'hC6; B = 8'h73; #100;
A = 8'hC6; B = 8'h74; #100;
A = 8'hC6; B = 8'h75; #100;
A = 8'hC6; B = 8'h76; #100;
A = 8'hC6; B = 8'h77; #100;
A = 8'hC6; B = 8'h78; #100;
A = 8'hC6; B = 8'h79; #100;
A = 8'hC6; B = 8'h7A; #100;
A = 8'hC6; B = 8'h7B; #100;
A = 8'hC6; B = 8'h7C; #100;
A = 8'hC6; B = 8'h7D; #100;
A = 8'hC6; B = 8'h7E; #100;
A = 8'hC6; B = 8'h7F; #100;
A = 8'hC6; B = 8'h80; #100;
A = 8'hC6; B = 8'h81; #100;
A = 8'hC6; B = 8'h82; #100;
A = 8'hC6; B = 8'h83; #100;
A = 8'hC6; B = 8'h84; #100;
A = 8'hC6; B = 8'h85; #100;
A = 8'hC6; B = 8'h86; #100;
A = 8'hC6; B = 8'h87; #100;
A = 8'hC6; B = 8'h88; #100;
A = 8'hC6; B = 8'h89; #100;
A = 8'hC6; B = 8'h8A; #100;
A = 8'hC6; B = 8'h8B; #100;
A = 8'hC6; B = 8'h8C; #100;
A = 8'hC6; B = 8'h8D; #100;
A = 8'hC6; B = 8'h8E; #100;
A = 8'hC6; B = 8'h8F; #100;
A = 8'hC6; B = 8'h90; #100;
A = 8'hC6; B = 8'h91; #100;
A = 8'hC6; B = 8'h92; #100;
A = 8'hC6; B = 8'h93; #100;
A = 8'hC6; B = 8'h94; #100;
A = 8'hC6; B = 8'h95; #100;
A = 8'hC6; B = 8'h96; #100;
A = 8'hC6; B = 8'h97; #100;
A = 8'hC6; B = 8'h98; #100;
A = 8'hC6; B = 8'h99; #100;
A = 8'hC6; B = 8'h9A; #100;
A = 8'hC6; B = 8'h9B; #100;
A = 8'hC6; B = 8'h9C; #100;
A = 8'hC6; B = 8'h9D; #100;
A = 8'hC6; B = 8'h9E; #100;
A = 8'hC6; B = 8'h9F; #100;
A = 8'hC6; B = 8'hA0; #100;
A = 8'hC6; B = 8'hA1; #100;
A = 8'hC6; B = 8'hA2; #100;
A = 8'hC6; B = 8'hA3; #100;
A = 8'hC6; B = 8'hA4; #100;
A = 8'hC6; B = 8'hA5; #100;
A = 8'hC6; B = 8'hA6; #100;
A = 8'hC6; B = 8'hA7; #100;
A = 8'hC6; B = 8'hA8; #100;
A = 8'hC6; B = 8'hA9; #100;
A = 8'hC6; B = 8'hAA; #100;
A = 8'hC6; B = 8'hAB; #100;
A = 8'hC6; B = 8'hAC; #100;
A = 8'hC6; B = 8'hAD; #100;
A = 8'hC6; B = 8'hAE; #100;
A = 8'hC6; B = 8'hAF; #100;
A = 8'hC6; B = 8'hB0; #100;
A = 8'hC6; B = 8'hB1; #100;
A = 8'hC6; B = 8'hB2; #100;
A = 8'hC6; B = 8'hB3; #100;
A = 8'hC6; B = 8'hB4; #100;
A = 8'hC6; B = 8'hB5; #100;
A = 8'hC6; B = 8'hB6; #100;
A = 8'hC6; B = 8'hB7; #100;
A = 8'hC6; B = 8'hB8; #100;
A = 8'hC6; B = 8'hB9; #100;
A = 8'hC6; B = 8'hBA; #100;
A = 8'hC6; B = 8'hBB; #100;
A = 8'hC6; B = 8'hBC; #100;
A = 8'hC6; B = 8'hBD; #100;
A = 8'hC6; B = 8'hBE; #100;
A = 8'hC6; B = 8'hBF; #100;
A = 8'hC6; B = 8'hC0; #100;
A = 8'hC6; B = 8'hC1; #100;
A = 8'hC6; B = 8'hC2; #100;
A = 8'hC6; B = 8'hC3; #100;
A = 8'hC6; B = 8'hC4; #100;
A = 8'hC6; B = 8'hC5; #100;
A = 8'hC6; B = 8'hC6; #100;
A = 8'hC6; B = 8'hC7; #100;
A = 8'hC6; B = 8'hC8; #100;
A = 8'hC6; B = 8'hC9; #100;
A = 8'hC6; B = 8'hCA; #100;
A = 8'hC6; B = 8'hCB; #100;
A = 8'hC6; B = 8'hCC; #100;
A = 8'hC6; B = 8'hCD; #100;
A = 8'hC6; B = 8'hCE; #100;
A = 8'hC6; B = 8'hCF; #100;
A = 8'hC6; B = 8'hD0; #100;
A = 8'hC6; B = 8'hD1; #100;
A = 8'hC6; B = 8'hD2; #100;
A = 8'hC6; B = 8'hD3; #100;
A = 8'hC6; B = 8'hD4; #100;
A = 8'hC6; B = 8'hD5; #100;
A = 8'hC6; B = 8'hD6; #100;
A = 8'hC6; B = 8'hD7; #100;
A = 8'hC6; B = 8'hD8; #100;
A = 8'hC6; B = 8'hD9; #100;
A = 8'hC6; B = 8'hDA; #100;
A = 8'hC6; B = 8'hDB; #100;
A = 8'hC6; B = 8'hDC; #100;
A = 8'hC6; B = 8'hDD; #100;
A = 8'hC6; B = 8'hDE; #100;
A = 8'hC6; B = 8'hDF; #100;
A = 8'hC6; B = 8'hE0; #100;
A = 8'hC6; B = 8'hE1; #100;
A = 8'hC6; B = 8'hE2; #100;
A = 8'hC6; B = 8'hE3; #100;
A = 8'hC6; B = 8'hE4; #100;
A = 8'hC6; B = 8'hE5; #100;
A = 8'hC6; B = 8'hE6; #100;
A = 8'hC6; B = 8'hE7; #100;
A = 8'hC6; B = 8'hE8; #100;
A = 8'hC6; B = 8'hE9; #100;
A = 8'hC6; B = 8'hEA; #100;
A = 8'hC6; B = 8'hEB; #100;
A = 8'hC6; B = 8'hEC; #100;
A = 8'hC6; B = 8'hED; #100;
A = 8'hC6; B = 8'hEE; #100;
A = 8'hC6; B = 8'hEF; #100;
A = 8'hC6; B = 8'hF0; #100;
A = 8'hC6; B = 8'hF1; #100;
A = 8'hC6; B = 8'hF2; #100;
A = 8'hC6; B = 8'hF3; #100;
A = 8'hC6; B = 8'hF4; #100;
A = 8'hC6; B = 8'hF5; #100;
A = 8'hC6; B = 8'hF6; #100;
A = 8'hC6; B = 8'hF7; #100;
A = 8'hC6; B = 8'hF8; #100;
A = 8'hC6; B = 8'hF9; #100;
A = 8'hC6; B = 8'hFA; #100;
A = 8'hC6; B = 8'hFB; #100;
A = 8'hC6; B = 8'hFC; #100;
A = 8'hC6; B = 8'hFD; #100;
A = 8'hC6; B = 8'hFE; #100;
A = 8'hC6; B = 8'hFF; #100;
A = 8'hC7; B = 8'h0; #100;
A = 8'hC7; B = 8'h1; #100;
A = 8'hC7; B = 8'h2; #100;
A = 8'hC7; B = 8'h3; #100;
A = 8'hC7; B = 8'h4; #100;
A = 8'hC7; B = 8'h5; #100;
A = 8'hC7; B = 8'h6; #100;
A = 8'hC7; B = 8'h7; #100;
A = 8'hC7; B = 8'h8; #100;
A = 8'hC7; B = 8'h9; #100;
A = 8'hC7; B = 8'hA; #100;
A = 8'hC7; B = 8'hB; #100;
A = 8'hC7; B = 8'hC; #100;
A = 8'hC7; B = 8'hD; #100;
A = 8'hC7; B = 8'hE; #100;
A = 8'hC7; B = 8'hF; #100;
A = 8'hC7; B = 8'h10; #100;
A = 8'hC7; B = 8'h11; #100;
A = 8'hC7; B = 8'h12; #100;
A = 8'hC7; B = 8'h13; #100;
A = 8'hC7; B = 8'h14; #100;
A = 8'hC7; B = 8'h15; #100;
A = 8'hC7; B = 8'h16; #100;
A = 8'hC7; B = 8'h17; #100;
A = 8'hC7; B = 8'h18; #100;
A = 8'hC7; B = 8'h19; #100;
A = 8'hC7; B = 8'h1A; #100;
A = 8'hC7; B = 8'h1B; #100;
A = 8'hC7; B = 8'h1C; #100;
A = 8'hC7; B = 8'h1D; #100;
A = 8'hC7; B = 8'h1E; #100;
A = 8'hC7; B = 8'h1F; #100;
A = 8'hC7; B = 8'h20; #100;
A = 8'hC7; B = 8'h21; #100;
A = 8'hC7; B = 8'h22; #100;
A = 8'hC7; B = 8'h23; #100;
A = 8'hC7; B = 8'h24; #100;
A = 8'hC7; B = 8'h25; #100;
A = 8'hC7; B = 8'h26; #100;
A = 8'hC7; B = 8'h27; #100;
A = 8'hC7; B = 8'h28; #100;
A = 8'hC7; B = 8'h29; #100;
A = 8'hC7; B = 8'h2A; #100;
A = 8'hC7; B = 8'h2B; #100;
A = 8'hC7; B = 8'h2C; #100;
A = 8'hC7; B = 8'h2D; #100;
A = 8'hC7; B = 8'h2E; #100;
A = 8'hC7; B = 8'h2F; #100;
A = 8'hC7; B = 8'h30; #100;
A = 8'hC7; B = 8'h31; #100;
A = 8'hC7; B = 8'h32; #100;
A = 8'hC7; B = 8'h33; #100;
A = 8'hC7; B = 8'h34; #100;
A = 8'hC7; B = 8'h35; #100;
A = 8'hC7; B = 8'h36; #100;
A = 8'hC7; B = 8'h37; #100;
A = 8'hC7; B = 8'h38; #100;
A = 8'hC7; B = 8'h39; #100;
A = 8'hC7; B = 8'h3A; #100;
A = 8'hC7; B = 8'h3B; #100;
A = 8'hC7; B = 8'h3C; #100;
A = 8'hC7; B = 8'h3D; #100;
A = 8'hC7; B = 8'h3E; #100;
A = 8'hC7; B = 8'h3F; #100;
A = 8'hC7; B = 8'h40; #100;
A = 8'hC7; B = 8'h41; #100;
A = 8'hC7; B = 8'h42; #100;
A = 8'hC7; B = 8'h43; #100;
A = 8'hC7; B = 8'h44; #100;
A = 8'hC7; B = 8'h45; #100;
A = 8'hC7; B = 8'h46; #100;
A = 8'hC7; B = 8'h47; #100;
A = 8'hC7; B = 8'h48; #100;
A = 8'hC7; B = 8'h49; #100;
A = 8'hC7; B = 8'h4A; #100;
A = 8'hC7; B = 8'h4B; #100;
A = 8'hC7; B = 8'h4C; #100;
A = 8'hC7; B = 8'h4D; #100;
A = 8'hC7; B = 8'h4E; #100;
A = 8'hC7; B = 8'h4F; #100;
A = 8'hC7; B = 8'h50; #100;
A = 8'hC7; B = 8'h51; #100;
A = 8'hC7; B = 8'h52; #100;
A = 8'hC7; B = 8'h53; #100;
A = 8'hC7; B = 8'h54; #100;
A = 8'hC7; B = 8'h55; #100;
A = 8'hC7; B = 8'h56; #100;
A = 8'hC7; B = 8'h57; #100;
A = 8'hC7; B = 8'h58; #100;
A = 8'hC7; B = 8'h59; #100;
A = 8'hC7; B = 8'h5A; #100;
A = 8'hC7; B = 8'h5B; #100;
A = 8'hC7; B = 8'h5C; #100;
A = 8'hC7; B = 8'h5D; #100;
A = 8'hC7; B = 8'h5E; #100;
A = 8'hC7; B = 8'h5F; #100;
A = 8'hC7; B = 8'h60; #100;
A = 8'hC7; B = 8'h61; #100;
A = 8'hC7; B = 8'h62; #100;
A = 8'hC7; B = 8'h63; #100;
A = 8'hC7; B = 8'h64; #100;
A = 8'hC7; B = 8'h65; #100;
A = 8'hC7; B = 8'h66; #100;
A = 8'hC7; B = 8'h67; #100;
A = 8'hC7; B = 8'h68; #100;
A = 8'hC7; B = 8'h69; #100;
A = 8'hC7; B = 8'h6A; #100;
A = 8'hC7; B = 8'h6B; #100;
A = 8'hC7; B = 8'h6C; #100;
A = 8'hC7; B = 8'h6D; #100;
A = 8'hC7; B = 8'h6E; #100;
A = 8'hC7; B = 8'h6F; #100;
A = 8'hC7; B = 8'h70; #100;
A = 8'hC7; B = 8'h71; #100;
A = 8'hC7; B = 8'h72; #100;
A = 8'hC7; B = 8'h73; #100;
A = 8'hC7; B = 8'h74; #100;
A = 8'hC7; B = 8'h75; #100;
A = 8'hC7; B = 8'h76; #100;
A = 8'hC7; B = 8'h77; #100;
A = 8'hC7; B = 8'h78; #100;
A = 8'hC7; B = 8'h79; #100;
A = 8'hC7; B = 8'h7A; #100;
A = 8'hC7; B = 8'h7B; #100;
A = 8'hC7; B = 8'h7C; #100;
A = 8'hC7; B = 8'h7D; #100;
A = 8'hC7; B = 8'h7E; #100;
A = 8'hC7; B = 8'h7F; #100;
A = 8'hC7; B = 8'h80; #100;
A = 8'hC7; B = 8'h81; #100;
A = 8'hC7; B = 8'h82; #100;
A = 8'hC7; B = 8'h83; #100;
A = 8'hC7; B = 8'h84; #100;
A = 8'hC7; B = 8'h85; #100;
A = 8'hC7; B = 8'h86; #100;
A = 8'hC7; B = 8'h87; #100;
A = 8'hC7; B = 8'h88; #100;
A = 8'hC7; B = 8'h89; #100;
A = 8'hC7; B = 8'h8A; #100;
A = 8'hC7; B = 8'h8B; #100;
A = 8'hC7; B = 8'h8C; #100;
A = 8'hC7; B = 8'h8D; #100;
A = 8'hC7; B = 8'h8E; #100;
A = 8'hC7; B = 8'h8F; #100;
A = 8'hC7; B = 8'h90; #100;
A = 8'hC7; B = 8'h91; #100;
A = 8'hC7; B = 8'h92; #100;
A = 8'hC7; B = 8'h93; #100;
A = 8'hC7; B = 8'h94; #100;
A = 8'hC7; B = 8'h95; #100;
A = 8'hC7; B = 8'h96; #100;
A = 8'hC7; B = 8'h97; #100;
A = 8'hC7; B = 8'h98; #100;
A = 8'hC7; B = 8'h99; #100;
A = 8'hC7; B = 8'h9A; #100;
A = 8'hC7; B = 8'h9B; #100;
A = 8'hC7; B = 8'h9C; #100;
A = 8'hC7; B = 8'h9D; #100;
A = 8'hC7; B = 8'h9E; #100;
A = 8'hC7; B = 8'h9F; #100;
A = 8'hC7; B = 8'hA0; #100;
A = 8'hC7; B = 8'hA1; #100;
A = 8'hC7; B = 8'hA2; #100;
A = 8'hC7; B = 8'hA3; #100;
A = 8'hC7; B = 8'hA4; #100;
A = 8'hC7; B = 8'hA5; #100;
A = 8'hC7; B = 8'hA6; #100;
A = 8'hC7; B = 8'hA7; #100;
A = 8'hC7; B = 8'hA8; #100;
A = 8'hC7; B = 8'hA9; #100;
A = 8'hC7; B = 8'hAA; #100;
A = 8'hC7; B = 8'hAB; #100;
A = 8'hC7; B = 8'hAC; #100;
A = 8'hC7; B = 8'hAD; #100;
A = 8'hC7; B = 8'hAE; #100;
A = 8'hC7; B = 8'hAF; #100;
A = 8'hC7; B = 8'hB0; #100;
A = 8'hC7; B = 8'hB1; #100;
A = 8'hC7; B = 8'hB2; #100;
A = 8'hC7; B = 8'hB3; #100;
A = 8'hC7; B = 8'hB4; #100;
A = 8'hC7; B = 8'hB5; #100;
A = 8'hC7; B = 8'hB6; #100;
A = 8'hC7; B = 8'hB7; #100;
A = 8'hC7; B = 8'hB8; #100;
A = 8'hC7; B = 8'hB9; #100;
A = 8'hC7; B = 8'hBA; #100;
A = 8'hC7; B = 8'hBB; #100;
A = 8'hC7; B = 8'hBC; #100;
A = 8'hC7; B = 8'hBD; #100;
A = 8'hC7; B = 8'hBE; #100;
A = 8'hC7; B = 8'hBF; #100;
A = 8'hC7; B = 8'hC0; #100;
A = 8'hC7; B = 8'hC1; #100;
A = 8'hC7; B = 8'hC2; #100;
A = 8'hC7; B = 8'hC3; #100;
A = 8'hC7; B = 8'hC4; #100;
A = 8'hC7; B = 8'hC5; #100;
A = 8'hC7; B = 8'hC6; #100;
A = 8'hC7; B = 8'hC7; #100;
A = 8'hC7; B = 8'hC8; #100;
A = 8'hC7; B = 8'hC9; #100;
A = 8'hC7; B = 8'hCA; #100;
A = 8'hC7; B = 8'hCB; #100;
A = 8'hC7; B = 8'hCC; #100;
A = 8'hC7; B = 8'hCD; #100;
A = 8'hC7; B = 8'hCE; #100;
A = 8'hC7; B = 8'hCF; #100;
A = 8'hC7; B = 8'hD0; #100;
A = 8'hC7; B = 8'hD1; #100;
A = 8'hC7; B = 8'hD2; #100;
A = 8'hC7; B = 8'hD3; #100;
A = 8'hC7; B = 8'hD4; #100;
A = 8'hC7; B = 8'hD5; #100;
A = 8'hC7; B = 8'hD6; #100;
A = 8'hC7; B = 8'hD7; #100;
A = 8'hC7; B = 8'hD8; #100;
A = 8'hC7; B = 8'hD9; #100;
A = 8'hC7; B = 8'hDA; #100;
A = 8'hC7; B = 8'hDB; #100;
A = 8'hC7; B = 8'hDC; #100;
A = 8'hC7; B = 8'hDD; #100;
A = 8'hC7; B = 8'hDE; #100;
A = 8'hC7; B = 8'hDF; #100;
A = 8'hC7; B = 8'hE0; #100;
A = 8'hC7; B = 8'hE1; #100;
A = 8'hC7; B = 8'hE2; #100;
A = 8'hC7; B = 8'hE3; #100;
A = 8'hC7; B = 8'hE4; #100;
A = 8'hC7; B = 8'hE5; #100;
A = 8'hC7; B = 8'hE6; #100;
A = 8'hC7; B = 8'hE7; #100;
A = 8'hC7; B = 8'hE8; #100;
A = 8'hC7; B = 8'hE9; #100;
A = 8'hC7; B = 8'hEA; #100;
A = 8'hC7; B = 8'hEB; #100;
A = 8'hC7; B = 8'hEC; #100;
A = 8'hC7; B = 8'hED; #100;
A = 8'hC7; B = 8'hEE; #100;
A = 8'hC7; B = 8'hEF; #100;
A = 8'hC7; B = 8'hF0; #100;
A = 8'hC7; B = 8'hF1; #100;
A = 8'hC7; B = 8'hF2; #100;
A = 8'hC7; B = 8'hF3; #100;
A = 8'hC7; B = 8'hF4; #100;
A = 8'hC7; B = 8'hF5; #100;
A = 8'hC7; B = 8'hF6; #100;
A = 8'hC7; B = 8'hF7; #100;
A = 8'hC7; B = 8'hF8; #100;
A = 8'hC7; B = 8'hF9; #100;
A = 8'hC7; B = 8'hFA; #100;
A = 8'hC7; B = 8'hFB; #100;
A = 8'hC7; B = 8'hFC; #100;
A = 8'hC7; B = 8'hFD; #100;
A = 8'hC7; B = 8'hFE; #100;
A = 8'hC7; B = 8'hFF; #100;
A = 8'hC8; B = 8'h0; #100;
A = 8'hC8; B = 8'h1; #100;
A = 8'hC8; B = 8'h2; #100;
A = 8'hC8; B = 8'h3; #100;
A = 8'hC8; B = 8'h4; #100;
A = 8'hC8; B = 8'h5; #100;
A = 8'hC8; B = 8'h6; #100;
A = 8'hC8; B = 8'h7; #100;
A = 8'hC8; B = 8'h8; #100;
A = 8'hC8; B = 8'h9; #100;
A = 8'hC8; B = 8'hA; #100;
A = 8'hC8; B = 8'hB; #100;
A = 8'hC8; B = 8'hC; #100;
A = 8'hC8; B = 8'hD; #100;
A = 8'hC8; B = 8'hE; #100;
A = 8'hC8; B = 8'hF; #100;
A = 8'hC8; B = 8'h10; #100;
A = 8'hC8; B = 8'h11; #100;
A = 8'hC8; B = 8'h12; #100;
A = 8'hC8; B = 8'h13; #100;
A = 8'hC8; B = 8'h14; #100;
A = 8'hC8; B = 8'h15; #100;
A = 8'hC8; B = 8'h16; #100;
A = 8'hC8; B = 8'h17; #100;
A = 8'hC8; B = 8'h18; #100;
A = 8'hC8; B = 8'h19; #100;
A = 8'hC8; B = 8'h1A; #100;
A = 8'hC8; B = 8'h1B; #100;
A = 8'hC8; B = 8'h1C; #100;
A = 8'hC8; B = 8'h1D; #100;
A = 8'hC8; B = 8'h1E; #100;
A = 8'hC8; B = 8'h1F; #100;
A = 8'hC8; B = 8'h20; #100;
A = 8'hC8; B = 8'h21; #100;
A = 8'hC8; B = 8'h22; #100;
A = 8'hC8; B = 8'h23; #100;
A = 8'hC8; B = 8'h24; #100;
A = 8'hC8; B = 8'h25; #100;
A = 8'hC8; B = 8'h26; #100;
A = 8'hC8; B = 8'h27; #100;
A = 8'hC8; B = 8'h28; #100;
A = 8'hC8; B = 8'h29; #100;
A = 8'hC8; B = 8'h2A; #100;
A = 8'hC8; B = 8'h2B; #100;
A = 8'hC8; B = 8'h2C; #100;
A = 8'hC8; B = 8'h2D; #100;
A = 8'hC8; B = 8'h2E; #100;
A = 8'hC8; B = 8'h2F; #100;
A = 8'hC8; B = 8'h30; #100;
A = 8'hC8; B = 8'h31; #100;
A = 8'hC8; B = 8'h32; #100;
A = 8'hC8; B = 8'h33; #100;
A = 8'hC8; B = 8'h34; #100;
A = 8'hC8; B = 8'h35; #100;
A = 8'hC8; B = 8'h36; #100;
A = 8'hC8; B = 8'h37; #100;
A = 8'hC8; B = 8'h38; #100;
A = 8'hC8; B = 8'h39; #100;
A = 8'hC8; B = 8'h3A; #100;
A = 8'hC8; B = 8'h3B; #100;
A = 8'hC8; B = 8'h3C; #100;
A = 8'hC8; B = 8'h3D; #100;
A = 8'hC8; B = 8'h3E; #100;
A = 8'hC8; B = 8'h3F; #100;
A = 8'hC8; B = 8'h40; #100;
A = 8'hC8; B = 8'h41; #100;
A = 8'hC8; B = 8'h42; #100;
A = 8'hC8; B = 8'h43; #100;
A = 8'hC8; B = 8'h44; #100;
A = 8'hC8; B = 8'h45; #100;
A = 8'hC8; B = 8'h46; #100;
A = 8'hC8; B = 8'h47; #100;
A = 8'hC8; B = 8'h48; #100;
A = 8'hC8; B = 8'h49; #100;
A = 8'hC8; B = 8'h4A; #100;
A = 8'hC8; B = 8'h4B; #100;
A = 8'hC8; B = 8'h4C; #100;
A = 8'hC8; B = 8'h4D; #100;
A = 8'hC8; B = 8'h4E; #100;
A = 8'hC8; B = 8'h4F; #100;
A = 8'hC8; B = 8'h50; #100;
A = 8'hC8; B = 8'h51; #100;
A = 8'hC8; B = 8'h52; #100;
A = 8'hC8; B = 8'h53; #100;
A = 8'hC8; B = 8'h54; #100;
A = 8'hC8; B = 8'h55; #100;
A = 8'hC8; B = 8'h56; #100;
A = 8'hC8; B = 8'h57; #100;
A = 8'hC8; B = 8'h58; #100;
A = 8'hC8; B = 8'h59; #100;
A = 8'hC8; B = 8'h5A; #100;
A = 8'hC8; B = 8'h5B; #100;
A = 8'hC8; B = 8'h5C; #100;
A = 8'hC8; B = 8'h5D; #100;
A = 8'hC8; B = 8'h5E; #100;
A = 8'hC8; B = 8'h5F; #100;
A = 8'hC8; B = 8'h60; #100;
A = 8'hC8; B = 8'h61; #100;
A = 8'hC8; B = 8'h62; #100;
A = 8'hC8; B = 8'h63; #100;
A = 8'hC8; B = 8'h64; #100;
A = 8'hC8; B = 8'h65; #100;
A = 8'hC8; B = 8'h66; #100;
A = 8'hC8; B = 8'h67; #100;
A = 8'hC8; B = 8'h68; #100;
A = 8'hC8; B = 8'h69; #100;
A = 8'hC8; B = 8'h6A; #100;
A = 8'hC8; B = 8'h6B; #100;
A = 8'hC8; B = 8'h6C; #100;
A = 8'hC8; B = 8'h6D; #100;
A = 8'hC8; B = 8'h6E; #100;
A = 8'hC8; B = 8'h6F; #100;
A = 8'hC8; B = 8'h70; #100;
A = 8'hC8; B = 8'h71; #100;
A = 8'hC8; B = 8'h72; #100;
A = 8'hC8; B = 8'h73; #100;
A = 8'hC8; B = 8'h74; #100;
A = 8'hC8; B = 8'h75; #100;
A = 8'hC8; B = 8'h76; #100;
A = 8'hC8; B = 8'h77; #100;
A = 8'hC8; B = 8'h78; #100;
A = 8'hC8; B = 8'h79; #100;
A = 8'hC8; B = 8'h7A; #100;
A = 8'hC8; B = 8'h7B; #100;
A = 8'hC8; B = 8'h7C; #100;
A = 8'hC8; B = 8'h7D; #100;
A = 8'hC8; B = 8'h7E; #100;
A = 8'hC8; B = 8'h7F; #100;
A = 8'hC8; B = 8'h80; #100;
A = 8'hC8; B = 8'h81; #100;
A = 8'hC8; B = 8'h82; #100;
A = 8'hC8; B = 8'h83; #100;
A = 8'hC8; B = 8'h84; #100;
A = 8'hC8; B = 8'h85; #100;
A = 8'hC8; B = 8'h86; #100;
A = 8'hC8; B = 8'h87; #100;
A = 8'hC8; B = 8'h88; #100;
A = 8'hC8; B = 8'h89; #100;
A = 8'hC8; B = 8'h8A; #100;
A = 8'hC8; B = 8'h8B; #100;
A = 8'hC8; B = 8'h8C; #100;
A = 8'hC8; B = 8'h8D; #100;
A = 8'hC8; B = 8'h8E; #100;
A = 8'hC8; B = 8'h8F; #100;
A = 8'hC8; B = 8'h90; #100;
A = 8'hC8; B = 8'h91; #100;
A = 8'hC8; B = 8'h92; #100;
A = 8'hC8; B = 8'h93; #100;
A = 8'hC8; B = 8'h94; #100;
A = 8'hC8; B = 8'h95; #100;
A = 8'hC8; B = 8'h96; #100;
A = 8'hC8; B = 8'h97; #100;
A = 8'hC8; B = 8'h98; #100;
A = 8'hC8; B = 8'h99; #100;
A = 8'hC8; B = 8'h9A; #100;
A = 8'hC8; B = 8'h9B; #100;
A = 8'hC8; B = 8'h9C; #100;
A = 8'hC8; B = 8'h9D; #100;
A = 8'hC8; B = 8'h9E; #100;
A = 8'hC8; B = 8'h9F; #100;
A = 8'hC8; B = 8'hA0; #100;
A = 8'hC8; B = 8'hA1; #100;
A = 8'hC8; B = 8'hA2; #100;
A = 8'hC8; B = 8'hA3; #100;
A = 8'hC8; B = 8'hA4; #100;
A = 8'hC8; B = 8'hA5; #100;
A = 8'hC8; B = 8'hA6; #100;
A = 8'hC8; B = 8'hA7; #100;
A = 8'hC8; B = 8'hA8; #100;
A = 8'hC8; B = 8'hA9; #100;
A = 8'hC8; B = 8'hAA; #100;
A = 8'hC8; B = 8'hAB; #100;
A = 8'hC8; B = 8'hAC; #100;
A = 8'hC8; B = 8'hAD; #100;
A = 8'hC8; B = 8'hAE; #100;
A = 8'hC8; B = 8'hAF; #100;
A = 8'hC8; B = 8'hB0; #100;
A = 8'hC8; B = 8'hB1; #100;
A = 8'hC8; B = 8'hB2; #100;
A = 8'hC8; B = 8'hB3; #100;
A = 8'hC8; B = 8'hB4; #100;
A = 8'hC8; B = 8'hB5; #100;
A = 8'hC8; B = 8'hB6; #100;
A = 8'hC8; B = 8'hB7; #100;
A = 8'hC8; B = 8'hB8; #100;
A = 8'hC8; B = 8'hB9; #100;
A = 8'hC8; B = 8'hBA; #100;
A = 8'hC8; B = 8'hBB; #100;
A = 8'hC8; B = 8'hBC; #100;
A = 8'hC8; B = 8'hBD; #100;
A = 8'hC8; B = 8'hBE; #100;
A = 8'hC8; B = 8'hBF; #100;
A = 8'hC8; B = 8'hC0; #100;
A = 8'hC8; B = 8'hC1; #100;
A = 8'hC8; B = 8'hC2; #100;
A = 8'hC8; B = 8'hC3; #100;
A = 8'hC8; B = 8'hC4; #100;
A = 8'hC8; B = 8'hC5; #100;
A = 8'hC8; B = 8'hC6; #100;
A = 8'hC8; B = 8'hC7; #100;
A = 8'hC8; B = 8'hC8; #100;
A = 8'hC8; B = 8'hC9; #100;
A = 8'hC8; B = 8'hCA; #100;
A = 8'hC8; B = 8'hCB; #100;
A = 8'hC8; B = 8'hCC; #100;
A = 8'hC8; B = 8'hCD; #100;
A = 8'hC8; B = 8'hCE; #100;
A = 8'hC8; B = 8'hCF; #100;
A = 8'hC8; B = 8'hD0; #100;
A = 8'hC8; B = 8'hD1; #100;
A = 8'hC8; B = 8'hD2; #100;
A = 8'hC8; B = 8'hD3; #100;
A = 8'hC8; B = 8'hD4; #100;
A = 8'hC8; B = 8'hD5; #100;
A = 8'hC8; B = 8'hD6; #100;
A = 8'hC8; B = 8'hD7; #100;
A = 8'hC8; B = 8'hD8; #100;
A = 8'hC8; B = 8'hD9; #100;
A = 8'hC8; B = 8'hDA; #100;
A = 8'hC8; B = 8'hDB; #100;
A = 8'hC8; B = 8'hDC; #100;
A = 8'hC8; B = 8'hDD; #100;
A = 8'hC8; B = 8'hDE; #100;
A = 8'hC8; B = 8'hDF; #100;
A = 8'hC8; B = 8'hE0; #100;
A = 8'hC8; B = 8'hE1; #100;
A = 8'hC8; B = 8'hE2; #100;
A = 8'hC8; B = 8'hE3; #100;
A = 8'hC8; B = 8'hE4; #100;
A = 8'hC8; B = 8'hE5; #100;
A = 8'hC8; B = 8'hE6; #100;
A = 8'hC8; B = 8'hE7; #100;
A = 8'hC8; B = 8'hE8; #100;
A = 8'hC8; B = 8'hE9; #100;
A = 8'hC8; B = 8'hEA; #100;
A = 8'hC8; B = 8'hEB; #100;
A = 8'hC8; B = 8'hEC; #100;
A = 8'hC8; B = 8'hED; #100;
A = 8'hC8; B = 8'hEE; #100;
A = 8'hC8; B = 8'hEF; #100;
A = 8'hC8; B = 8'hF0; #100;
A = 8'hC8; B = 8'hF1; #100;
A = 8'hC8; B = 8'hF2; #100;
A = 8'hC8; B = 8'hF3; #100;
A = 8'hC8; B = 8'hF4; #100;
A = 8'hC8; B = 8'hF5; #100;
A = 8'hC8; B = 8'hF6; #100;
A = 8'hC8; B = 8'hF7; #100;
A = 8'hC8; B = 8'hF8; #100;
A = 8'hC8; B = 8'hF9; #100;
A = 8'hC8; B = 8'hFA; #100;
A = 8'hC8; B = 8'hFB; #100;
A = 8'hC8; B = 8'hFC; #100;
A = 8'hC8; B = 8'hFD; #100;
A = 8'hC8; B = 8'hFE; #100;
A = 8'hC8; B = 8'hFF; #100;
A = 8'hC9; B = 8'h0; #100;
A = 8'hC9; B = 8'h1; #100;
A = 8'hC9; B = 8'h2; #100;
A = 8'hC9; B = 8'h3; #100;
A = 8'hC9; B = 8'h4; #100;
A = 8'hC9; B = 8'h5; #100;
A = 8'hC9; B = 8'h6; #100;
A = 8'hC9; B = 8'h7; #100;
A = 8'hC9; B = 8'h8; #100;
A = 8'hC9; B = 8'h9; #100;
A = 8'hC9; B = 8'hA; #100;
A = 8'hC9; B = 8'hB; #100;
A = 8'hC9; B = 8'hC; #100;
A = 8'hC9; B = 8'hD; #100;
A = 8'hC9; B = 8'hE; #100;
A = 8'hC9; B = 8'hF; #100;
A = 8'hC9; B = 8'h10; #100;
A = 8'hC9; B = 8'h11; #100;
A = 8'hC9; B = 8'h12; #100;
A = 8'hC9; B = 8'h13; #100;
A = 8'hC9; B = 8'h14; #100;
A = 8'hC9; B = 8'h15; #100;
A = 8'hC9; B = 8'h16; #100;
A = 8'hC9; B = 8'h17; #100;
A = 8'hC9; B = 8'h18; #100;
A = 8'hC9; B = 8'h19; #100;
A = 8'hC9; B = 8'h1A; #100;
A = 8'hC9; B = 8'h1B; #100;
A = 8'hC9; B = 8'h1C; #100;
A = 8'hC9; B = 8'h1D; #100;
A = 8'hC9; B = 8'h1E; #100;
A = 8'hC9; B = 8'h1F; #100;
A = 8'hC9; B = 8'h20; #100;
A = 8'hC9; B = 8'h21; #100;
A = 8'hC9; B = 8'h22; #100;
A = 8'hC9; B = 8'h23; #100;
A = 8'hC9; B = 8'h24; #100;
A = 8'hC9; B = 8'h25; #100;
A = 8'hC9; B = 8'h26; #100;
A = 8'hC9; B = 8'h27; #100;
A = 8'hC9; B = 8'h28; #100;
A = 8'hC9; B = 8'h29; #100;
A = 8'hC9; B = 8'h2A; #100;
A = 8'hC9; B = 8'h2B; #100;
A = 8'hC9; B = 8'h2C; #100;
A = 8'hC9; B = 8'h2D; #100;
A = 8'hC9; B = 8'h2E; #100;
A = 8'hC9; B = 8'h2F; #100;
A = 8'hC9; B = 8'h30; #100;
A = 8'hC9; B = 8'h31; #100;
A = 8'hC9; B = 8'h32; #100;
A = 8'hC9; B = 8'h33; #100;
A = 8'hC9; B = 8'h34; #100;
A = 8'hC9; B = 8'h35; #100;
A = 8'hC9; B = 8'h36; #100;
A = 8'hC9; B = 8'h37; #100;
A = 8'hC9; B = 8'h38; #100;
A = 8'hC9; B = 8'h39; #100;
A = 8'hC9; B = 8'h3A; #100;
A = 8'hC9; B = 8'h3B; #100;
A = 8'hC9; B = 8'h3C; #100;
A = 8'hC9; B = 8'h3D; #100;
A = 8'hC9; B = 8'h3E; #100;
A = 8'hC9; B = 8'h3F; #100;
A = 8'hC9; B = 8'h40; #100;
A = 8'hC9; B = 8'h41; #100;
A = 8'hC9; B = 8'h42; #100;
A = 8'hC9; B = 8'h43; #100;
A = 8'hC9; B = 8'h44; #100;
A = 8'hC9; B = 8'h45; #100;
A = 8'hC9; B = 8'h46; #100;
A = 8'hC9; B = 8'h47; #100;
A = 8'hC9; B = 8'h48; #100;
A = 8'hC9; B = 8'h49; #100;
A = 8'hC9; B = 8'h4A; #100;
A = 8'hC9; B = 8'h4B; #100;
A = 8'hC9; B = 8'h4C; #100;
A = 8'hC9; B = 8'h4D; #100;
A = 8'hC9; B = 8'h4E; #100;
A = 8'hC9; B = 8'h4F; #100;
A = 8'hC9; B = 8'h50; #100;
A = 8'hC9; B = 8'h51; #100;
A = 8'hC9; B = 8'h52; #100;
A = 8'hC9; B = 8'h53; #100;
A = 8'hC9; B = 8'h54; #100;
A = 8'hC9; B = 8'h55; #100;
A = 8'hC9; B = 8'h56; #100;
A = 8'hC9; B = 8'h57; #100;
A = 8'hC9; B = 8'h58; #100;
A = 8'hC9; B = 8'h59; #100;
A = 8'hC9; B = 8'h5A; #100;
A = 8'hC9; B = 8'h5B; #100;
A = 8'hC9; B = 8'h5C; #100;
A = 8'hC9; B = 8'h5D; #100;
A = 8'hC9; B = 8'h5E; #100;
A = 8'hC9; B = 8'h5F; #100;
A = 8'hC9; B = 8'h60; #100;
A = 8'hC9; B = 8'h61; #100;
A = 8'hC9; B = 8'h62; #100;
A = 8'hC9; B = 8'h63; #100;
A = 8'hC9; B = 8'h64; #100;
A = 8'hC9; B = 8'h65; #100;
A = 8'hC9; B = 8'h66; #100;
A = 8'hC9; B = 8'h67; #100;
A = 8'hC9; B = 8'h68; #100;
A = 8'hC9; B = 8'h69; #100;
A = 8'hC9; B = 8'h6A; #100;
A = 8'hC9; B = 8'h6B; #100;
A = 8'hC9; B = 8'h6C; #100;
A = 8'hC9; B = 8'h6D; #100;
A = 8'hC9; B = 8'h6E; #100;
A = 8'hC9; B = 8'h6F; #100;
A = 8'hC9; B = 8'h70; #100;
A = 8'hC9; B = 8'h71; #100;
A = 8'hC9; B = 8'h72; #100;
A = 8'hC9; B = 8'h73; #100;
A = 8'hC9; B = 8'h74; #100;
A = 8'hC9; B = 8'h75; #100;
A = 8'hC9; B = 8'h76; #100;
A = 8'hC9; B = 8'h77; #100;
A = 8'hC9; B = 8'h78; #100;
A = 8'hC9; B = 8'h79; #100;
A = 8'hC9; B = 8'h7A; #100;
A = 8'hC9; B = 8'h7B; #100;
A = 8'hC9; B = 8'h7C; #100;
A = 8'hC9; B = 8'h7D; #100;
A = 8'hC9; B = 8'h7E; #100;
A = 8'hC9; B = 8'h7F; #100;
A = 8'hC9; B = 8'h80; #100;
A = 8'hC9; B = 8'h81; #100;
A = 8'hC9; B = 8'h82; #100;
A = 8'hC9; B = 8'h83; #100;
A = 8'hC9; B = 8'h84; #100;
A = 8'hC9; B = 8'h85; #100;
A = 8'hC9; B = 8'h86; #100;
A = 8'hC9; B = 8'h87; #100;
A = 8'hC9; B = 8'h88; #100;
A = 8'hC9; B = 8'h89; #100;
A = 8'hC9; B = 8'h8A; #100;
A = 8'hC9; B = 8'h8B; #100;
A = 8'hC9; B = 8'h8C; #100;
A = 8'hC9; B = 8'h8D; #100;
A = 8'hC9; B = 8'h8E; #100;
A = 8'hC9; B = 8'h8F; #100;
A = 8'hC9; B = 8'h90; #100;
A = 8'hC9; B = 8'h91; #100;
A = 8'hC9; B = 8'h92; #100;
A = 8'hC9; B = 8'h93; #100;
A = 8'hC9; B = 8'h94; #100;
A = 8'hC9; B = 8'h95; #100;
A = 8'hC9; B = 8'h96; #100;
A = 8'hC9; B = 8'h97; #100;
A = 8'hC9; B = 8'h98; #100;
A = 8'hC9; B = 8'h99; #100;
A = 8'hC9; B = 8'h9A; #100;
A = 8'hC9; B = 8'h9B; #100;
A = 8'hC9; B = 8'h9C; #100;
A = 8'hC9; B = 8'h9D; #100;
A = 8'hC9; B = 8'h9E; #100;
A = 8'hC9; B = 8'h9F; #100;
A = 8'hC9; B = 8'hA0; #100;
A = 8'hC9; B = 8'hA1; #100;
A = 8'hC9; B = 8'hA2; #100;
A = 8'hC9; B = 8'hA3; #100;
A = 8'hC9; B = 8'hA4; #100;
A = 8'hC9; B = 8'hA5; #100;
A = 8'hC9; B = 8'hA6; #100;
A = 8'hC9; B = 8'hA7; #100;
A = 8'hC9; B = 8'hA8; #100;
A = 8'hC9; B = 8'hA9; #100;
A = 8'hC9; B = 8'hAA; #100;
A = 8'hC9; B = 8'hAB; #100;
A = 8'hC9; B = 8'hAC; #100;
A = 8'hC9; B = 8'hAD; #100;
A = 8'hC9; B = 8'hAE; #100;
A = 8'hC9; B = 8'hAF; #100;
A = 8'hC9; B = 8'hB0; #100;
A = 8'hC9; B = 8'hB1; #100;
A = 8'hC9; B = 8'hB2; #100;
A = 8'hC9; B = 8'hB3; #100;
A = 8'hC9; B = 8'hB4; #100;
A = 8'hC9; B = 8'hB5; #100;
A = 8'hC9; B = 8'hB6; #100;
A = 8'hC9; B = 8'hB7; #100;
A = 8'hC9; B = 8'hB8; #100;
A = 8'hC9; B = 8'hB9; #100;
A = 8'hC9; B = 8'hBA; #100;
A = 8'hC9; B = 8'hBB; #100;
A = 8'hC9; B = 8'hBC; #100;
A = 8'hC9; B = 8'hBD; #100;
A = 8'hC9; B = 8'hBE; #100;
A = 8'hC9; B = 8'hBF; #100;
A = 8'hC9; B = 8'hC0; #100;
A = 8'hC9; B = 8'hC1; #100;
A = 8'hC9; B = 8'hC2; #100;
A = 8'hC9; B = 8'hC3; #100;
A = 8'hC9; B = 8'hC4; #100;
A = 8'hC9; B = 8'hC5; #100;
A = 8'hC9; B = 8'hC6; #100;
A = 8'hC9; B = 8'hC7; #100;
A = 8'hC9; B = 8'hC8; #100;
A = 8'hC9; B = 8'hC9; #100;
A = 8'hC9; B = 8'hCA; #100;
A = 8'hC9; B = 8'hCB; #100;
A = 8'hC9; B = 8'hCC; #100;
A = 8'hC9; B = 8'hCD; #100;
A = 8'hC9; B = 8'hCE; #100;
A = 8'hC9; B = 8'hCF; #100;
A = 8'hC9; B = 8'hD0; #100;
A = 8'hC9; B = 8'hD1; #100;
A = 8'hC9; B = 8'hD2; #100;
A = 8'hC9; B = 8'hD3; #100;
A = 8'hC9; B = 8'hD4; #100;
A = 8'hC9; B = 8'hD5; #100;
A = 8'hC9; B = 8'hD6; #100;
A = 8'hC9; B = 8'hD7; #100;
A = 8'hC9; B = 8'hD8; #100;
A = 8'hC9; B = 8'hD9; #100;
A = 8'hC9; B = 8'hDA; #100;
A = 8'hC9; B = 8'hDB; #100;
A = 8'hC9; B = 8'hDC; #100;
A = 8'hC9; B = 8'hDD; #100;
A = 8'hC9; B = 8'hDE; #100;
A = 8'hC9; B = 8'hDF; #100;
A = 8'hC9; B = 8'hE0; #100;
A = 8'hC9; B = 8'hE1; #100;
A = 8'hC9; B = 8'hE2; #100;
A = 8'hC9; B = 8'hE3; #100;
A = 8'hC9; B = 8'hE4; #100;
A = 8'hC9; B = 8'hE5; #100;
A = 8'hC9; B = 8'hE6; #100;
A = 8'hC9; B = 8'hE7; #100;
A = 8'hC9; B = 8'hE8; #100;
A = 8'hC9; B = 8'hE9; #100;
A = 8'hC9; B = 8'hEA; #100;
A = 8'hC9; B = 8'hEB; #100;
A = 8'hC9; B = 8'hEC; #100;
A = 8'hC9; B = 8'hED; #100;
A = 8'hC9; B = 8'hEE; #100;
A = 8'hC9; B = 8'hEF; #100;
A = 8'hC9; B = 8'hF0; #100;
A = 8'hC9; B = 8'hF1; #100;
A = 8'hC9; B = 8'hF2; #100;
A = 8'hC9; B = 8'hF3; #100;
A = 8'hC9; B = 8'hF4; #100;
A = 8'hC9; B = 8'hF5; #100;
A = 8'hC9; B = 8'hF6; #100;
A = 8'hC9; B = 8'hF7; #100;
A = 8'hC9; B = 8'hF8; #100;
A = 8'hC9; B = 8'hF9; #100;
A = 8'hC9; B = 8'hFA; #100;
A = 8'hC9; B = 8'hFB; #100;
A = 8'hC9; B = 8'hFC; #100;
A = 8'hC9; B = 8'hFD; #100;
A = 8'hC9; B = 8'hFE; #100;
A = 8'hC9; B = 8'hFF; #100;
A = 8'hCA; B = 8'h0; #100;
A = 8'hCA; B = 8'h1; #100;
A = 8'hCA; B = 8'h2; #100;
A = 8'hCA; B = 8'h3; #100;
A = 8'hCA; B = 8'h4; #100;
A = 8'hCA; B = 8'h5; #100;
A = 8'hCA; B = 8'h6; #100;
A = 8'hCA; B = 8'h7; #100;
A = 8'hCA; B = 8'h8; #100;
A = 8'hCA; B = 8'h9; #100;
A = 8'hCA; B = 8'hA; #100;
A = 8'hCA; B = 8'hB; #100;
A = 8'hCA; B = 8'hC; #100;
A = 8'hCA; B = 8'hD; #100;
A = 8'hCA; B = 8'hE; #100;
A = 8'hCA; B = 8'hF; #100;
A = 8'hCA; B = 8'h10; #100;
A = 8'hCA; B = 8'h11; #100;
A = 8'hCA; B = 8'h12; #100;
A = 8'hCA; B = 8'h13; #100;
A = 8'hCA; B = 8'h14; #100;
A = 8'hCA; B = 8'h15; #100;
A = 8'hCA; B = 8'h16; #100;
A = 8'hCA; B = 8'h17; #100;
A = 8'hCA; B = 8'h18; #100;
A = 8'hCA; B = 8'h19; #100;
A = 8'hCA; B = 8'h1A; #100;
A = 8'hCA; B = 8'h1B; #100;
A = 8'hCA; B = 8'h1C; #100;
A = 8'hCA; B = 8'h1D; #100;
A = 8'hCA; B = 8'h1E; #100;
A = 8'hCA; B = 8'h1F; #100;
A = 8'hCA; B = 8'h20; #100;
A = 8'hCA; B = 8'h21; #100;
A = 8'hCA; B = 8'h22; #100;
A = 8'hCA; B = 8'h23; #100;
A = 8'hCA; B = 8'h24; #100;
A = 8'hCA; B = 8'h25; #100;
A = 8'hCA; B = 8'h26; #100;
A = 8'hCA; B = 8'h27; #100;
A = 8'hCA; B = 8'h28; #100;
A = 8'hCA; B = 8'h29; #100;
A = 8'hCA; B = 8'h2A; #100;
A = 8'hCA; B = 8'h2B; #100;
A = 8'hCA; B = 8'h2C; #100;
A = 8'hCA; B = 8'h2D; #100;
A = 8'hCA; B = 8'h2E; #100;
A = 8'hCA; B = 8'h2F; #100;
A = 8'hCA; B = 8'h30; #100;
A = 8'hCA; B = 8'h31; #100;
A = 8'hCA; B = 8'h32; #100;
A = 8'hCA; B = 8'h33; #100;
A = 8'hCA; B = 8'h34; #100;
A = 8'hCA; B = 8'h35; #100;
A = 8'hCA; B = 8'h36; #100;
A = 8'hCA; B = 8'h37; #100;
A = 8'hCA; B = 8'h38; #100;
A = 8'hCA; B = 8'h39; #100;
A = 8'hCA; B = 8'h3A; #100;
A = 8'hCA; B = 8'h3B; #100;
A = 8'hCA; B = 8'h3C; #100;
A = 8'hCA; B = 8'h3D; #100;
A = 8'hCA; B = 8'h3E; #100;
A = 8'hCA; B = 8'h3F; #100;
A = 8'hCA; B = 8'h40; #100;
A = 8'hCA; B = 8'h41; #100;
A = 8'hCA; B = 8'h42; #100;
A = 8'hCA; B = 8'h43; #100;
A = 8'hCA; B = 8'h44; #100;
A = 8'hCA; B = 8'h45; #100;
A = 8'hCA; B = 8'h46; #100;
A = 8'hCA; B = 8'h47; #100;
A = 8'hCA; B = 8'h48; #100;
A = 8'hCA; B = 8'h49; #100;
A = 8'hCA; B = 8'h4A; #100;
A = 8'hCA; B = 8'h4B; #100;
A = 8'hCA; B = 8'h4C; #100;
A = 8'hCA; B = 8'h4D; #100;
A = 8'hCA; B = 8'h4E; #100;
A = 8'hCA; B = 8'h4F; #100;
A = 8'hCA; B = 8'h50; #100;
A = 8'hCA; B = 8'h51; #100;
A = 8'hCA; B = 8'h52; #100;
A = 8'hCA; B = 8'h53; #100;
A = 8'hCA; B = 8'h54; #100;
A = 8'hCA; B = 8'h55; #100;
A = 8'hCA; B = 8'h56; #100;
A = 8'hCA; B = 8'h57; #100;
A = 8'hCA; B = 8'h58; #100;
A = 8'hCA; B = 8'h59; #100;
A = 8'hCA; B = 8'h5A; #100;
A = 8'hCA; B = 8'h5B; #100;
A = 8'hCA; B = 8'h5C; #100;
A = 8'hCA; B = 8'h5D; #100;
A = 8'hCA; B = 8'h5E; #100;
A = 8'hCA; B = 8'h5F; #100;
A = 8'hCA; B = 8'h60; #100;
A = 8'hCA; B = 8'h61; #100;
A = 8'hCA; B = 8'h62; #100;
A = 8'hCA; B = 8'h63; #100;
A = 8'hCA; B = 8'h64; #100;
A = 8'hCA; B = 8'h65; #100;
A = 8'hCA; B = 8'h66; #100;
A = 8'hCA; B = 8'h67; #100;
A = 8'hCA; B = 8'h68; #100;
A = 8'hCA; B = 8'h69; #100;
A = 8'hCA; B = 8'h6A; #100;
A = 8'hCA; B = 8'h6B; #100;
A = 8'hCA; B = 8'h6C; #100;
A = 8'hCA; B = 8'h6D; #100;
A = 8'hCA; B = 8'h6E; #100;
A = 8'hCA; B = 8'h6F; #100;
A = 8'hCA; B = 8'h70; #100;
A = 8'hCA; B = 8'h71; #100;
A = 8'hCA; B = 8'h72; #100;
A = 8'hCA; B = 8'h73; #100;
A = 8'hCA; B = 8'h74; #100;
A = 8'hCA; B = 8'h75; #100;
A = 8'hCA; B = 8'h76; #100;
A = 8'hCA; B = 8'h77; #100;
A = 8'hCA; B = 8'h78; #100;
A = 8'hCA; B = 8'h79; #100;
A = 8'hCA; B = 8'h7A; #100;
A = 8'hCA; B = 8'h7B; #100;
A = 8'hCA; B = 8'h7C; #100;
A = 8'hCA; B = 8'h7D; #100;
A = 8'hCA; B = 8'h7E; #100;
A = 8'hCA; B = 8'h7F; #100;
A = 8'hCA; B = 8'h80; #100;
A = 8'hCA; B = 8'h81; #100;
A = 8'hCA; B = 8'h82; #100;
A = 8'hCA; B = 8'h83; #100;
A = 8'hCA; B = 8'h84; #100;
A = 8'hCA; B = 8'h85; #100;
A = 8'hCA; B = 8'h86; #100;
A = 8'hCA; B = 8'h87; #100;
A = 8'hCA; B = 8'h88; #100;
A = 8'hCA; B = 8'h89; #100;
A = 8'hCA; B = 8'h8A; #100;
A = 8'hCA; B = 8'h8B; #100;
A = 8'hCA; B = 8'h8C; #100;
A = 8'hCA; B = 8'h8D; #100;
A = 8'hCA; B = 8'h8E; #100;
A = 8'hCA; B = 8'h8F; #100;
A = 8'hCA; B = 8'h90; #100;
A = 8'hCA; B = 8'h91; #100;
A = 8'hCA; B = 8'h92; #100;
A = 8'hCA; B = 8'h93; #100;
A = 8'hCA; B = 8'h94; #100;
A = 8'hCA; B = 8'h95; #100;
A = 8'hCA; B = 8'h96; #100;
A = 8'hCA; B = 8'h97; #100;
A = 8'hCA; B = 8'h98; #100;
A = 8'hCA; B = 8'h99; #100;
A = 8'hCA; B = 8'h9A; #100;
A = 8'hCA; B = 8'h9B; #100;
A = 8'hCA; B = 8'h9C; #100;
A = 8'hCA; B = 8'h9D; #100;
A = 8'hCA; B = 8'h9E; #100;
A = 8'hCA; B = 8'h9F; #100;
A = 8'hCA; B = 8'hA0; #100;
A = 8'hCA; B = 8'hA1; #100;
A = 8'hCA; B = 8'hA2; #100;
A = 8'hCA; B = 8'hA3; #100;
A = 8'hCA; B = 8'hA4; #100;
A = 8'hCA; B = 8'hA5; #100;
A = 8'hCA; B = 8'hA6; #100;
A = 8'hCA; B = 8'hA7; #100;
A = 8'hCA; B = 8'hA8; #100;
A = 8'hCA; B = 8'hA9; #100;
A = 8'hCA; B = 8'hAA; #100;
A = 8'hCA; B = 8'hAB; #100;
A = 8'hCA; B = 8'hAC; #100;
A = 8'hCA; B = 8'hAD; #100;
A = 8'hCA; B = 8'hAE; #100;
A = 8'hCA; B = 8'hAF; #100;
A = 8'hCA; B = 8'hB0; #100;
A = 8'hCA; B = 8'hB1; #100;
A = 8'hCA; B = 8'hB2; #100;
A = 8'hCA; B = 8'hB3; #100;
A = 8'hCA; B = 8'hB4; #100;
A = 8'hCA; B = 8'hB5; #100;
A = 8'hCA; B = 8'hB6; #100;
A = 8'hCA; B = 8'hB7; #100;
A = 8'hCA; B = 8'hB8; #100;
A = 8'hCA; B = 8'hB9; #100;
A = 8'hCA; B = 8'hBA; #100;
A = 8'hCA; B = 8'hBB; #100;
A = 8'hCA; B = 8'hBC; #100;
A = 8'hCA; B = 8'hBD; #100;
A = 8'hCA; B = 8'hBE; #100;
A = 8'hCA; B = 8'hBF; #100;
A = 8'hCA; B = 8'hC0; #100;
A = 8'hCA; B = 8'hC1; #100;
A = 8'hCA; B = 8'hC2; #100;
A = 8'hCA; B = 8'hC3; #100;
A = 8'hCA; B = 8'hC4; #100;
A = 8'hCA; B = 8'hC5; #100;
A = 8'hCA; B = 8'hC6; #100;
A = 8'hCA; B = 8'hC7; #100;
A = 8'hCA; B = 8'hC8; #100;
A = 8'hCA; B = 8'hC9; #100;
A = 8'hCA; B = 8'hCA; #100;
A = 8'hCA; B = 8'hCB; #100;
A = 8'hCA; B = 8'hCC; #100;
A = 8'hCA; B = 8'hCD; #100;
A = 8'hCA; B = 8'hCE; #100;
A = 8'hCA; B = 8'hCF; #100;
A = 8'hCA; B = 8'hD0; #100;
A = 8'hCA; B = 8'hD1; #100;
A = 8'hCA; B = 8'hD2; #100;
A = 8'hCA; B = 8'hD3; #100;
A = 8'hCA; B = 8'hD4; #100;
A = 8'hCA; B = 8'hD5; #100;
A = 8'hCA; B = 8'hD6; #100;
A = 8'hCA; B = 8'hD7; #100;
A = 8'hCA; B = 8'hD8; #100;
A = 8'hCA; B = 8'hD9; #100;
A = 8'hCA; B = 8'hDA; #100;
A = 8'hCA; B = 8'hDB; #100;
A = 8'hCA; B = 8'hDC; #100;
A = 8'hCA; B = 8'hDD; #100;
A = 8'hCA; B = 8'hDE; #100;
A = 8'hCA; B = 8'hDF; #100;
A = 8'hCA; B = 8'hE0; #100;
A = 8'hCA; B = 8'hE1; #100;
A = 8'hCA; B = 8'hE2; #100;
A = 8'hCA; B = 8'hE3; #100;
A = 8'hCA; B = 8'hE4; #100;
A = 8'hCA; B = 8'hE5; #100;
A = 8'hCA; B = 8'hE6; #100;
A = 8'hCA; B = 8'hE7; #100;
A = 8'hCA; B = 8'hE8; #100;
A = 8'hCA; B = 8'hE9; #100;
A = 8'hCA; B = 8'hEA; #100;
A = 8'hCA; B = 8'hEB; #100;
A = 8'hCA; B = 8'hEC; #100;
A = 8'hCA; B = 8'hED; #100;
A = 8'hCA; B = 8'hEE; #100;
A = 8'hCA; B = 8'hEF; #100;
A = 8'hCA; B = 8'hF0; #100;
A = 8'hCA; B = 8'hF1; #100;
A = 8'hCA; B = 8'hF2; #100;
A = 8'hCA; B = 8'hF3; #100;
A = 8'hCA; B = 8'hF4; #100;
A = 8'hCA; B = 8'hF5; #100;
A = 8'hCA; B = 8'hF6; #100;
A = 8'hCA; B = 8'hF7; #100;
A = 8'hCA; B = 8'hF8; #100;
A = 8'hCA; B = 8'hF9; #100;
A = 8'hCA; B = 8'hFA; #100;
A = 8'hCA; B = 8'hFB; #100;
A = 8'hCA; B = 8'hFC; #100;
A = 8'hCA; B = 8'hFD; #100;
A = 8'hCA; B = 8'hFE; #100;
A = 8'hCA; B = 8'hFF; #100;
A = 8'hCB; B = 8'h0; #100;
A = 8'hCB; B = 8'h1; #100;
A = 8'hCB; B = 8'h2; #100;
A = 8'hCB; B = 8'h3; #100;
A = 8'hCB; B = 8'h4; #100;
A = 8'hCB; B = 8'h5; #100;
A = 8'hCB; B = 8'h6; #100;
A = 8'hCB; B = 8'h7; #100;
A = 8'hCB; B = 8'h8; #100;
A = 8'hCB; B = 8'h9; #100;
A = 8'hCB; B = 8'hA; #100;
A = 8'hCB; B = 8'hB; #100;
A = 8'hCB; B = 8'hC; #100;
A = 8'hCB; B = 8'hD; #100;
A = 8'hCB; B = 8'hE; #100;
A = 8'hCB; B = 8'hF; #100;
A = 8'hCB; B = 8'h10; #100;
A = 8'hCB; B = 8'h11; #100;
A = 8'hCB; B = 8'h12; #100;
A = 8'hCB; B = 8'h13; #100;
A = 8'hCB; B = 8'h14; #100;
A = 8'hCB; B = 8'h15; #100;
A = 8'hCB; B = 8'h16; #100;
A = 8'hCB; B = 8'h17; #100;
A = 8'hCB; B = 8'h18; #100;
A = 8'hCB; B = 8'h19; #100;
A = 8'hCB; B = 8'h1A; #100;
A = 8'hCB; B = 8'h1B; #100;
A = 8'hCB; B = 8'h1C; #100;
A = 8'hCB; B = 8'h1D; #100;
A = 8'hCB; B = 8'h1E; #100;
A = 8'hCB; B = 8'h1F; #100;
A = 8'hCB; B = 8'h20; #100;
A = 8'hCB; B = 8'h21; #100;
A = 8'hCB; B = 8'h22; #100;
A = 8'hCB; B = 8'h23; #100;
A = 8'hCB; B = 8'h24; #100;
A = 8'hCB; B = 8'h25; #100;
A = 8'hCB; B = 8'h26; #100;
A = 8'hCB; B = 8'h27; #100;
A = 8'hCB; B = 8'h28; #100;
A = 8'hCB; B = 8'h29; #100;
A = 8'hCB; B = 8'h2A; #100;
A = 8'hCB; B = 8'h2B; #100;
A = 8'hCB; B = 8'h2C; #100;
A = 8'hCB; B = 8'h2D; #100;
A = 8'hCB; B = 8'h2E; #100;
A = 8'hCB; B = 8'h2F; #100;
A = 8'hCB; B = 8'h30; #100;
A = 8'hCB; B = 8'h31; #100;
A = 8'hCB; B = 8'h32; #100;
A = 8'hCB; B = 8'h33; #100;
A = 8'hCB; B = 8'h34; #100;
A = 8'hCB; B = 8'h35; #100;
A = 8'hCB; B = 8'h36; #100;
A = 8'hCB; B = 8'h37; #100;
A = 8'hCB; B = 8'h38; #100;
A = 8'hCB; B = 8'h39; #100;
A = 8'hCB; B = 8'h3A; #100;
A = 8'hCB; B = 8'h3B; #100;
A = 8'hCB; B = 8'h3C; #100;
A = 8'hCB; B = 8'h3D; #100;
A = 8'hCB; B = 8'h3E; #100;
A = 8'hCB; B = 8'h3F; #100;
A = 8'hCB; B = 8'h40; #100;
A = 8'hCB; B = 8'h41; #100;
A = 8'hCB; B = 8'h42; #100;
A = 8'hCB; B = 8'h43; #100;
A = 8'hCB; B = 8'h44; #100;
A = 8'hCB; B = 8'h45; #100;
A = 8'hCB; B = 8'h46; #100;
A = 8'hCB; B = 8'h47; #100;
A = 8'hCB; B = 8'h48; #100;
A = 8'hCB; B = 8'h49; #100;
A = 8'hCB; B = 8'h4A; #100;
A = 8'hCB; B = 8'h4B; #100;
A = 8'hCB; B = 8'h4C; #100;
A = 8'hCB; B = 8'h4D; #100;
A = 8'hCB; B = 8'h4E; #100;
A = 8'hCB; B = 8'h4F; #100;
A = 8'hCB; B = 8'h50; #100;
A = 8'hCB; B = 8'h51; #100;
A = 8'hCB; B = 8'h52; #100;
A = 8'hCB; B = 8'h53; #100;
A = 8'hCB; B = 8'h54; #100;
A = 8'hCB; B = 8'h55; #100;
A = 8'hCB; B = 8'h56; #100;
A = 8'hCB; B = 8'h57; #100;
A = 8'hCB; B = 8'h58; #100;
A = 8'hCB; B = 8'h59; #100;
A = 8'hCB; B = 8'h5A; #100;
A = 8'hCB; B = 8'h5B; #100;
A = 8'hCB; B = 8'h5C; #100;
A = 8'hCB; B = 8'h5D; #100;
A = 8'hCB; B = 8'h5E; #100;
A = 8'hCB; B = 8'h5F; #100;
A = 8'hCB; B = 8'h60; #100;
A = 8'hCB; B = 8'h61; #100;
A = 8'hCB; B = 8'h62; #100;
A = 8'hCB; B = 8'h63; #100;
A = 8'hCB; B = 8'h64; #100;
A = 8'hCB; B = 8'h65; #100;
A = 8'hCB; B = 8'h66; #100;
A = 8'hCB; B = 8'h67; #100;
A = 8'hCB; B = 8'h68; #100;
A = 8'hCB; B = 8'h69; #100;
A = 8'hCB; B = 8'h6A; #100;
A = 8'hCB; B = 8'h6B; #100;
A = 8'hCB; B = 8'h6C; #100;
A = 8'hCB; B = 8'h6D; #100;
A = 8'hCB; B = 8'h6E; #100;
A = 8'hCB; B = 8'h6F; #100;
A = 8'hCB; B = 8'h70; #100;
A = 8'hCB; B = 8'h71; #100;
A = 8'hCB; B = 8'h72; #100;
A = 8'hCB; B = 8'h73; #100;
A = 8'hCB; B = 8'h74; #100;
A = 8'hCB; B = 8'h75; #100;
A = 8'hCB; B = 8'h76; #100;
A = 8'hCB; B = 8'h77; #100;
A = 8'hCB; B = 8'h78; #100;
A = 8'hCB; B = 8'h79; #100;
A = 8'hCB; B = 8'h7A; #100;
A = 8'hCB; B = 8'h7B; #100;
A = 8'hCB; B = 8'h7C; #100;
A = 8'hCB; B = 8'h7D; #100;
A = 8'hCB; B = 8'h7E; #100;
A = 8'hCB; B = 8'h7F; #100;
A = 8'hCB; B = 8'h80; #100;
A = 8'hCB; B = 8'h81; #100;
A = 8'hCB; B = 8'h82; #100;
A = 8'hCB; B = 8'h83; #100;
A = 8'hCB; B = 8'h84; #100;
A = 8'hCB; B = 8'h85; #100;
A = 8'hCB; B = 8'h86; #100;
A = 8'hCB; B = 8'h87; #100;
A = 8'hCB; B = 8'h88; #100;
A = 8'hCB; B = 8'h89; #100;
A = 8'hCB; B = 8'h8A; #100;
A = 8'hCB; B = 8'h8B; #100;
A = 8'hCB; B = 8'h8C; #100;
A = 8'hCB; B = 8'h8D; #100;
A = 8'hCB; B = 8'h8E; #100;
A = 8'hCB; B = 8'h8F; #100;
A = 8'hCB; B = 8'h90; #100;
A = 8'hCB; B = 8'h91; #100;
A = 8'hCB; B = 8'h92; #100;
A = 8'hCB; B = 8'h93; #100;
A = 8'hCB; B = 8'h94; #100;
A = 8'hCB; B = 8'h95; #100;
A = 8'hCB; B = 8'h96; #100;
A = 8'hCB; B = 8'h97; #100;
A = 8'hCB; B = 8'h98; #100;
A = 8'hCB; B = 8'h99; #100;
A = 8'hCB; B = 8'h9A; #100;
A = 8'hCB; B = 8'h9B; #100;
A = 8'hCB; B = 8'h9C; #100;
A = 8'hCB; B = 8'h9D; #100;
A = 8'hCB; B = 8'h9E; #100;
A = 8'hCB; B = 8'h9F; #100;
A = 8'hCB; B = 8'hA0; #100;
A = 8'hCB; B = 8'hA1; #100;
A = 8'hCB; B = 8'hA2; #100;
A = 8'hCB; B = 8'hA3; #100;
A = 8'hCB; B = 8'hA4; #100;
A = 8'hCB; B = 8'hA5; #100;
A = 8'hCB; B = 8'hA6; #100;
A = 8'hCB; B = 8'hA7; #100;
A = 8'hCB; B = 8'hA8; #100;
A = 8'hCB; B = 8'hA9; #100;
A = 8'hCB; B = 8'hAA; #100;
A = 8'hCB; B = 8'hAB; #100;
A = 8'hCB; B = 8'hAC; #100;
A = 8'hCB; B = 8'hAD; #100;
A = 8'hCB; B = 8'hAE; #100;
A = 8'hCB; B = 8'hAF; #100;
A = 8'hCB; B = 8'hB0; #100;
A = 8'hCB; B = 8'hB1; #100;
A = 8'hCB; B = 8'hB2; #100;
A = 8'hCB; B = 8'hB3; #100;
A = 8'hCB; B = 8'hB4; #100;
A = 8'hCB; B = 8'hB5; #100;
A = 8'hCB; B = 8'hB6; #100;
A = 8'hCB; B = 8'hB7; #100;
A = 8'hCB; B = 8'hB8; #100;
A = 8'hCB; B = 8'hB9; #100;
A = 8'hCB; B = 8'hBA; #100;
A = 8'hCB; B = 8'hBB; #100;
A = 8'hCB; B = 8'hBC; #100;
A = 8'hCB; B = 8'hBD; #100;
A = 8'hCB; B = 8'hBE; #100;
A = 8'hCB; B = 8'hBF; #100;
A = 8'hCB; B = 8'hC0; #100;
A = 8'hCB; B = 8'hC1; #100;
A = 8'hCB; B = 8'hC2; #100;
A = 8'hCB; B = 8'hC3; #100;
A = 8'hCB; B = 8'hC4; #100;
A = 8'hCB; B = 8'hC5; #100;
A = 8'hCB; B = 8'hC6; #100;
A = 8'hCB; B = 8'hC7; #100;
A = 8'hCB; B = 8'hC8; #100;
A = 8'hCB; B = 8'hC9; #100;
A = 8'hCB; B = 8'hCA; #100;
A = 8'hCB; B = 8'hCB; #100;
A = 8'hCB; B = 8'hCC; #100;
A = 8'hCB; B = 8'hCD; #100;
A = 8'hCB; B = 8'hCE; #100;
A = 8'hCB; B = 8'hCF; #100;
A = 8'hCB; B = 8'hD0; #100;
A = 8'hCB; B = 8'hD1; #100;
A = 8'hCB; B = 8'hD2; #100;
A = 8'hCB; B = 8'hD3; #100;
A = 8'hCB; B = 8'hD4; #100;
A = 8'hCB; B = 8'hD5; #100;
A = 8'hCB; B = 8'hD6; #100;
A = 8'hCB; B = 8'hD7; #100;
A = 8'hCB; B = 8'hD8; #100;
A = 8'hCB; B = 8'hD9; #100;
A = 8'hCB; B = 8'hDA; #100;
A = 8'hCB; B = 8'hDB; #100;
A = 8'hCB; B = 8'hDC; #100;
A = 8'hCB; B = 8'hDD; #100;
A = 8'hCB; B = 8'hDE; #100;
A = 8'hCB; B = 8'hDF; #100;
A = 8'hCB; B = 8'hE0; #100;
A = 8'hCB; B = 8'hE1; #100;
A = 8'hCB; B = 8'hE2; #100;
A = 8'hCB; B = 8'hE3; #100;
A = 8'hCB; B = 8'hE4; #100;
A = 8'hCB; B = 8'hE5; #100;
A = 8'hCB; B = 8'hE6; #100;
A = 8'hCB; B = 8'hE7; #100;
A = 8'hCB; B = 8'hE8; #100;
A = 8'hCB; B = 8'hE9; #100;
A = 8'hCB; B = 8'hEA; #100;
A = 8'hCB; B = 8'hEB; #100;
A = 8'hCB; B = 8'hEC; #100;
A = 8'hCB; B = 8'hED; #100;
A = 8'hCB; B = 8'hEE; #100;
A = 8'hCB; B = 8'hEF; #100;
A = 8'hCB; B = 8'hF0; #100;
A = 8'hCB; B = 8'hF1; #100;
A = 8'hCB; B = 8'hF2; #100;
A = 8'hCB; B = 8'hF3; #100;
A = 8'hCB; B = 8'hF4; #100;
A = 8'hCB; B = 8'hF5; #100;
A = 8'hCB; B = 8'hF6; #100;
A = 8'hCB; B = 8'hF7; #100;
A = 8'hCB; B = 8'hF8; #100;
A = 8'hCB; B = 8'hF9; #100;
A = 8'hCB; B = 8'hFA; #100;
A = 8'hCB; B = 8'hFB; #100;
A = 8'hCB; B = 8'hFC; #100;
A = 8'hCB; B = 8'hFD; #100;
A = 8'hCB; B = 8'hFE; #100;
A = 8'hCB; B = 8'hFF; #100;
A = 8'hCC; B = 8'h0; #100;
A = 8'hCC; B = 8'h1; #100;
A = 8'hCC; B = 8'h2; #100;
A = 8'hCC; B = 8'h3; #100;
A = 8'hCC; B = 8'h4; #100;
A = 8'hCC; B = 8'h5; #100;
A = 8'hCC; B = 8'h6; #100;
A = 8'hCC; B = 8'h7; #100;
A = 8'hCC; B = 8'h8; #100;
A = 8'hCC; B = 8'h9; #100;
A = 8'hCC; B = 8'hA; #100;
A = 8'hCC; B = 8'hB; #100;
A = 8'hCC; B = 8'hC; #100;
A = 8'hCC; B = 8'hD; #100;
A = 8'hCC; B = 8'hE; #100;
A = 8'hCC; B = 8'hF; #100;
A = 8'hCC; B = 8'h10; #100;
A = 8'hCC; B = 8'h11; #100;
A = 8'hCC; B = 8'h12; #100;
A = 8'hCC; B = 8'h13; #100;
A = 8'hCC; B = 8'h14; #100;
A = 8'hCC; B = 8'h15; #100;
A = 8'hCC; B = 8'h16; #100;
A = 8'hCC; B = 8'h17; #100;
A = 8'hCC; B = 8'h18; #100;
A = 8'hCC; B = 8'h19; #100;
A = 8'hCC; B = 8'h1A; #100;
A = 8'hCC; B = 8'h1B; #100;
A = 8'hCC; B = 8'h1C; #100;
A = 8'hCC; B = 8'h1D; #100;
A = 8'hCC; B = 8'h1E; #100;
A = 8'hCC; B = 8'h1F; #100;
A = 8'hCC; B = 8'h20; #100;
A = 8'hCC; B = 8'h21; #100;
A = 8'hCC; B = 8'h22; #100;
A = 8'hCC; B = 8'h23; #100;
A = 8'hCC; B = 8'h24; #100;
A = 8'hCC; B = 8'h25; #100;
A = 8'hCC; B = 8'h26; #100;
A = 8'hCC; B = 8'h27; #100;
A = 8'hCC; B = 8'h28; #100;
A = 8'hCC; B = 8'h29; #100;
A = 8'hCC; B = 8'h2A; #100;
A = 8'hCC; B = 8'h2B; #100;
A = 8'hCC; B = 8'h2C; #100;
A = 8'hCC; B = 8'h2D; #100;
A = 8'hCC; B = 8'h2E; #100;
A = 8'hCC; B = 8'h2F; #100;
A = 8'hCC; B = 8'h30; #100;
A = 8'hCC; B = 8'h31; #100;
A = 8'hCC; B = 8'h32; #100;
A = 8'hCC; B = 8'h33; #100;
A = 8'hCC; B = 8'h34; #100;
A = 8'hCC; B = 8'h35; #100;
A = 8'hCC; B = 8'h36; #100;
A = 8'hCC; B = 8'h37; #100;
A = 8'hCC; B = 8'h38; #100;
A = 8'hCC; B = 8'h39; #100;
A = 8'hCC; B = 8'h3A; #100;
A = 8'hCC; B = 8'h3B; #100;
A = 8'hCC; B = 8'h3C; #100;
A = 8'hCC; B = 8'h3D; #100;
A = 8'hCC; B = 8'h3E; #100;
A = 8'hCC; B = 8'h3F; #100;
A = 8'hCC; B = 8'h40; #100;
A = 8'hCC; B = 8'h41; #100;
A = 8'hCC; B = 8'h42; #100;
A = 8'hCC; B = 8'h43; #100;
A = 8'hCC; B = 8'h44; #100;
A = 8'hCC; B = 8'h45; #100;
A = 8'hCC; B = 8'h46; #100;
A = 8'hCC; B = 8'h47; #100;
A = 8'hCC; B = 8'h48; #100;
A = 8'hCC; B = 8'h49; #100;
A = 8'hCC; B = 8'h4A; #100;
A = 8'hCC; B = 8'h4B; #100;
A = 8'hCC; B = 8'h4C; #100;
A = 8'hCC; B = 8'h4D; #100;
A = 8'hCC; B = 8'h4E; #100;
A = 8'hCC; B = 8'h4F; #100;
A = 8'hCC; B = 8'h50; #100;
A = 8'hCC; B = 8'h51; #100;
A = 8'hCC; B = 8'h52; #100;
A = 8'hCC; B = 8'h53; #100;
A = 8'hCC; B = 8'h54; #100;
A = 8'hCC; B = 8'h55; #100;
A = 8'hCC; B = 8'h56; #100;
A = 8'hCC; B = 8'h57; #100;
A = 8'hCC; B = 8'h58; #100;
A = 8'hCC; B = 8'h59; #100;
A = 8'hCC; B = 8'h5A; #100;
A = 8'hCC; B = 8'h5B; #100;
A = 8'hCC; B = 8'h5C; #100;
A = 8'hCC; B = 8'h5D; #100;
A = 8'hCC; B = 8'h5E; #100;
A = 8'hCC; B = 8'h5F; #100;
A = 8'hCC; B = 8'h60; #100;
A = 8'hCC; B = 8'h61; #100;
A = 8'hCC; B = 8'h62; #100;
A = 8'hCC; B = 8'h63; #100;
A = 8'hCC; B = 8'h64; #100;
A = 8'hCC; B = 8'h65; #100;
A = 8'hCC; B = 8'h66; #100;
A = 8'hCC; B = 8'h67; #100;
A = 8'hCC; B = 8'h68; #100;
A = 8'hCC; B = 8'h69; #100;
A = 8'hCC; B = 8'h6A; #100;
A = 8'hCC; B = 8'h6B; #100;
A = 8'hCC; B = 8'h6C; #100;
A = 8'hCC; B = 8'h6D; #100;
A = 8'hCC; B = 8'h6E; #100;
A = 8'hCC; B = 8'h6F; #100;
A = 8'hCC; B = 8'h70; #100;
A = 8'hCC; B = 8'h71; #100;
A = 8'hCC; B = 8'h72; #100;
A = 8'hCC; B = 8'h73; #100;
A = 8'hCC; B = 8'h74; #100;
A = 8'hCC; B = 8'h75; #100;
A = 8'hCC; B = 8'h76; #100;
A = 8'hCC; B = 8'h77; #100;
A = 8'hCC; B = 8'h78; #100;
A = 8'hCC; B = 8'h79; #100;
A = 8'hCC; B = 8'h7A; #100;
A = 8'hCC; B = 8'h7B; #100;
A = 8'hCC; B = 8'h7C; #100;
A = 8'hCC; B = 8'h7D; #100;
A = 8'hCC; B = 8'h7E; #100;
A = 8'hCC; B = 8'h7F; #100;
A = 8'hCC; B = 8'h80; #100;
A = 8'hCC; B = 8'h81; #100;
A = 8'hCC; B = 8'h82; #100;
A = 8'hCC; B = 8'h83; #100;
A = 8'hCC; B = 8'h84; #100;
A = 8'hCC; B = 8'h85; #100;
A = 8'hCC; B = 8'h86; #100;
A = 8'hCC; B = 8'h87; #100;
A = 8'hCC; B = 8'h88; #100;
A = 8'hCC; B = 8'h89; #100;
A = 8'hCC; B = 8'h8A; #100;
A = 8'hCC; B = 8'h8B; #100;
A = 8'hCC; B = 8'h8C; #100;
A = 8'hCC; B = 8'h8D; #100;
A = 8'hCC; B = 8'h8E; #100;
A = 8'hCC; B = 8'h8F; #100;
A = 8'hCC; B = 8'h90; #100;
A = 8'hCC; B = 8'h91; #100;
A = 8'hCC; B = 8'h92; #100;
A = 8'hCC; B = 8'h93; #100;
A = 8'hCC; B = 8'h94; #100;
A = 8'hCC; B = 8'h95; #100;
A = 8'hCC; B = 8'h96; #100;
A = 8'hCC; B = 8'h97; #100;
A = 8'hCC; B = 8'h98; #100;
A = 8'hCC; B = 8'h99; #100;
A = 8'hCC; B = 8'h9A; #100;
A = 8'hCC; B = 8'h9B; #100;
A = 8'hCC; B = 8'h9C; #100;
A = 8'hCC; B = 8'h9D; #100;
A = 8'hCC; B = 8'h9E; #100;
A = 8'hCC; B = 8'h9F; #100;
A = 8'hCC; B = 8'hA0; #100;
A = 8'hCC; B = 8'hA1; #100;
A = 8'hCC; B = 8'hA2; #100;
A = 8'hCC; B = 8'hA3; #100;
A = 8'hCC; B = 8'hA4; #100;
A = 8'hCC; B = 8'hA5; #100;
A = 8'hCC; B = 8'hA6; #100;
A = 8'hCC; B = 8'hA7; #100;
A = 8'hCC; B = 8'hA8; #100;
A = 8'hCC; B = 8'hA9; #100;
A = 8'hCC; B = 8'hAA; #100;
A = 8'hCC; B = 8'hAB; #100;
A = 8'hCC; B = 8'hAC; #100;
A = 8'hCC; B = 8'hAD; #100;
A = 8'hCC; B = 8'hAE; #100;
A = 8'hCC; B = 8'hAF; #100;
A = 8'hCC; B = 8'hB0; #100;
A = 8'hCC; B = 8'hB1; #100;
A = 8'hCC; B = 8'hB2; #100;
A = 8'hCC; B = 8'hB3; #100;
A = 8'hCC; B = 8'hB4; #100;
A = 8'hCC; B = 8'hB5; #100;
A = 8'hCC; B = 8'hB6; #100;
A = 8'hCC; B = 8'hB7; #100;
A = 8'hCC; B = 8'hB8; #100;
A = 8'hCC; B = 8'hB9; #100;
A = 8'hCC; B = 8'hBA; #100;
A = 8'hCC; B = 8'hBB; #100;
A = 8'hCC; B = 8'hBC; #100;
A = 8'hCC; B = 8'hBD; #100;
A = 8'hCC; B = 8'hBE; #100;
A = 8'hCC; B = 8'hBF; #100;
A = 8'hCC; B = 8'hC0; #100;
A = 8'hCC; B = 8'hC1; #100;
A = 8'hCC; B = 8'hC2; #100;
A = 8'hCC; B = 8'hC3; #100;
A = 8'hCC; B = 8'hC4; #100;
A = 8'hCC; B = 8'hC5; #100;
A = 8'hCC; B = 8'hC6; #100;
A = 8'hCC; B = 8'hC7; #100;
A = 8'hCC; B = 8'hC8; #100;
A = 8'hCC; B = 8'hC9; #100;
A = 8'hCC; B = 8'hCA; #100;
A = 8'hCC; B = 8'hCB; #100;
A = 8'hCC; B = 8'hCC; #100;
A = 8'hCC; B = 8'hCD; #100;
A = 8'hCC; B = 8'hCE; #100;
A = 8'hCC; B = 8'hCF; #100;
A = 8'hCC; B = 8'hD0; #100;
A = 8'hCC; B = 8'hD1; #100;
A = 8'hCC; B = 8'hD2; #100;
A = 8'hCC; B = 8'hD3; #100;
A = 8'hCC; B = 8'hD4; #100;
A = 8'hCC; B = 8'hD5; #100;
A = 8'hCC; B = 8'hD6; #100;
A = 8'hCC; B = 8'hD7; #100;
A = 8'hCC; B = 8'hD8; #100;
A = 8'hCC; B = 8'hD9; #100;
A = 8'hCC; B = 8'hDA; #100;
A = 8'hCC; B = 8'hDB; #100;
A = 8'hCC; B = 8'hDC; #100;
A = 8'hCC; B = 8'hDD; #100;
A = 8'hCC; B = 8'hDE; #100;
A = 8'hCC; B = 8'hDF; #100;
A = 8'hCC; B = 8'hE0; #100;
A = 8'hCC; B = 8'hE1; #100;
A = 8'hCC; B = 8'hE2; #100;
A = 8'hCC; B = 8'hE3; #100;
A = 8'hCC; B = 8'hE4; #100;
A = 8'hCC; B = 8'hE5; #100;
A = 8'hCC; B = 8'hE6; #100;
A = 8'hCC; B = 8'hE7; #100;
A = 8'hCC; B = 8'hE8; #100;
A = 8'hCC; B = 8'hE9; #100;
A = 8'hCC; B = 8'hEA; #100;
A = 8'hCC; B = 8'hEB; #100;
A = 8'hCC; B = 8'hEC; #100;
A = 8'hCC; B = 8'hED; #100;
A = 8'hCC; B = 8'hEE; #100;
A = 8'hCC; B = 8'hEF; #100;
A = 8'hCC; B = 8'hF0; #100;
A = 8'hCC; B = 8'hF1; #100;
A = 8'hCC; B = 8'hF2; #100;
A = 8'hCC; B = 8'hF3; #100;
A = 8'hCC; B = 8'hF4; #100;
A = 8'hCC; B = 8'hF5; #100;
A = 8'hCC; B = 8'hF6; #100;
A = 8'hCC; B = 8'hF7; #100;
A = 8'hCC; B = 8'hF8; #100;
A = 8'hCC; B = 8'hF9; #100;
A = 8'hCC; B = 8'hFA; #100;
A = 8'hCC; B = 8'hFB; #100;
A = 8'hCC; B = 8'hFC; #100;
A = 8'hCC; B = 8'hFD; #100;
A = 8'hCC; B = 8'hFE; #100;
A = 8'hCC; B = 8'hFF; #100;
A = 8'hCD; B = 8'h0; #100;
A = 8'hCD; B = 8'h1; #100;
A = 8'hCD; B = 8'h2; #100;
A = 8'hCD; B = 8'h3; #100;
A = 8'hCD; B = 8'h4; #100;
A = 8'hCD; B = 8'h5; #100;
A = 8'hCD; B = 8'h6; #100;
A = 8'hCD; B = 8'h7; #100;
A = 8'hCD; B = 8'h8; #100;
A = 8'hCD; B = 8'h9; #100;
A = 8'hCD; B = 8'hA; #100;
A = 8'hCD; B = 8'hB; #100;
A = 8'hCD; B = 8'hC; #100;
A = 8'hCD; B = 8'hD; #100;
A = 8'hCD; B = 8'hE; #100;
A = 8'hCD; B = 8'hF; #100;
A = 8'hCD; B = 8'h10; #100;
A = 8'hCD; B = 8'h11; #100;
A = 8'hCD; B = 8'h12; #100;
A = 8'hCD; B = 8'h13; #100;
A = 8'hCD; B = 8'h14; #100;
A = 8'hCD; B = 8'h15; #100;
A = 8'hCD; B = 8'h16; #100;
A = 8'hCD; B = 8'h17; #100;
A = 8'hCD; B = 8'h18; #100;
A = 8'hCD; B = 8'h19; #100;
A = 8'hCD; B = 8'h1A; #100;
A = 8'hCD; B = 8'h1B; #100;
A = 8'hCD; B = 8'h1C; #100;
A = 8'hCD; B = 8'h1D; #100;
A = 8'hCD; B = 8'h1E; #100;
A = 8'hCD; B = 8'h1F; #100;
A = 8'hCD; B = 8'h20; #100;
A = 8'hCD; B = 8'h21; #100;
A = 8'hCD; B = 8'h22; #100;
A = 8'hCD; B = 8'h23; #100;
A = 8'hCD; B = 8'h24; #100;
A = 8'hCD; B = 8'h25; #100;
A = 8'hCD; B = 8'h26; #100;
A = 8'hCD; B = 8'h27; #100;
A = 8'hCD; B = 8'h28; #100;
A = 8'hCD; B = 8'h29; #100;
A = 8'hCD; B = 8'h2A; #100;
A = 8'hCD; B = 8'h2B; #100;
A = 8'hCD; B = 8'h2C; #100;
A = 8'hCD; B = 8'h2D; #100;
A = 8'hCD; B = 8'h2E; #100;
A = 8'hCD; B = 8'h2F; #100;
A = 8'hCD; B = 8'h30; #100;
A = 8'hCD; B = 8'h31; #100;
A = 8'hCD; B = 8'h32; #100;
A = 8'hCD; B = 8'h33; #100;
A = 8'hCD; B = 8'h34; #100;
A = 8'hCD; B = 8'h35; #100;
A = 8'hCD; B = 8'h36; #100;
A = 8'hCD; B = 8'h37; #100;
A = 8'hCD; B = 8'h38; #100;
A = 8'hCD; B = 8'h39; #100;
A = 8'hCD; B = 8'h3A; #100;
A = 8'hCD; B = 8'h3B; #100;
A = 8'hCD; B = 8'h3C; #100;
A = 8'hCD; B = 8'h3D; #100;
A = 8'hCD; B = 8'h3E; #100;
A = 8'hCD; B = 8'h3F; #100;
A = 8'hCD; B = 8'h40; #100;
A = 8'hCD; B = 8'h41; #100;
A = 8'hCD; B = 8'h42; #100;
A = 8'hCD; B = 8'h43; #100;
A = 8'hCD; B = 8'h44; #100;
A = 8'hCD; B = 8'h45; #100;
A = 8'hCD; B = 8'h46; #100;
A = 8'hCD; B = 8'h47; #100;
A = 8'hCD; B = 8'h48; #100;
A = 8'hCD; B = 8'h49; #100;
A = 8'hCD; B = 8'h4A; #100;
A = 8'hCD; B = 8'h4B; #100;
A = 8'hCD; B = 8'h4C; #100;
A = 8'hCD; B = 8'h4D; #100;
A = 8'hCD; B = 8'h4E; #100;
A = 8'hCD; B = 8'h4F; #100;
A = 8'hCD; B = 8'h50; #100;
A = 8'hCD; B = 8'h51; #100;
A = 8'hCD; B = 8'h52; #100;
A = 8'hCD; B = 8'h53; #100;
A = 8'hCD; B = 8'h54; #100;
A = 8'hCD; B = 8'h55; #100;
A = 8'hCD; B = 8'h56; #100;
A = 8'hCD; B = 8'h57; #100;
A = 8'hCD; B = 8'h58; #100;
A = 8'hCD; B = 8'h59; #100;
A = 8'hCD; B = 8'h5A; #100;
A = 8'hCD; B = 8'h5B; #100;
A = 8'hCD; B = 8'h5C; #100;
A = 8'hCD; B = 8'h5D; #100;
A = 8'hCD; B = 8'h5E; #100;
A = 8'hCD; B = 8'h5F; #100;
A = 8'hCD; B = 8'h60; #100;
A = 8'hCD; B = 8'h61; #100;
A = 8'hCD; B = 8'h62; #100;
A = 8'hCD; B = 8'h63; #100;
A = 8'hCD; B = 8'h64; #100;
A = 8'hCD; B = 8'h65; #100;
A = 8'hCD; B = 8'h66; #100;
A = 8'hCD; B = 8'h67; #100;
A = 8'hCD; B = 8'h68; #100;
A = 8'hCD; B = 8'h69; #100;
A = 8'hCD; B = 8'h6A; #100;
A = 8'hCD; B = 8'h6B; #100;
A = 8'hCD; B = 8'h6C; #100;
A = 8'hCD; B = 8'h6D; #100;
A = 8'hCD; B = 8'h6E; #100;
A = 8'hCD; B = 8'h6F; #100;
A = 8'hCD; B = 8'h70; #100;
A = 8'hCD; B = 8'h71; #100;
A = 8'hCD; B = 8'h72; #100;
A = 8'hCD; B = 8'h73; #100;
A = 8'hCD; B = 8'h74; #100;
A = 8'hCD; B = 8'h75; #100;
A = 8'hCD; B = 8'h76; #100;
A = 8'hCD; B = 8'h77; #100;
A = 8'hCD; B = 8'h78; #100;
A = 8'hCD; B = 8'h79; #100;
A = 8'hCD; B = 8'h7A; #100;
A = 8'hCD; B = 8'h7B; #100;
A = 8'hCD; B = 8'h7C; #100;
A = 8'hCD; B = 8'h7D; #100;
A = 8'hCD; B = 8'h7E; #100;
A = 8'hCD; B = 8'h7F; #100;
A = 8'hCD; B = 8'h80; #100;
A = 8'hCD; B = 8'h81; #100;
A = 8'hCD; B = 8'h82; #100;
A = 8'hCD; B = 8'h83; #100;
A = 8'hCD; B = 8'h84; #100;
A = 8'hCD; B = 8'h85; #100;
A = 8'hCD; B = 8'h86; #100;
A = 8'hCD; B = 8'h87; #100;
A = 8'hCD; B = 8'h88; #100;
A = 8'hCD; B = 8'h89; #100;
A = 8'hCD; B = 8'h8A; #100;
A = 8'hCD; B = 8'h8B; #100;
A = 8'hCD; B = 8'h8C; #100;
A = 8'hCD; B = 8'h8D; #100;
A = 8'hCD; B = 8'h8E; #100;
A = 8'hCD; B = 8'h8F; #100;
A = 8'hCD; B = 8'h90; #100;
A = 8'hCD; B = 8'h91; #100;
A = 8'hCD; B = 8'h92; #100;
A = 8'hCD; B = 8'h93; #100;
A = 8'hCD; B = 8'h94; #100;
A = 8'hCD; B = 8'h95; #100;
A = 8'hCD; B = 8'h96; #100;
A = 8'hCD; B = 8'h97; #100;
A = 8'hCD; B = 8'h98; #100;
A = 8'hCD; B = 8'h99; #100;
A = 8'hCD; B = 8'h9A; #100;
A = 8'hCD; B = 8'h9B; #100;
A = 8'hCD; B = 8'h9C; #100;
A = 8'hCD; B = 8'h9D; #100;
A = 8'hCD; B = 8'h9E; #100;
A = 8'hCD; B = 8'h9F; #100;
A = 8'hCD; B = 8'hA0; #100;
A = 8'hCD; B = 8'hA1; #100;
A = 8'hCD; B = 8'hA2; #100;
A = 8'hCD; B = 8'hA3; #100;
A = 8'hCD; B = 8'hA4; #100;
A = 8'hCD; B = 8'hA5; #100;
A = 8'hCD; B = 8'hA6; #100;
A = 8'hCD; B = 8'hA7; #100;
A = 8'hCD; B = 8'hA8; #100;
A = 8'hCD; B = 8'hA9; #100;
A = 8'hCD; B = 8'hAA; #100;
A = 8'hCD; B = 8'hAB; #100;
A = 8'hCD; B = 8'hAC; #100;
A = 8'hCD; B = 8'hAD; #100;
A = 8'hCD; B = 8'hAE; #100;
A = 8'hCD; B = 8'hAF; #100;
A = 8'hCD; B = 8'hB0; #100;
A = 8'hCD; B = 8'hB1; #100;
A = 8'hCD; B = 8'hB2; #100;
A = 8'hCD; B = 8'hB3; #100;
A = 8'hCD; B = 8'hB4; #100;
A = 8'hCD; B = 8'hB5; #100;
A = 8'hCD; B = 8'hB6; #100;
A = 8'hCD; B = 8'hB7; #100;
A = 8'hCD; B = 8'hB8; #100;
A = 8'hCD; B = 8'hB9; #100;
A = 8'hCD; B = 8'hBA; #100;
A = 8'hCD; B = 8'hBB; #100;
A = 8'hCD; B = 8'hBC; #100;
A = 8'hCD; B = 8'hBD; #100;
A = 8'hCD; B = 8'hBE; #100;
A = 8'hCD; B = 8'hBF; #100;
A = 8'hCD; B = 8'hC0; #100;
A = 8'hCD; B = 8'hC1; #100;
A = 8'hCD; B = 8'hC2; #100;
A = 8'hCD; B = 8'hC3; #100;
A = 8'hCD; B = 8'hC4; #100;
A = 8'hCD; B = 8'hC5; #100;
A = 8'hCD; B = 8'hC6; #100;
A = 8'hCD; B = 8'hC7; #100;
A = 8'hCD; B = 8'hC8; #100;
A = 8'hCD; B = 8'hC9; #100;
A = 8'hCD; B = 8'hCA; #100;
A = 8'hCD; B = 8'hCB; #100;
A = 8'hCD; B = 8'hCC; #100;
A = 8'hCD; B = 8'hCD; #100;
A = 8'hCD; B = 8'hCE; #100;
A = 8'hCD; B = 8'hCF; #100;
A = 8'hCD; B = 8'hD0; #100;
A = 8'hCD; B = 8'hD1; #100;
A = 8'hCD; B = 8'hD2; #100;
A = 8'hCD; B = 8'hD3; #100;
A = 8'hCD; B = 8'hD4; #100;
A = 8'hCD; B = 8'hD5; #100;
A = 8'hCD; B = 8'hD6; #100;
A = 8'hCD; B = 8'hD7; #100;
A = 8'hCD; B = 8'hD8; #100;
A = 8'hCD; B = 8'hD9; #100;
A = 8'hCD; B = 8'hDA; #100;
A = 8'hCD; B = 8'hDB; #100;
A = 8'hCD; B = 8'hDC; #100;
A = 8'hCD; B = 8'hDD; #100;
A = 8'hCD; B = 8'hDE; #100;
A = 8'hCD; B = 8'hDF; #100;
A = 8'hCD; B = 8'hE0; #100;
A = 8'hCD; B = 8'hE1; #100;
A = 8'hCD; B = 8'hE2; #100;
A = 8'hCD; B = 8'hE3; #100;
A = 8'hCD; B = 8'hE4; #100;
A = 8'hCD; B = 8'hE5; #100;
A = 8'hCD; B = 8'hE6; #100;
A = 8'hCD; B = 8'hE7; #100;
A = 8'hCD; B = 8'hE8; #100;
A = 8'hCD; B = 8'hE9; #100;
A = 8'hCD; B = 8'hEA; #100;
A = 8'hCD; B = 8'hEB; #100;
A = 8'hCD; B = 8'hEC; #100;
A = 8'hCD; B = 8'hED; #100;
A = 8'hCD; B = 8'hEE; #100;
A = 8'hCD; B = 8'hEF; #100;
A = 8'hCD; B = 8'hF0; #100;
A = 8'hCD; B = 8'hF1; #100;
A = 8'hCD; B = 8'hF2; #100;
A = 8'hCD; B = 8'hF3; #100;
A = 8'hCD; B = 8'hF4; #100;
A = 8'hCD; B = 8'hF5; #100;
A = 8'hCD; B = 8'hF6; #100;
A = 8'hCD; B = 8'hF7; #100;
A = 8'hCD; B = 8'hF8; #100;
A = 8'hCD; B = 8'hF9; #100;
A = 8'hCD; B = 8'hFA; #100;
A = 8'hCD; B = 8'hFB; #100;
A = 8'hCD; B = 8'hFC; #100;
A = 8'hCD; B = 8'hFD; #100;
A = 8'hCD; B = 8'hFE; #100;
A = 8'hCD; B = 8'hFF; #100;
A = 8'hCE; B = 8'h0; #100;
A = 8'hCE; B = 8'h1; #100;
A = 8'hCE; B = 8'h2; #100;
A = 8'hCE; B = 8'h3; #100;
A = 8'hCE; B = 8'h4; #100;
A = 8'hCE; B = 8'h5; #100;
A = 8'hCE; B = 8'h6; #100;
A = 8'hCE; B = 8'h7; #100;
A = 8'hCE; B = 8'h8; #100;
A = 8'hCE; B = 8'h9; #100;
A = 8'hCE; B = 8'hA; #100;
A = 8'hCE; B = 8'hB; #100;
A = 8'hCE; B = 8'hC; #100;
A = 8'hCE; B = 8'hD; #100;
A = 8'hCE; B = 8'hE; #100;
A = 8'hCE; B = 8'hF; #100;
A = 8'hCE; B = 8'h10; #100;
A = 8'hCE; B = 8'h11; #100;
A = 8'hCE; B = 8'h12; #100;
A = 8'hCE; B = 8'h13; #100;
A = 8'hCE; B = 8'h14; #100;
A = 8'hCE; B = 8'h15; #100;
A = 8'hCE; B = 8'h16; #100;
A = 8'hCE; B = 8'h17; #100;
A = 8'hCE; B = 8'h18; #100;
A = 8'hCE; B = 8'h19; #100;
A = 8'hCE; B = 8'h1A; #100;
A = 8'hCE; B = 8'h1B; #100;
A = 8'hCE; B = 8'h1C; #100;
A = 8'hCE; B = 8'h1D; #100;
A = 8'hCE; B = 8'h1E; #100;
A = 8'hCE; B = 8'h1F; #100;
A = 8'hCE; B = 8'h20; #100;
A = 8'hCE; B = 8'h21; #100;
A = 8'hCE; B = 8'h22; #100;
A = 8'hCE; B = 8'h23; #100;
A = 8'hCE; B = 8'h24; #100;
A = 8'hCE; B = 8'h25; #100;
A = 8'hCE; B = 8'h26; #100;
A = 8'hCE; B = 8'h27; #100;
A = 8'hCE; B = 8'h28; #100;
A = 8'hCE; B = 8'h29; #100;
A = 8'hCE; B = 8'h2A; #100;
A = 8'hCE; B = 8'h2B; #100;
A = 8'hCE; B = 8'h2C; #100;
A = 8'hCE; B = 8'h2D; #100;
A = 8'hCE; B = 8'h2E; #100;
A = 8'hCE; B = 8'h2F; #100;
A = 8'hCE; B = 8'h30; #100;
A = 8'hCE; B = 8'h31; #100;
A = 8'hCE; B = 8'h32; #100;
A = 8'hCE; B = 8'h33; #100;
A = 8'hCE; B = 8'h34; #100;
A = 8'hCE; B = 8'h35; #100;
A = 8'hCE; B = 8'h36; #100;
A = 8'hCE; B = 8'h37; #100;
A = 8'hCE; B = 8'h38; #100;
A = 8'hCE; B = 8'h39; #100;
A = 8'hCE; B = 8'h3A; #100;
A = 8'hCE; B = 8'h3B; #100;
A = 8'hCE; B = 8'h3C; #100;
A = 8'hCE; B = 8'h3D; #100;
A = 8'hCE; B = 8'h3E; #100;
A = 8'hCE; B = 8'h3F; #100;
A = 8'hCE; B = 8'h40; #100;
A = 8'hCE; B = 8'h41; #100;
A = 8'hCE; B = 8'h42; #100;
A = 8'hCE; B = 8'h43; #100;
A = 8'hCE; B = 8'h44; #100;
A = 8'hCE; B = 8'h45; #100;
A = 8'hCE; B = 8'h46; #100;
A = 8'hCE; B = 8'h47; #100;
A = 8'hCE; B = 8'h48; #100;
A = 8'hCE; B = 8'h49; #100;
A = 8'hCE; B = 8'h4A; #100;
A = 8'hCE; B = 8'h4B; #100;
A = 8'hCE; B = 8'h4C; #100;
A = 8'hCE; B = 8'h4D; #100;
A = 8'hCE; B = 8'h4E; #100;
A = 8'hCE; B = 8'h4F; #100;
A = 8'hCE; B = 8'h50; #100;
A = 8'hCE; B = 8'h51; #100;
A = 8'hCE; B = 8'h52; #100;
A = 8'hCE; B = 8'h53; #100;
A = 8'hCE; B = 8'h54; #100;
A = 8'hCE; B = 8'h55; #100;
A = 8'hCE; B = 8'h56; #100;
A = 8'hCE; B = 8'h57; #100;
A = 8'hCE; B = 8'h58; #100;
A = 8'hCE; B = 8'h59; #100;
A = 8'hCE; B = 8'h5A; #100;
A = 8'hCE; B = 8'h5B; #100;
A = 8'hCE; B = 8'h5C; #100;
A = 8'hCE; B = 8'h5D; #100;
A = 8'hCE; B = 8'h5E; #100;
A = 8'hCE; B = 8'h5F; #100;
A = 8'hCE; B = 8'h60; #100;
A = 8'hCE; B = 8'h61; #100;
A = 8'hCE; B = 8'h62; #100;
A = 8'hCE; B = 8'h63; #100;
A = 8'hCE; B = 8'h64; #100;
A = 8'hCE; B = 8'h65; #100;
A = 8'hCE; B = 8'h66; #100;
A = 8'hCE; B = 8'h67; #100;
A = 8'hCE; B = 8'h68; #100;
A = 8'hCE; B = 8'h69; #100;
A = 8'hCE; B = 8'h6A; #100;
A = 8'hCE; B = 8'h6B; #100;
A = 8'hCE; B = 8'h6C; #100;
A = 8'hCE; B = 8'h6D; #100;
A = 8'hCE; B = 8'h6E; #100;
A = 8'hCE; B = 8'h6F; #100;
A = 8'hCE; B = 8'h70; #100;
A = 8'hCE; B = 8'h71; #100;
A = 8'hCE; B = 8'h72; #100;
A = 8'hCE; B = 8'h73; #100;
A = 8'hCE; B = 8'h74; #100;
A = 8'hCE; B = 8'h75; #100;
A = 8'hCE; B = 8'h76; #100;
A = 8'hCE; B = 8'h77; #100;
A = 8'hCE; B = 8'h78; #100;
A = 8'hCE; B = 8'h79; #100;
A = 8'hCE; B = 8'h7A; #100;
A = 8'hCE; B = 8'h7B; #100;
A = 8'hCE; B = 8'h7C; #100;
A = 8'hCE; B = 8'h7D; #100;
A = 8'hCE; B = 8'h7E; #100;
A = 8'hCE; B = 8'h7F; #100;
A = 8'hCE; B = 8'h80; #100;
A = 8'hCE; B = 8'h81; #100;
A = 8'hCE; B = 8'h82; #100;
A = 8'hCE; B = 8'h83; #100;
A = 8'hCE; B = 8'h84; #100;
A = 8'hCE; B = 8'h85; #100;
A = 8'hCE; B = 8'h86; #100;
A = 8'hCE; B = 8'h87; #100;
A = 8'hCE; B = 8'h88; #100;
A = 8'hCE; B = 8'h89; #100;
A = 8'hCE; B = 8'h8A; #100;
A = 8'hCE; B = 8'h8B; #100;
A = 8'hCE; B = 8'h8C; #100;
A = 8'hCE; B = 8'h8D; #100;
A = 8'hCE; B = 8'h8E; #100;
A = 8'hCE; B = 8'h8F; #100;
A = 8'hCE; B = 8'h90; #100;
A = 8'hCE; B = 8'h91; #100;
A = 8'hCE; B = 8'h92; #100;
A = 8'hCE; B = 8'h93; #100;
A = 8'hCE; B = 8'h94; #100;
A = 8'hCE; B = 8'h95; #100;
A = 8'hCE; B = 8'h96; #100;
A = 8'hCE; B = 8'h97; #100;
A = 8'hCE; B = 8'h98; #100;
A = 8'hCE; B = 8'h99; #100;
A = 8'hCE; B = 8'h9A; #100;
A = 8'hCE; B = 8'h9B; #100;
A = 8'hCE; B = 8'h9C; #100;
A = 8'hCE; B = 8'h9D; #100;
A = 8'hCE; B = 8'h9E; #100;
A = 8'hCE; B = 8'h9F; #100;
A = 8'hCE; B = 8'hA0; #100;
A = 8'hCE; B = 8'hA1; #100;
A = 8'hCE; B = 8'hA2; #100;
A = 8'hCE; B = 8'hA3; #100;
A = 8'hCE; B = 8'hA4; #100;
A = 8'hCE; B = 8'hA5; #100;
A = 8'hCE; B = 8'hA6; #100;
A = 8'hCE; B = 8'hA7; #100;
A = 8'hCE; B = 8'hA8; #100;
A = 8'hCE; B = 8'hA9; #100;
A = 8'hCE; B = 8'hAA; #100;
A = 8'hCE; B = 8'hAB; #100;
A = 8'hCE; B = 8'hAC; #100;
A = 8'hCE; B = 8'hAD; #100;
A = 8'hCE; B = 8'hAE; #100;
A = 8'hCE; B = 8'hAF; #100;
A = 8'hCE; B = 8'hB0; #100;
A = 8'hCE; B = 8'hB1; #100;
A = 8'hCE; B = 8'hB2; #100;
A = 8'hCE; B = 8'hB3; #100;
A = 8'hCE; B = 8'hB4; #100;
A = 8'hCE; B = 8'hB5; #100;
A = 8'hCE; B = 8'hB6; #100;
A = 8'hCE; B = 8'hB7; #100;
A = 8'hCE; B = 8'hB8; #100;
A = 8'hCE; B = 8'hB9; #100;
A = 8'hCE; B = 8'hBA; #100;
A = 8'hCE; B = 8'hBB; #100;
A = 8'hCE; B = 8'hBC; #100;
A = 8'hCE; B = 8'hBD; #100;
A = 8'hCE; B = 8'hBE; #100;
A = 8'hCE; B = 8'hBF; #100;
A = 8'hCE; B = 8'hC0; #100;
A = 8'hCE; B = 8'hC1; #100;
A = 8'hCE; B = 8'hC2; #100;
A = 8'hCE; B = 8'hC3; #100;
A = 8'hCE; B = 8'hC4; #100;
A = 8'hCE; B = 8'hC5; #100;
A = 8'hCE; B = 8'hC6; #100;
A = 8'hCE; B = 8'hC7; #100;
A = 8'hCE; B = 8'hC8; #100;
A = 8'hCE; B = 8'hC9; #100;
A = 8'hCE; B = 8'hCA; #100;
A = 8'hCE; B = 8'hCB; #100;
A = 8'hCE; B = 8'hCC; #100;
A = 8'hCE; B = 8'hCD; #100;
A = 8'hCE; B = 8'hCE; #100;
A = 8'hCE; B = 8'hCF; #100;
A = 8'hCE; B = 8'hD0; #100;
A = 8'hCE; B = 8'hD1; #100;
A = 8'hCE; B = 8'hD2; #100;
A = 8'hCE; B = 8'hD3; #100;
A = 8'hCE; B = 8'hD4; #100;
A = 8'hCE; B = 8'hD5; #100;
A = 8'hCE; B = 8'hD6; #100;
A = 8'hCE; B = 8'hD7; #100;
A = 8'hCE; B = 8'hD8; #100;
A = 8'hCE; B = 8'hD9; #100;
A = 8'hCE; B = 8'hDA; #100;
A = 8'hCE; B = 8'hDB; #100;
A = 8'hCE; B = 8'hDC; #100;
A = 8'hCE; B = 8'hDD; #100;
A = 8'hCE; B = 8'hDE; #100;
A = 8'hCE; B = 8'hDF; #100;
A = 8'hCE; B = 8'hE0; #100;
A = 8'hCE; B = 8'hE1; #100;
A = 8'hCE; B = 8'hE2; #100;
A = 8'hCE; B = 8'hE3; #100;
A = 8'hCE; B = 8'hE4; #100;
A = 8'hCE; B = 8'hE5; #100;
A = 8'hCE; B = 8'hE6; #100;
A = 8'hCE; B = 8'hE7; #100;
A = 8'hCE; B = 8'hE8; #100;
A = 8'hCE; B = 8'hE9; #100;
A = 8'hCE; B = 8'hEA; #100;
A = 8'hCE; B = 8'hEB; #100;
A = 8'hCE; B = 8'hEC; #100;
A = 8'hCE; B = 8'hED; #100;
A = 8'hCE; B = 8'hEE; #100;
A = 8'hCE; B = 8'hEF; #100;
A = 8'hCE; B = 8'hF0; #100;
A = 8'hCE; B = 8'hF1; #100;
A = 8'hCE; B = 8'hF2; #100;
A = 8'hCE; B = 8'hF3; #100;
A = 8'hCE; B = 8'hF4; #100;
A = 8'hCE; B = 8'hF5; #100;
A = 8'hCE; B = 8'hF6; #100;
A = 8'hCE; B = 8'hF7; #100;
A = 8'hCE; B = 8'hF8; #100;
A = 8'hCE; B = 8'hF9; #100;
A = 8'hCE; B = 8'hFA; #100;
A = 8'hCE; B = 8'hFB; #100;
A = 8'hCE; B = 8'hFC; #100;
A = 8'hCE; B = 8'hFD; #100;
A = 8'hCE; B = 8'hFE; #100;
A = 8'hCE; B = 8'hFF; #100;
A = 8'hCF; B = 8'h0; #100;
A = 8'hCF; B = 8'h1; #100;
A = 8'hCF; B = 8'h2; #100;
A = 8'hCF; B = 8'h3; #100;
A = 8'hCF; B = 8'h4; #100;
A = 8'hCF; B = 8'h5; #100;
A = 8'hCF; B = 8'h6; #100;
A = 8'hCF; B = 8'h7; #100;
A = 8'hCF; B = 8'h8; #100;
A = 8'hCF; B = 8'h9; #100;
A = 8'hCF; B = 8'hA; #100;
A = 8'hCF; B = 8'hB; #100;
A = 8'hCF; B = 8'hC; #100;
A = 8'hCF; B = 8'hD; #100;
A = 8'hCF; B = 8'hE; #100;
A = 8'hCF; B = 8'hF; #100;
A = 8'hCF; B = 8'h10; #100;
A = 8'hCF; B = 8'h11; #100;
A = 8'hCF; B = 8'h12; #100;
A = 8'hCF; B = 8'h13; #100;
A = 8'hCF; B = 8'h14; #100;
A = 8'hCF; B = 8'h15; #100;
A = 8'hCF; B = 8'h16; #100;
A = 8'hCF; B = 8'h17; #100;
A = 8'hCF; B = 8'h18; #100;
A = 8'hCF; B = 8'h19; #100;
A = 8'hCF; B = 8'h1A; #100;
A = 8'hCF; B = 8'h1B; #100;
A = 8'hCF; B = 8'h1C; #100;
A = 8'hCF; B = 8'h1D; #100;
A = 8'hCF; B = 8'h1E; #100;
A = 8'hCF; B = 8'h1F; #100;
A = 8'hCF; B = 8'h20; #100;
A = 8'hCF; B = 8'h21; #100;
A = 8'hCF; B = 8'h22; #100;
A = 8'hCF; B = 8'h23; #100;
A = 8'hCF; B = 8'h24; #100;
A = 8'hCF; B = 8'h25; #100;
A = 8'hCF; B = 8'h26; #100;
A = 8'hCF; B = 8'h27; #100;
A = 8'hCF; B = 8'h28; #100;
A = 8'hCF; B = 8'h29; #100;
A = 8'hCF; B = 8'h2A; #100;
A = 8'hCF; B = 8'h2B; #100;
A = 8'hCF; B = 8'h2C; #100;
A = 8'hCF; B = 8'h2D; #100;
A = 8'hCF; B = 8'h2E; #100;
A = 8'hCF; B = 8'h2F; #100;
A = 8'hCF; B = 8'h30; #100;
A = 8'hCF; B = 8'h31; #100;
A = 8'hCF; B = 8'h32; #100;
A = 8'hCF; B = 8'h33; #100;
A = 8'hCF; B = 8'h34; #100;
A = 8'hCF; B = 8'h35; #100;
A = 8'hCF; B = 8'h36; #100;
A = 8'hCF; B = 8'h37; #100;
A = 8'hCF; B = 8'h38; #100;
A = 8'hCF; B = 8'h39; #100;
A = 8'hCF; B = 8'h3A; #100;
A = 8'hCF; B = 8'h3B; #100;
A = 8'hCF; B = 8'h3C; #100;
A = 8'hCF; B = 8'h3D; #100;
A = 8'hCF; B = 8'h3E; #100;
A = 8'hCF; B = 8'h3F; #100;
A = 8'hCF; B = 8'h40; #100;
A = 8'hCF; B = 8'h41; #100;
A = 8'hCF; B = 8'h42; #100;
A = 8'hCF; B = 8'h43; #100;
A = 8'hCF; B = 8'h44; #100;
A = 8'hCF; B = 8'h45; #100;
A = 8'hCF; B = 8'h46; #100;
A = 8'hCF; B = 8'h47; #100;
A = 8'hCF; B = 8'h48; #100;
A = 8'hCF; B = 8'h49; #100;
A = 8'hCF; B = 8'h4A; #100;
A = 8'hCF; B = 8'h4B; #100;
A = 8'hCF; B = 8'h4C; #100;
A = 8'hCF; B = 8'h4D; #100;
A = 8'hCF; B = 8'h4E; #100;
A = 8'hCF; B = 8'h4F; #100;
A = 8'hCF; B = 8'h50; #100;
A = 8'hCF; B = 8'h51; #100;
A = 8'hCF; B = 8'h52; #100;
A = 8'hCF; B = 8'h53; #100;
A = 8'hCF; B = 8'h54; #100;
A = 8'hCF; B = 8'h55; #100;
A = 8'hCF; B = 8'h56; #100;
A = 8'hCF; B = 8'h57; #100;
A = 8'hCF; B = 8'h58; #100;
A = 8'hCF; B = 8'h59; #100;
A = 8'hCF; B = 8'h5A; #100;
A = 8'hCF; B = 8'h5B; #100;
A = 8'hCF; B = 8'h5C; #100;
A = 8'hCF; B = 8'h5D; #100;
A = 8'hCF; B = 8'h5E; #100;
A = 8'hCF; B = 8'h5F; #100;
A = 8'hCF; B = 8'h60; #100;
A = 8'hCF; B = 8'h61; #100;
A = 8'hCF; B = 8'h62; #100;
A = 8'hCF; B = 8'h63; #100;
A = 8'hCF; B = 8'h64; #100;
A = 8'hCF; B = 8'h65; #100;
A = 8'hCF; B = 8'h66; #100;
A = 8'hCF; B = 8'h67; #100;
A = 8'hCF; B = 8'h68; #100;
A = 8'hCF; B = 8'h69; #100;
A = 8'hCF; B = 8'h6A; #100;
A = 8'hCF; B = 8'h6B; #100;
A = 8'hCF; B = 8'h6C; #100;
A = 8'hCF; B = 8'h6D; #100;
A = 8'hCF; B = 8'h6E; #100;
A = 8'hCF; B = 8'h6F; #100;
A = 8'hCF; B = 8'h70; #100;
A = 8'hCF; B = 8'h71; #100;
A = 8'hCF; B = 8'h72; #100;
A = 8'hCF; B = 8'h73; #100;
A = 8'hCF; B = 8'h74; #100;
A = 8'hCF; B = 8'h75; #100;
A = 8'hCF; B = 8'h76; #100;
A = 8'hCF; B = 8'h77; #100;
A = 8'hCF; B = 8'h78; #100;
A = 8'hCF; B = 8'h79; #100;
A = 8'hCF; B = 8'h7A; #100;
A = 8'hCF; B = 8'h7B; #100;
A = 8'hCF; B = 8'h7C; #100;
A = 8'hCF; B = 8'h7D; #100;
A = 8'hCF; B = 8'h7E; #100;
A = 8'hCF; B = 8'h7F; #100;
A = 8'hCF; B = 8'h80; #100;
A = 8'hCF; B = 8'h81; #100;
A = 8'hCF; B = 8'h82; #100;
A = 8'hCF; B = 8'h83; #100;
A = 8'hCF; B = 8'h84; #100;
A = 8'hCF; B = 8'h85; #100;
A = 8'hCF; B = 8'h86; #100;
A = 8'hCF; B = 8'h87; #100;
A = 8'hCF; B = 8'h88; #100;
A = 8'hCF; B = 8'h89; #100;
A = 8'hCF; B = 8'h8A; #100;
A = 8'hCF; B = 8'h8B; #100;
A = 8'hCF; B = 8'h8C; #100;
A = 8'hCF; B = 8'h8D; #100;
A = 8'hCF; B = 8'h8E; #100;
A = 8'hCF; B = 8'h8F; #100;
A = 8'hCF; B = 8'h90; #100;
A = 8'hCF; B = 8'h91; #100;
A = 8'hCF; B = 8'h92; #100;
A = 8'hCF; B = 8'h93; #100;
A = 8'hCF; B = 8'h94; #100;
A = 8'hCF; B = 8'h95; #100;
A = 8'hCF; B = 8'h96; #100;
A = 8'hCF; B = 8'h97; #100;
A = 8'hCF; B = 8'h98; #100;
A = 8'hCF; B = 8'h99; #100;
A = 8'hCF; B = 8'h9A; #100;
A = 8'hCF; B = 8'h9B; #100;
A = 8'hCF; B = 8'h9C; #100;
A = 8'hCF; B = 8'h9D; #100;
A = 8'hCF; B = 8'h9E; #100;
A = 8'hCF; B = 8'h9F; #100;
A = 8'hCF; B = 8'hA0; #100;
A = 8'hCF; B = 8'hA1; #100;
A = 8'hCF; B = 8'hA2; #100;
A = 8'hCF; B = 8'hA3; #100;
A = 8'hCF; B = 8'hA4; #100;
A = 8'hCF; B = 8'hA5; #100;
A = 8'hCF; B = 8'hA6; #100;
A = 8'hCF; B = 8'hA7; #100;
A = 8'hCF; B = 8'hA8; #100;
A = 8'hCF; B = 8'hA9; #100;
A = 8'hCF; B = 8'hAA; #100;
A = 8'hCF; B = 8'hAB; #100;
A = 8'hCF; B = 8'hAC; #100;
A = 8'hCF; B = 8'hAD; #100;
A = 8'hCF; B = 8'hAE; #100;
A = 8'hCF; B = 8'hAF; #100;
A = 8'hCF; B = 8'hB0; #100;
A = 8'hCF; B = 8'hB1; #100;
A = 8'hCF; B = 8'hB2; #100;
A = 8'hCF; B = 8'hB3; #100;
A = 8'hCF; B = 8'hB4; #100;
A = 8'hCF; B = 8'hB5; #100;
A = 8'hCF; B = 8'hB6; #100;
A = 8'hCF; B = 8'hB7; #100;
A = 8'hCF; B = 8'hB8; #100;
A = 8'hCF; B = 8'hB9; #100;
A = 8'hCF; B = 8'hBA; #100;
A = 8'hCF; B = 8'hBB; #100;
A = 8'hCF; B = 8'hBC; #100;
A = 8'hCF; B = 8'hBD; #100;
A = 8'hCF; B = 8'hBE; #100;
A = 8'hCF; B = 8'hBF; #100;
A = 8'hCF; B = 8'hC0; #100;
A = 8'hCF; B = 8'hC1; #100;
A = 8'hCF; B = 8'hC2; #100;
A = 8'hCF; B = 8'hC3; #100;
A = 8'hCF; B = 8'hC4; #100;
A = 8'hCF; B = 8'hC5; #100;
A = 8'hCF; B = 8'hC6; #100;
A = 8'hCF; B = 8'hC7; #100;
A = 8'hCF; B = 8'hC8; #100;
A = 8'hCF; B = 8'hC9; #100;
A = 8'hCF; B = 8'hCA; #100;
A = 8'hCF; B = 8'hCB; #100;
A = 8'hCF; B = 8'hCC; #100;
A = 8'hCF; B = 8'hCD; #100;
A = 8'hCF; B = 8'hCE; #100;
A = 8'hCF; B = 8'hCF; #100;
A = 8'hCF; B = 8'hD0; #100;
A = 8'hCF; B = 8'hD1; #100;
A = 8'hCF; B = 8'hD2; #100;
A = 8'hCF; B = 8'hD3; #100;
A = 8'hCF; B = 8'hD4; #100;
A = 8'hCF; B = 8'hD5; #100;
A = 8'hCF; B = 8'hD6; #100;
A = 8'hCF; B = 8'hD7; #100;
A = 8'hCF; B = 8'hD8; #100;
A = 8'hCF; B = 8'hD9; #100;
A = 8'hCF; B = 8'hDA; #100;
A = 8'hCF; B = 8'hDB; #100;
A = 8'hCF; B = 8'hDC; #100;
A = 8'hCF; B = 8'hDD; #100;
A = 8'hCF; B = 8'hDE; #100;
A = 8'hCF; B = 8'hDF; #100;
A = 8'hCF; B = 8'hE0; #100;
A = 8'hCF; B = 8'hE1; #100;
A = 8'hCF; B = 8'hE2; #100;
A = 8'hCF; B = 8'hE3; #100;
A = 8'hCF; B = 8'hE4; #100;
A = 8'hCF; B = 8'hE5; #100;
A = 8'hCF; B = 8'hE6; #100;
A = 8'hCF; B = 8'hE7; #100;
A = 8'hCF; B = 8'hE8; #100;
A = 8'hCF; B = 8'hE9; #100;
A = 8'hCF; B = 8'hEA; #100;
A = 8'hCF; B = 8'hEB; #100;
A = 8'hCF; B = 8'hEC; #100;
A = 8'hCF; B = 8'hED; #100;
A = 8'hCF; B = 8'hEE; #100;
A = 8'hCF; B = 8'hEF; #100;
A = 8'hCF; B = 8'hF0; #100;
A = 8'hCF; B = 8'hF1; #100;
A = 8'hCF; B = 8'hF2; #100;
A = 8'hCF; B = 8'hF3; #100;
A = 8'hCF; B = 8'hF4; #100;
A = 8'hCF; B = 8'hF5; #100;
A = 8'hCF; B = 8'hF6; #100;
A = 8'hCF; B = 8'hF7; #100;
A = 8'hCF; B = 8'hF8; #100;
A = 8'hCF; B = 8'hF9; #100;
A = 8'hCF; B = 8'hFA; #100;
A = 8'hCF; B = 8'hFB; #100;
A = 8'hCF; B = 8'hFC; #100;
A = 8'hCF; B = 8'hFD; #100;
A = 8'hCF; B = 8'hFE; #100;
A = 8'hCF; B = 8'hFF; #100;
A = 8'hD0; B = 8'h0; #100;
A = 8'hD0; B = 8'h1; #100;
A = 8'hD0; B = 8'h2; #100;
A = 8'hD0; B = 8'h3; #100;
A = 8'hD0; B = 8'h4; #100;
A = 8'hD0; B = 8'h5; #100;
A = 8'hD0; B = 8'h6; #100;
A = 8'hD0; B = 8'h7; #100;
A = 8'hD0; B = 8'h8; #100;
A = 8'hD0; B = 8'h9; #100;
A = 8'hD0; B = 8'hA; #100;
A = 8'hD0; B = 8'hB; #100;
A = 8'hD0; B = 8'hC; #100;
A = 8'hD0; B = 8'hD; #100;
A = 8'hD0; B = 8'hE; #100;
A = 8'hD0; B = 8'hF; #100;
A = 8'hD0; B = 8'h10; #100;
A = 8'hD0; B = 8'h11; #100;
A = 8'hD0; B = 8'h12; #100;
A = 8'hD0; B = 8'h13; #100;
A = 8'hD0; B = 8'h14; #100;
A = 8'hD0; B = 8'h15; #100;
A = 8'hD0; B = 8'h16; #100;
A = 8'hD0; B = 8'h17; #100;
A = 8'hD0; B = 8'h18; #100;
A = 8'hD0; B = 8'h19; #100;
A = 8'hD0; B = 8'h1A; #100;
A = 8'hD0; B = 8'h1B; #100;
A = 8'hD0; B = 8'h1C; #100;
A = 8'hD0; B = 8'h1D; #100;
A = 8'hD0; B = 8'h1E; #100;
A = 8'hD0; B = 8'h1F; #100;
A = 8'hD0; B = 8'h20; #100;
A = 8'hD0; B = 8'h21; #100;
A = 8'hD0; B = 8'h22; #100;
A = 8'hD0; B = 8'h23; #100;
A = 8'hD0; B = 8'h24; #100;
A = 8'hD0; B = 8'h25; #100;
A = 8'hD0; B = 8'h26; #100;
A = 8'hD0; B = 8'h27; #100;
A = 8'hD0; B = 8'h28; #100;
A = 8'hD0; B = 8'h29; #100;
A = 8'hD0; B = 8'h2A; #100;
A = 8'hD0; B = 8'h2B; #100;
A = 8'hD0; B = 8'h2C; #100;
A = 8'hD0; B = 8'h2D; #100;
A = 8'hD0; B = 8'h2E; #100;
A = 8'hD0; B = 8'h2F; #100;
A = 8'hD0; B = 8'h30; #100;
A = 8'hD0; B = 8'h31; #100;
A = 8'hD0; B = 8'h32; #100;
A = 8'hD0; B = 8'h33; #100;
A = 8'hD0; B = 8'h34; #100;
A = 8'hD0; B = 8'h35; #100;
A = 8'hD0; B = 8'h36; #100;
A = 8'hD0; B = 8'h37; #100;
A = 8'hD0; B = 8'h38; #100;
A = 8'hD0; B = 8'h39; #100;
A = 8'hD0; B = 8'h3A; #100;
A = 8'hD0; B = 8'h3B; #100;
A = 8'hD0; B = 8'h3C; #100;
A = 8'hD0; B = 8'h3D; #100;
A = 8'hD0; B = 8'h3E; #100;
A = 8'hD0; B = 8'h3F; #100;
A = 8'hD0; B = 8'h40; #100;
A = 8'hD0; B = 8'h41; #100;
A = 8'hD0; B = 8'h42; #100;
A = 8'hD0; B = 8'h43; #100;
A = 8'hD0; B = 8'h44; #100;
A = 8'hD0; B = 8'h45; #100;
A = 8'hD0; B = 8'h46; #100;
A = 8'hD0; B = 8'h47; #100;
A = 8'hD0; B = 8'h48; #100;
A = 8'hD0; B = 8'h49; #100;
A = 8'hD0; B = 8'h4A; #100;
A = 8'hD0; B = 8'h4B; #100;
A = 8'hD0; B = 8'h4C; #100;
A = 8'hD0; B = 8'h4D; #100;
A = 8'hD0; B = 8'h4E; #100;
A = 8'hD0; B = 8'h4F; #100;
A = 8'hD0; B = 8'h50; #100;
A = 8'hD0; B = 8'h51; #100;
A = 8'hD0; B = 8'h52; #100;
A = 8'hD0; B = 8'h53; #100;
A = 8'hD0; B = 8'h54; #100;
A = 8'hD0; B = 8'h55; #100;
A = 8'hD0; B = 8'h56; #100;
A = 8'hD0; B = 8'h57; #100;
A = 8'hD0; B = 8'h58; #100;
A = 8'hD0; B = 8'h59; #100;
A = 8'hD0; B = 8'h5A; #100;
A = 8'hD0; B = 8'h5B; #100;
A = 8'hD0; B = 8'h5C; #100;
A = 8'hD0; B = 8'h5D; #100;
A = 8'hD0; B = 8'h5E; #100;
A = 8'hD0; B = 8'h5F; #100;
A = 8'hD0; B = 8'h60; #100;
A = 8'hD0; B = 8'h61; #100;
A = 8'hD0; B = 8'h62; #100;
A = 8'hD0; B = 8'h63; #100;
A = 8'hD0; B = 8'h64; #100;
A = 8'hD0; B = 8'h65; #100;
A = 8'hD0; B = 8'h66; #100;
A = 8'hD0; B = 8'h67; #100;
A = 8'hD0; B = 8'h68; #100;
A = 8'hD0; B = 8'h69; #100;
A = 8'hD0; B = 8'h6A; #100;
A = 8'hD0; B = 8'h6B; #100;
A = 8'hD0; B = 8'h6C; #100;
A = 8'hD0; B = 8'h6D; #100;
A = 8'hD0; B = 8'h6E; #100;
A = 8'hD0; B = 8'h6F; #100;
A = 8'hD0; B = 8'h70; #100;
A = 8'hD0; B = 8'h71; #100;
A = 8'hD0; B = 8'h72; #100;
A = 8'hD0; B = 8'h73; #100;
A = 8'hD0; B = 8'h74; #100;
A = 8'hD0; B = 8'h75; #100;
A = 8'hD0; B = 8'h76; #100;
A = 8'hD0; B = 8'h77; #100;
A = 8'hD0; B = 8'h78; #100;
A = 8'hD0; B = 8'h79; #100;
A = 8'hD0; B = 8'h7A; #100;
A = 8'hD0; B = 8'h7B; #100;
A = 8'hD0; B = 8'h7C; #100;
A = 8'hD0; B = 8'h7D; #100;
A = 8'hD0; B = 8'h7E; #100;
A = 8'hD0; B = 8'h7F; #100;
A = 8'hD0; B = 8'h80; #100;
A = 8'hD0; B = 8'h81; #100;
A = 8'hD0; B = 8'h82; #100;
A = 8'hD0; B = 8'h83; #100;
A = 8'hD0; B = 8'h84; #100;
A = 8'hD0; B = 8'h85; #100;
A = 8'hD0; B = 8'h86; #100;
A = 8'hD0; B = 8'h87; #100;
A = 8'hD0; B = 8'h88; #100;
A = 8'hD0; B = 8'h89; #100;
A = 8'hD0; B = 8'h8A; #100;
A = 8'hD0; B = 8'h8B; #100;
A = 8'hD0; B = 8'h8C; #100;
A = 8'hD0; B = 8'h8D; #100;
A = 8'hD0; B = 8'h8E; #100;
A = 8'hD0; B = 8'h8F; #100;
A = 8'hD0; B = 8'h90; #100;
A = 8'hD0; B = 8'h91; #100;
A = 8'hD0; B = 8'h92; #100;
A = 8'hD0; B = 8'h93; #100;
A = 8'hD0; B = 8'h94; #100;
A = 8'hD0; B = 8'h95; #100;
A = 8'hD0; B = 8'h96; #100;
A = 8'hD0; B = 8'h97; #100;
A = 8'hD0; B = 8'h98; #100;
A = 8'hD0; B = 8'h99; #100;
A = 8'hD0; B = 8'h9A; #100;
A = 8'hD0; B = 8'h9B; #100;
A = 8'hD0; B = 8'h9C; #100;
A = 8'hD0; B = 8'h9D; #100;
A = 8'hD0; B = 8'h9E; #100;
A = 8'hD0; B = 8'h9F; #100;
A = 8'hD0; B = 8'hA0; #100;
A = 8'hD0; B = 8'hA1; #100;
A = 8'hD0; B = 8'hA2; #100;
A = 8'hD0; B = 8'hA3; #100;
A = 8'hD0; B = 8'hA4; #100;
A = 8'hD0; B = 8'hA5; #100;
A = 8'hD0; B = 8'hA6; #100;
A = 8'hD0; B = 8'hA7; #100;
A = 8'hD0; B = 8'hA8; #100;
A = 8'hD0; B = 8'hA9; #100;
A = 8'hD0; B = 8'hAA; #100;
A = 8'hD0; B = 8'hAB; #100;
A = 8'hD0; B = 8'hAC; #100;
A = 8'hD0; B = 8'hAD; #100;
A = 8'hD0; B = 8'hAE; #100;
A = 8'hD0; B = 8'hAF; #100;
A = 8'hD0; B = 8'hB0; #100;
A = 8'hD0; B = 8'hB1; #100;
A = 8'hD0; B = 8'hB2; #100;
A = 8'hD0; B = 8'hB3; #100;
A = 8'hD0; B = 8'hB4; #100;
A = 8'hD0; B = 8'hB5; #100;
A = 8'hD0; B = 8'hB6; #100;
A = 8'hD0; B = 8'hB7; #100;
A = 8'hD0; B = 8'hB8; #100;
A = 8'hD0; B = 8'hB9; #100;
A = 8'hD0; B = 8'hBA; #100;
A = 8'hD0; B = 8'hBB; #100;
A = 8'hD0; B = 8'hBC; #100;
A = 8'hD0; B = 8'hBD; #100;
A = 8'hD0; B = 8'hBE; #100;
A = 8'hD0; B = 8'hBF; #100;
A = 8'hD0; B = 8'hC0; #100;
A = 8'hD0; B = 8'hC1; #100;
A = 8'hD0; B = 8'hC2; #100;
A = 8'hD0; B = 8'hC3; #100;
A = 8'hD0; B = 8'hC4; #100;
A = 8'hD0; B = 8'hC5; #100;
A = 8'hD0; B = 8'hC6; #100;
A = 8'hD0; B = 8'hC7; #100;
A = 8'hD0; B = 8'hC8; #100;
A = 8'hD0; B = 8'hC9; #100;
A = 8'hD0; B = 8'hCA; #100;
A = 8'hD0; B = 8'hCB; #100;
A = 8'hD0; B = 8'hCC; #100;
A = 8'hD0; B = 8'hCD; #100;
A = 8'hD0; B = 8'hCE; #100;
A = 8'hD0; B = 8'hCF; #100;
A = 8'hD0; B = 8'hD0; #100;
A = 8'hD0; B = 8'hD1; #100;
A = 8'hD0; B = 8'hD2; #100;
A = 8'hD0; B = 8'hD3; #100;
A = 8'hD0; B = 8'hD4; #100;
A = 8'hD0; B = 8'hD5; #100;
A = 8'hD0; B = 8'hD6; #100;
A = 8'hD0; B = 8'hD7; #100;
A = 8'hD0; B = 8'hD8; #100;
A = 8'hD0; B = 8'hD9; #100;
A = 8'hD0; B = 8'hDA; #100;
A = 8'hD0; B = 8'hDB; #100;
A = 8'hD0; B = 8'hDC; #100;
A = 8'hD0; B = 8'hDD; #100;
A = 8'hD0; B = 8'hDE; #100;
A = 8'hD0; B = 8'hDF; #100;
A = 8'hD0; B = 8'hE0; #100;
A = 8'hD0; B = 8'hE1; #100;
A = 8'hD0; B = 8'hE2; #100;
A = 8'hD0; B = 8'hE3; #100;
A = 8'hD0; B = 8'hE4; #100;
A = 8'hD0; B = 8'hE5; #100;
A = 8'hD0; B = 8'hE6; #100;
A = 8'hD0; B = 8'hE7; #100;
A = 8'hD0; B = 8'hE8; #100;
A = 8'hD0; B = 8'hE9; #100;
A = 8'hD0; B = 8'hEA; #100;
A = 8'hD0; B = 8'hEB; #100;
A = 8'hD0; B = 8'hEC; #100;
A = 8'hD0; B = 8'hED; #100;
A = 8'hD0; B = 8'hEE; #100;
A = 8'hD0; B = 8'hEF; #100;
A = 8'hD0; B = 8'hF0; #100;
A = 8'hD0; B = 8'hF1; #100;
A = 8'hD0; B = 8'hF2; #100;
A = 8'hD0; B = 8'hF3; #100;
A = 8'hD0; B = 8'hF4; #100;
A = 8'hD0; B = 8'hF5; #100;
A = 8'hD0; B = 8'hF6; #100;
A = 8'hD0; B = 8'hF7; #100;
A = 8'hD0; B = 8'hF8; #100;
A = 8'hD0; B = 8'hF9; #100;
A = 8'hD0; B = 8'hFA; #100;
A = 8'hD0; B = 8'hFB; #100;
A = 8'hD0; B = 8'hFC; #100;
A = 8'hD0; B = 8'hFD; #100;
A = 8'hD0; B = 8'hFE; #100;
A = 8'hD0; B = 8'hFF; #100;
A = 8'hD1; B = 8'h0; #100;
A = 8'hD1; B = 8'h1; #100;
A = 8'hD1; B = 8'h2; #100;
A = 8'hD1; B = 8'h3; #100;
A = 8'hD1; B = 8'h4; #100;
A = 8'hD1; B = 8'h5; #100;
A = 8'hD1; B = 8'h6; #100;
A = 8'hD1; B = 8'h7; #100;
A = 8'hD1; B = 8'h8; #100;
A = 8'hD1; B = 8'h9; #100;
A = 8'hD1; B = 8'hA; #100;
A = 8'hD1; B = 8'hB; #100;
A = 8'hD1; B = 8'hC; #100;
A = 8'hD1; B = 8'hD; #100;
A = 8'hD1; B = 8'hE; #100;
A = 8'hD1; B = 8'hF; #100;
A = 8'hD1; B = 8'h10; #100;
A = 8'hD1; B = 8'h11; #100;
A = 8'hD1; B = 8'h12; #100;
A = 8'hD1; B = 8'h13; #100;
A = 8'hD1; B = 8'h14; #100;
A = 8'hD1; B = 8'h15; #100;
A = 8'hD1; B = 8'h16; #100;
A = 8'hD1; B = 8'h17; #100;
A = 8'hD1; B = 8'h18; #100;
A = 8'hD1; B = 8'h19; #100;
A = 8'hD1; B = 8'h1A; #100;
A = 8'hD1; B = 8'h1B; #100;
A = 8'hD1; B = 8'h1C; #100;
A = 8'hD1; B = 8'h1D; #100;
A = 8'hD1; B = 8'h1E; #100;
A = 8'hD1; B = 8'h1F; #100;
A = 8'hD1; B = 8'h20; #100;
A = 8'hD1; B = 8'h21; #100;
A = 8'hD1; B = 8'h22; #100;
A = 8'hD1; B = 8'h23; #100;
A = 8'hD1; B = 8'h24; #100;
A = 8'hD1; B = 8'h25; #100;
A = 8'hD1; B = 8'h26; #100;
A = 8'hD1; B = 8'h27; #100;
A = 8'hD1; B = 8'h28; #100;
A = 8'hD1; B = 8'h29; #100;
A = 8'hD1; B = 8'h2A; #100;
A = 8'hD1; B = 8'h2B; #100;
A = 8'hD1; B = 8'h2C; #100;
A = 8'hD1; B = 8'h2D; #100;
A = 8'hD1; B = 8'h2E; #100;
A = 8'hD1; B = 8'h2F; #100;
A = 8'hD1; B = 8'h30; #100;
A = 8'hD1; B = 8'h31; #100;
A = 8'hD1; B = 8'h32; #100;
A = 8'hD1; B = 8'h33; #100;
A = 8'hD1; B = 8'h34; #100;
A = 8'hD1; B = 8'h35; #100;
A = 8'hD1; B = 8'h36; #100;
A = 8'hD1; B = 8'h37; #100;
A = 8'hD1; B = 8'h38; #100;
A = 8'hD1; B = 8'h39; #100;
A = 8'hD1; B = 8'h3A; #100;
A = 8'hD1; B = 8'h3B; #100;
A = 8'hD1; B = 8'h3C; #100;
A = 8'hD1; B = 8'h3D; #100;
A = 8'hD1; B = 8'h3E; #100;
A = 8'hD1; B = 8'h3F; #100;
A = 8'hD1; B = 8'h40; #100;
A = 8'hD1; B = 8'h41; #100;
A = 8'hD1; B = 8'h42; #100;
A = 8'hD1; B = 8'h43; #100;
A = 8'hD1; B = 8'h44; #100;
A = 8'hD1; B = 8'h45; #100;
A = 8'hD1; B = 8'h46; #100;
A = 8'hD1; B = 8'h47; #100;
A = 8'hD1; B = 8'h48; #100;
A = 8'hD1; B = 8'h49; #100;
A = 8'hD1; B = 8'h4A; #100;
A = 8'hD1; B = 8'h4B; #100;
A = 8'hD1; B = 8'h4C; #100;
A = 8'hD1; B = 8'h4D; #100;
A = 8'hD1; B = 8'h4E; #100;
A = 8'hD1; B = 8'h4F; #100;
A = 8'hD1; B = 8'h50; #100;
A = 8'hD1; B = 8'h51; #100;
A = 8'hD1; B = 8'h52; #100;
A = 8'hD1; B = 8'h53; #100;
A = 8'hD1; B = 8'h54; #100;
A = 8'hD1; B = 8'h55; #100;
A = 8'hD1; B = 8'h56; #100;
A = 8'hD1; B = 8'h57; #100;
A = 8'hD1; B = 8'h58; #100;
A = 8'hD1; B = 8'h59; #100;
A = 8'hD1; B = 8'h5A; #100;
A = 8'hD1; B = 8'h5B; #100;
A = 8'hD1; B = 8'h5C; #100;
A = 8'hD1; B = 8'h5D; #100;
A = 8'hD1; B = 8'h5E; #100;
A = 8'hD1; B = 8'h5F; #100;
A = 8'hD1; B = 8'h60; #100;
A = 8'hD1; B = 8'h61; #100;
A = 8'hD1; B = 8'h62; #100;
A = 8'hD1; B = 8'h63; #100;
A = 8'hD1; B = 8'h64; #100;
A = 8'hD1; B = 8'h65; #100;
A = 8'hD1; B = 8'h66; #100;
A = 8'hD1; B = 8'h67; #100;
A = 8'hD1; B = 8'h68; #100;
A = 8'hD1; B = 8'h69; #100;
A = 8'hD1; B = 8'h6A; #100;
A = 8'hD1; B = 8'h6B; #100;
A = 8'hD1; B = 8'h6C; #100;
A = 8'hD1; B = 8'h6D; #100;
A = 8'hD1; B = 8'h6E; #100;
A = 8'hD1; B = 8'h6F; #100;
A = 8'hD1; B = 8'h70; #100;
A = 8'hD1; B = 8'h71; #100;
A = 8'hD1; B = 8'h72; #100;
A = 8'hD1; B = 8'h73; #100;
A = 8'hD1; B = 8'h74; #100;
A = 8'hD1; B = 8'h75; #100;
A = 8'hD1; B = 8'h76; #100;
A = 8'hD1; B = 8'h77; #100;
A = 8'hD1; B = 8'h78; #100;
A = 8'hD1; B = 8'h79; #100;
A = 8'hD1; B = 8'h7A; #100;
A = 8'hD1; B = 8'h7B; #100;
A = 8'hD1; B = 8'h7C; #100;
A = 8'hD1; B = 8'h7D; #100;
A = 8'hD1; B = 8'h7E; #100;
A = 8'hD1; B = 8'h7F; #100;
A = 8'hD1; B = 8'h80; #100;
A = 8'hD1; B = 8'h81; #100;
A = 8'hD1; B = 8'h82; #100;
A = 8'hD1; B = 8'h83; #100;
A = 8'hD1; B = 8'h84; #100;
A = 8'hD1; B = 8'h85; #100;
A = 8'hD1; B = 8'h86; #100;
A = 8'hD1; B = 8'h87; #100;
A = 8'hD1; B = 8'h88; #100;
A = 8'hD1; B = 8'h89; #100;
A = 8'hD1; B = 8'h8A; #100;
A = 8'hD1; B = 8'h8B; #100;
A = 8'hD1; B = 8'h8C; #100;
A = 8'hD1; B = 8'h8D; #100;
A = 8'hD1; B = 8'h8E; #100;
A = 8'hD1; B = 8'h8F; #100;
A = 8'hD1; B = 8'h90; #100;
A = 8'hD1; B = 8'h91; #100;
A = 8'hD1; B = 8'h92; #100;
A = 8'hD1; B = 8'h93; #100;
A = 8'hD1; B = 8'h94; #100;
A = 8'hD1; B = 8'h95; #100;
A = 8'hD1; B = 8'h96; #100;
A = 8'hD1; B = 8'h97; #100;
A = 8'hD1; B = 8'h98; #100;
A = 8'hD1; B = 8'h99; #100;
A = 8'hD1; B = 8'h9A; #100;
A = 8'hD1; B = 8'h9B; #100;
A = 8'hD1; B = 8'h9C; #100;
A = 8'hD1; B = 8'h9D; #100;
A = 8'hD1; B = 8'h9E; #100;
A = 8'hD1; B = 8'h9F; #100;
A = 8'hD1; B = 8'hA0; #100;
A = 8'hD1; B = 8'hA1; #100;
A = 8'hD1; B = 8'hA2; #100;
A = 8'hD1; B = 8'hA3; #100;
A = 8'hD1; B = 8'hA4; #100;
A = 8'hD1; B = 8'hA5; #100;
A = 8'hD1; B = 8'hA6; #100;
A = 8'hD1; B = 8'hA7; #100;
A = 8'hD1; B = 8'hA8; #100;
A = 8'hD1; B = 8'hA9; #100;
A = 8'hD1; B = 8'hAA; #100;
A = 8'hD1; B = 8'hAB; #100;
A = 8'hD1; B = 8'hAC; #100;
A = 8'hD1; B = 8'hAD; #100;
A = 8'hD1; B = 8'hAE; #100;
A = 8'hD1; B = 8'hAF; #100;
A = 8'hD1; B = 8'hB0; #100;
A = 8'hD1; B = 8'hB1; #100;
A = 8'hD1; B = 8'hB2; #100;
A = 8'hD1; B = 8'hB3; #100;
A = 8'hD1; B = 8'hB4; #100;
A = 8'hD1; B = 8'hB5; #100;
A = 8'hD1; B = 8'hB6; #100;
A = 8'hD1; B = 8'hB7; #100;
A = 8'hD1; B = 8'hB8; #100;
A = 8'hD1; B = 8'hB9; #100;
A = 8'hD1; B = 8'hBA; #100;
A = 8'hD1; B = 8'hBB; #100;
A = 8'hD1; B = 8'hBC; #100;
A = 8'hD1; B = 8'hBD; #100;
A = 8'hD1; B = 8'hBE; #100;
A = 8'hD1; B = 8'hBF; #100;
A = 8'hD1; B = 8'hC0; #100;
A = 8'hD1; B = 8'hC1; #100;
A = 8'hD1; B = 8'hC2; #100;
A = 8'hD1; B = 8'hC3; #100;
A = 8'hD1; B = 8'hC4; #100;
A = 8'hD1; B = 8'hC5; #100;
A = 8'hD1; B = 8'hC6; #100;
A = 8'hD1; B = 8'hC7; #100;
A = 8'hD1; B = 8'hC8; #100;
A = 8'hD1; B = 8'hC9; #100;
A = 8'hD1; B = 8'hCA; #100;
A = 8'hD1; B = 8'hCB; #100;
A = 8'hD1; B = 8'hCC; #100;
A = 8'hD1; B = 8'hCD; #100;
A = 8'hD1; B = 8'hCE; #100;
A = 8'hD1; B = 8'hCF; #100;
A = 8'hD1; B = 8'hD0; #100;
A = 8'hD1; B = 8'hD1; #100;
A = 8'hD1; B = 8'hD2; #100;
A = 8'hD1; B = 8'hD3; #100;
A = 8'hD1; B = 8'hD4; #100;
A = 8'hD1; B = 8'hD5; #100;
A = 8'hD1; B = 8'hD6; #100;
A = 8'hD1; B = 8'hD7; #100;
A = 8'hD1; B = 8'hD8; #100;
A = 8'hD1; B = 8'hD9; #100;
A = 8'hD1; B = 8'hDA; #100;
A = 8'hD1; B = 8'hDB; #100;
A = 8'hD1; B = 8'hDC; #100;
A = 8'hD1; B = 8'hDD; #100;
A = 8'hD1; B = 8'hDE; #100;
A = 8'hD1; B = 8'hDF; #100;
A = 8'hD1; B = 8'hE0; #100;
A = 8'hD1; B = 8'hE1; #100;
A = 8'hD1; B = 8'hE2; #100;
A = 8'hD1; B = 8'hE3; #100;
A = 8'hD1; B = 8'hE4; #100;
A = 8'hD1; B = 8'hE5; #100;
A = 8'hD1; B = 8'hE6; #100;
A = 8'hD1; B = 8'hE7; #100;
A = 8'hD1; B = 8'hE8; #100;
A = 8'hD1; B = 8'hE9; #100;
A = 8'hD1; B = 8'hEA; #100;
A = 8'hD1; B = 8'hEB; #100;
A = 8'hD1; B = 8'hEC; #100;
A = 8'hD1; B = 8'hED; #100;
A = 8'hD1; B = 8'hEE; #100;
A = 8'hD1; B = 8'hEF; #100;
A = 8'hD1; B = 8'hF0; #100;
A = 8'hD1; B = 8'hF1; #100;
A = 8'hD1; B = 8'hF2; #100;
A = 8'hD1; B = 8'hF3; #100;
A = 8'hD1; B = 8'hF4; #100;
A = 8'hD1; B = 8'hF5; #100;
A = 8'hD1; B = 8'hF6; #100;
A = 8'hD1; B = 8'hF7; #100;
A = 8'hD1; B = 8'hF8; #100;
A = 8'hD1; B = 8'hF9; #100;
A = 8'hD1; B = 8'hFA; #100;
A = 8'hD1; B = 8'hFB; #100;
A = 8'hD1; B = 8'hFC; #100;
A = 8'hD1; B = 8'hFD; #100;
A = 8'hD1; B = 8'hFE; #100;
A = 8'hD1; B = 8'hFF; #100;
A = 8'hD2; B = 8'h0; #100;
A = 8'hD2; B = 8'h1; #100;
A = 8'hD2; B = 8'h2; #100;
A = 8'hD2; B = 8'h3; #100;
A = 8'hD2; B = 8'h4; #100;
A = 8'hD2; B = 8'h5; #100;
A = 8'hD2; B = 8'h6; #100;
A = 8'hD2; B = 8'h7; #100;
A = 8'hD2; B = 8'h8; #100;
A = 8'hD2; B = 8'h9; #100;
A = 8'hD2; B = 8'hA; #100;
A = 8'hD2; B = 8'hB; #100;
A = 8'hD2; B = 8'hC; #100;
A = 8'hD2; B = 8'hD; #100;
A = 8'hD2; B = 8'hE; #100;
A = 8'hD2; B = 8'hF; #100;
A = 8'hD2; B = 8'h10; #100;
A = 8'hD2; B = 8'h11; #100;
A = 8'hD2; B = 8'h12; #100;
A = 8'hD2; B = 8'h13; #100;
A = 8'hD2; B = 8'h14; #100;
A = 8'hD2; B = 8'h15; #100;
A = 8'hD2; B = 8'h16; #100;
A = 8'hD2; B = 8'h17; #100;
A = 8'hD2; B = 8'h18; #100;
A = 8'hD2; B = 8'h19; #100;
A = 8'hD2; B = 8'h1A; #100;
A = 8'hD2; B = 8'h1B; #100;
A = 8'hD2; B = 8'h1C; #100;
A = 8'hD2; B = 8'h1D; #100;
A = 8'hD2; B = 8'h1E; #100;
A = 8'hD2; B = 8'h1F; #100;
A = 8'hD2; B = 8'h20; #100;
A = 8'hD2; B = 8'h21; #100;
A = 8'hD2; B = 8'h22; #100;
A = 8'hD2; B = 8'h23; #100;
A = 8'hD2; B = 8'h24; #100;
A = 8'hD2; B = 8'h25; #100;
A = 8'hD2; B = 8'h26; #100;
A = 8'hD2; B = 8'h27; #100;
A = 8'hD2; B = 8'h28; #100;
A = 8'hD2; B = 8'h29; #100;
A = 8'hD2; B = 8'h2A; #100;
A = 8'hD2; B = 8'h2B; #100;
A = 8'hD2; B = 8'h2C; #100;
A = 8'hD2; B = 8'h2D; #100;
A = 8'hD2; B = 8'h2E; #100;
A = 8'hD2; B = 8'h2F; #100;
A = 8'hD2; B = 8'h30; #100;
A = 8'hD2; B = 8'h31; #100;
A = 8'hD2; B = 8'h32; #100;
A = 8'hD2; B = 8'h33; #100;
A = 8'hD2; B = 8'h34; #100;
A = 8'hD2; B = 8'h35; #100;
A = 8'hD2; B = 8'h36; #100;
A = 8'hD2; B = 8'h37; #100;
A = 8'hD2; B = 8'h38; #100;
A = 8'hD2; B = 8'h39; #100;
A = 8'hD2; B = 8'h3A; #100;
A = 8'hD2; B = 8'h3B; #100;
A = 8'hD2; B = 8'h3C; #100;
A = 8'hD2; B = 8'h3D; #100;
A = 8'hD2; B = 8'h3E; #100;
A = 8'hD2; B = 8'h3F; #100;
A = 8'hD2; B = 8'h40; #100;
A = 8'hD2; B = 8'h41; #100;
A = 8'hD2; B = 8'h42; #100;
A = 8'hD2; B = 8'h43; #100;
A = 8'hD2; B = 8'h44; #100;
A = 8'hD2; B = 8'h45; #100;
A = 8'hD2; B = 8'h46; #100;
A = 8'hD2; B = 8'h47; #100;
A = 8'hD2; B = 8'h48; #100;
A = 8'hD2; B = 8'h49; #100;
A = 8'hD2; B = 8'h4A; #100;
A = 8'hD2; B = 8'h4B; #100;
A = 8'hD2; B = 8'h4C; #100;
A = 8'hD2; B = 8'h4D; #100;
A = 8'hD2; B = 8'h4E; #100;
A = 8'hD2; B = 8'h4F; #100;
A = 8'hD2; B = 8'h50; #100;
A = 8'hD2; B = 8'h51; #100;
A = 8'hD2; B = 8'h52; #100;
A = 8'hD2; B = 8'h53; #100;
A = 8'hD2; B = 8'h54; #100;
A = 8'hD2; B = 8'h55; #100;
A = 8'hD2; B = 8'h56; #100;
A = 8'hD2; B = 8'h57; #100;
A = 8'hD2; B = 8'h58; #100;
A = 8'hD2; B = 8'h59; #100;
A = 8'hD2; B = 8'h5A; #100;
A = 8'hD2; B = 8'h5B; #100;
A = 8'hD2; B = 8'h5C; #100;
A = 8'hD2; B = 8'h5D; #100;
A = 8'hD2; B = 8'h5E; #100;
A = 8'hD2; B = 8'h5F; #100;
A = 8'hD2; B = 8'h60; #100;
A = 8'hD2; B = 8'h61; #100;
A = 8'hD2; B = 8'h62; #100;
A = 8'hD2; B = 8'h63; #100;
A = 8'hD2; B = 8'h64; #100;
A = 8'hD2; B = 8'h65; #100;
A = 8'hD2; B = 8'h66; #100;
A = 8'hD2; B = 8'h67; #100;
A = 8'hD2; B = 8'h68; #100;
A = 8'hD2; B = 8'h69; #100;
A = 8'hD2; B = 8'h6A; #100;
A = 8'hD2; B = 8'h6B; #100;
A = 8'hD2; B = 8'h6C; #100;
A = 8'hD2; B = 8'h6D; #100;
A = 8'hD2; B = 8'h6E; #100;
A = 8'hD2; B = 8'h6F; #100;
A = 8'hD2; B = 8'h70; #100;
A = 8'hD2; B = 8'h71; #100;
A = 8'hD2; B = 8'h72; #100;
A = 8'hD2; B = 8'h73; #100;
A = 8'hD2; B = 8'h74; #100;
A = 8'hD2; B = 8'h75; #100;
A = 8'hD2; B = 8'h76; #100;
A = 8'hD2; B = 8'h77; #100;
A = 8'hD2; B = 8'h78; #100;
A = 8'hD2; B = 8'h79; #100;
A = 8'hD2; B = 8'h7A; #100;
A = 8'hD2; B = 8'h7B; #100;
A = 8'hD2; B = 8'h7C; #100;
A = 8'hD2; B = 8'h7D; #100;
A = 8'hD2; B = 8'h7E; #100;
A = 8'hD2; B = 8'h7F; #100;
A = 8'hD2; B = 8'h80; #100;
A = 8'hD2; B = 8'h81; #100;
A = 8'hD2; B = 8'h82; #100;
A = 8'hD2; B = 8'h83; #100;
A = 8'hD2; B = 8'h84; #100;
A = 8'hD2; B = 8'h85; #100;
A = 8'hD2; B = 8'h86; #100;
A = 8'hD2; B = 8'h87; #100;
A = 8'hD2; B = 8'h88; #100;
A = 8'hD2; B = 8'h89; #100;
A = 8'hD2; B = 8'h8A; #100;
A = 8'hD2; B = 8'h8B; #100;
A = 8'hD2; B = 8'h8C; #100;
A = 8'hD2; B = 8'h8D; #100;
A = 8'hD2; B = 8'h8E; #100;
A = 8'hD2; B = 8'h8F; #100;
A = 8'hD2; B = 8'h90; #100;
A = 8'hD2; B = 8'h91; #100;
A = 8'hD2; B = 8'h92; #100;
A = 8'hD2; B = 8'h93; #100;
A = 8'hD2; B = 8'h94; #100;
A = 8'hD2; B = 8'h95; #100;
A = 8'hD2; B = 8'h96; #100;
A = 8'hD2; B = 8'h97; #100;
A = 8'hD2; B = 8'h98; #100;
A = 8'hD2; B = 8'h99; #100;
A = 8'hD2; B = 8'h9A; #100;
A = 8'hD2; B = 8'h9B; #100;
A = 8'hD2; B = 8'h9C; #100;
A = 8'hD2; B = 8'h9D; #100;
A = 8'hD2; B = 8'h9E; #100;
A = 8'hD2; B = 8'h9F; #100;
A = 8'hD2; B = 8'hA0; #100;
A = 8'hD2; B = 8'hA1; #100;
A = 8'hD2; B = 8'hA2; #100;
A = 8'hD2; B = 8'hA3; #100;
A = 8'hD2; B = 8'hA4; #100;
A = 8'hD2; B = 8'hA5; #100;
A = 8'hD2; B = 8'hA6; #100;
A = 8'hD2; B = 8'hA7; #100;
A = 8'hD2; B = 8'hA8; #100;
A = 8'hD2; B = 8'hA9; #100;
A = 8'hD2; B = 8'hAA; #100;
A = 8'hD2; B = 8'hAB; #100;
A = 8'hD2; B = 8'hAC; #100;
A = 8'hD2; B = 8'hAD; #100;
A = 8'hD2; B = 8'hAE; #100;
A = 8'hD2; B = 8'hAF; #100;
A = 8'hD2; B = 8'hB0; #100;
A = 8'hD2; B = 8'hB1; #100;
A = 8'hD2; B = 8'hB2; #100;
A = 8'hD2; B = 8'hB3; #100;
A = 8'hD2; B = 8'hB4; #100;
A = 8'hD2; B = 8'hB5; #100;
A = 8'hD2; B = 8'hB6; #100;
A = 8'hD2; B = 8'hB7; #100;
A = 8'hD2; B = 8'hB8; #100;
A = 8'hD2; B = 8'hB9; #100;
A = 8'hD2; B = 8'hBA; #100;
A = 8'hD2; B = 8'hBB; #100;
A = 8'hD2; B = 8'hBC; #100;
A = 8'hD2; B = 8'hBD; #100;
A = 8'hD2; B = 8'hBE; #100;
A = 8'hD2; B = 8'hBF; #100;
A = 8'hD2; B = 8'hC0; #100;
A = 8'hD2; B = 8'hC1; #100;
A = 8'hD2; B = 8'hC2; #100;
A = 8'hD2; B = 8'hC3; #100;
A = 8'hD2; B = 8'hC4; #100;
A = 8'hD2; B = 8'hC5; #100;
A = 8'hD2; B = 8'hC6; #100;
A = 8'hD2; B = 8'hC7; #100;
A = 8'hD2; B = 8'hC8; #100;
A = 8'hD2; B = 8'hC9; #100;
A = 8'hD2; B = 8'hCA; #100;
A = 8'hD2; B = 8'hCB; #100;
A = 8'hD2; B = 8'hCC; #100;
A = 8'hD2; B = 8'hCD; #100;
A = 8'hD2; B = 8'hCE; #100;
A = 8'hD2; B = 8'hCF; #100;
A = 8'hD2; B = 8'hD0; #100;
A = 8'hD2; B = 8'hD1; #100;
A = 8'hD2; B = 8'hD2; #100;
A = 8'hD2; B = 8'hD3; #100;
A = 8'hD2; B = 8'hD4; #100;
A = 8'hD2; B = 8'hD5; #100;
A = 8'hD2; B = 8'hD6; #100;
A = 8'hD2; B = 8'hD7; #100;
A = 8'hD2; B = 8'hD8; #100;
A = 8'hD2; B = 8'hD9; #100;
A = 8'hD2; B = 8'hDA; #100;
A = 8'hD2; B = 8'hDB; #100;
A = 8'hD2; B = 8'hDC; #100;
A = 8'hD2; B = 8'hDD; #100;
A = 8'hD2; B = 8'hDE; #100;
A = 8'hD2; B = 8'hDF; #100;
A = 8'hD2; B = 8'hE0; #100;
A = 8'hD2; B = 8'hE1; #100;
A = 8'hD2; B = 8'hE2; #100;
A = 8'hD2; B = 8'hE3; #100;
A = 8'hD2; B = 8'hE4; #100;
A = 8'hD2; B = 8'hE5; #100;
A = 8'hD2; B = 8'hE6; #100;
A = 8'hD2; B = 8'hE7; #100;
A = 8'hD2; B = 8'hE8; #100;
A = 8'hD2; B = 8'hE9; #100;
A = 8'hD2; B = 8'hEA; #100;
A = 8'hD2; B = 8'hEB; #100;
A = 8'hD2; B = 8'hEC; #100;
A = 8'hD2; B = 8'hED; #100;
A = 8'hD2; B = 8'hEE; #100;
A = 8'hD2; B = 8'hEF; #100;
A = 8'hD2; B = 8'hF0; #100;
A = 8'hD2; B = 8'hF1; #100;
A = 8'hD2; B = 8'hF2; #100;
A = 8'hD2; B = 8'hF3; #100;
A = 8'hD2; B = 8'hF4; #100;
A = 8'hD2; B = 8'hF5; #100;
A = 8'hD2; B = 8'hF6; #100;
A = 8'hD2; B = 8'hF7; #100;
A = 8'hD2; B = 8'hF8; #100;
A = 8'hD2; B = 8'hF9; #100;
A = 8'hD2; B = 8'hFA; #100;
A = 8'hD2; B = 8'hFB; #100;
A = 8'hD2; B = 8'hFC; #100;
A = 8'hD2; B = 8'hFD; #100;
A = 8'hD2; B = 8'hFE; #100;
A = 8'hD2; B = 8'hFF; #100;
A = 8'hD3; B = 8'h0; #100;
A = 8'hD3; B = 8'h1; #100;
A = 8'hD3; B = 8'h2; #100;
A = 8'hD3; B = 8'h3; #100;
A = 8'hD3; B = 8'h4; #100;
A = 8'hD3; B = 8'h5; #100;
A = 8'hD3; B = 8'h6; #100;
A = 8'hD3; B = 8'h7; #100;
A = 8'hD3; B = 8'h8; #100;
A = 8'hD3; B = 8'h9; #100;
A = 8'hD3; B = 8'hA; #100;
A = 8'hD3; B = 8'hB; #100;
A = 8'hD3; B = 8'hC; #100;
A = 8'hD3; B = 8'hD; #100;
A = 8'hD3; B = 8'hE; #100;
A = 8'hD3; B = 8'hF; #100;
A = 8'hD3; B = 8'h10; #100;
A = 8'hD3; B = 8'h11; #100;
A = 8'hD3; B = 8'h12; #100;
A = 8'hD3; B = 8'h13; #100;
A = 8'hD3; B = 8'h14; #100;
A = 8'hD3; B = 8'h15; #100;
A = 8'hD3; B = 8'h16; #100;
A = 8'hD3; B = 8'h17; #100;
A = 8'hD3; B = 8'h18; #100;
A = 8'hD3; B = 8'h19; #100;
A = 8'hD3; B = 8'h1A; #100;
A = 8'hD3; B = 8'h1B; #100;
A = 8'hD3; B = 8'h1C; #100;
A = 8'hD3; B = 8'h1D; #100;
A = 8'hD3; B = 8'h1E; #100;
A = 8'hD3; B = 8'h1F; #100;
A = 8'hD3; B = 8'h20; #100;
A = 8'hD3; B = 8'h21; #100;
A = 8'hD3; B = 8'h22; #100;
A = 8'hD3; B = 8'h23; #100;
A = 8'hD3; B = 8'h24; #100;
A = 8'hD3; B = 8'h25; #100;
A = 8'hD3; B = 8'h26; #100;
A = 8'hD3; B = 8'h27; #100;
A = 8'hD3; B = 8'h28; #100;
A = 8'hD3; B = 8'h29; #100;
A = 8'hD3; B = 8'h2A; #100;
A = 8'hD3; B = 8'h2B; #100;
A = 8'hD3; B = 8'h2C; #100;
A = 8'hD3; B = 8'h2D; #100;
A = 8'hD3; B = 8'h2E; #100;
A = 8'hD3; B = 8'h2F; #100;
A = 8'hD3; B = 8'h30; #100;
A = 8'hD3; B = 8'h31; #100;
A = 8'hD3; B = 8'h32; #100;
A = 8'hD3; B = 8'h33; #100;
A = 8'hD3; B = 8'h34; #100;
A = 8'hD3; B = 8'h35; #100;
A = 8'hD3; B = 8'h36; #100;
A = 8'hD3; B = 8'h37; #100;
A = 8'hD3; B = 8'h38; #100;
A = 8'hD3; B = 8'h39; #100;
A = 8'hD3; B = 8'h3A; #100;
A = 8'hD3; B = 8'h3B; #100;
A = 8'hD3; B = 8'h3C; #100;
A = 8'hD3; B = 8'h3D; #100;
A = 8'hD3; B = 8'h3E; #100;
A = 8'hD3; B = 8'h3F; #100;
A = 8'hD3; B = 8'h40; #100;
A = 8'hD3; B = 8'h41; #100;
A = 8'hD3; B = 8'h42; #100;
A = 8'hD3; B = 8'h43; #100;
A = 8'hD3; B = 8'h44; #100;
A = 8'hD3; B = 8'h45; #100;
A = 8'hD3; B = 8'h46; #100;
A = 8'hD3; B = 8'h47; #100;
A = 8'hD3; B = 8'h48; #100;
A = 8'hD3; B = 8'h49; #100;
A = 8'hD3; B = 8'h4A; #100;
A = 8'hD3; B = 8'h4B; #100;
A = 8'hD3; B = 8'h4C; #100;
A = 8'hD3; B = 8'h4D; #100;
A = 8'hD3; B = 8'h4E; #100;
A = 8'hD3; B = 8'h4F; #100;
A = 8'hD3; B = 8'h50; #100;
A = 8'hD3; B = 8'h51; #100;
A = 8'hD3; B = 8'h52; #100;
A = 8'hD3; B = 8'h53; #100;
A = 8'hD3; B = 8'h54; #100;
A = 8'hD3; B = 8'h55; #100;
A = 8'hD3; B = 8'h56; #100;
A = 8'hD3; B = 8'h57; #100;
A = 8'hD3; B = 8'h58; #100;
A = 8'hD3; B = 8'h59; #100;
A = 8'hD3; B = 8'h5A; #100;
A = 8'hD3; B = 8'h5B; #100;
A = 8'hD3; B = 8'h5C; #100;
A = 8'hD3; B = 8'h5D; #100;
A = 8'hD3; B = 8'h5E; #100;
A = 8'hD3; B = 8'h5F; #100;
A = 8'hD3; B = 8'h60; #100;
A = 8'hD3; B = 8'h61; #100;
A = 8'hD3; B = 8'h62; #100;
A = 8'hD3; B = 8'h63; #100;
A = 8'hD3; B = 8'h64; #100;
A = 8'hD3; B = 8'h65; #100;
A = 8'hD3; B = 8'h66; #100;
A = 8'hD3; B = 8'h67; #100;
A = 8'hD3; B = 8'h68; #100;
A = 8'hD3; B = 8'h69; #100;
A = 8'hD3; B = 8'h6A; #100;
A = 8'hD3; B = 8'h6B; #100;
A = 8'hD3; B = 8'h6C; #100;
A = 8'hD3; B = 8'h6D; #100;
A = 8'hD3; B = 8'h6E; #100;
A = 8'hD3; B = 8'h6F; #100;
A = 8'hD3; B = 8'h70; #100;
A = 8'hD3; B = 8'h71; #100;
A = 8'hD3; B = 8'h72; #100;
A = 8'hD3; B = 8'h73; #100;
A = 8'hD3; B = 8'h74; #100;
A = 8'hD3; B = 8'h75; #100;
A = 8'hD3; B = 8'h76; #100;
A = 8'hD3; B = 8'h77; #100;
A = 8'hD3; B = 8'h78; #100;
A = 8'hD3; B = 8'h79; #100;
A = 8'hD3; B = 8'h7A; #100;
A = 8'hD3; B = 8'h7B; #100;
A = 8'hD3; B = 8'h7C; #100;
A = 8'hD3; B = 8'h7D; #100;
A = 8'hD3; B = 8'h7E; #100;
A = 8'hD3; B = 8'h7F; #100;
A = 8'hD3; B = 8'h80; #100;
A = 8'hD3; B = 8'h81; #100;
A = 8'hD3; B = 8'h82; #100;
A = 8'hD3; B = 8'h83; #100;
A = 8'hD3; B = 8'h84; #100;
A = 8'hD3; B = 8'h85; #100;
A = 8'hD3; B = 8'h86; #100;
A = 8'hD3; B = 8'h87; #100;
A = 8'hD3; B = 8'h88; #100;
A = 8'hD3; B = 8'h89; #100;
A = 8'hD3; B = 8'h8A; #100;
A = 8'hD3; B = 8'h8B; #100;
A = 8'hD3; B = 8'h8C; #100;
A = 8'hD3; B = 8'h8D; #100;
A = 8'hD3; B = 8'h8E; #100;
A = 8'hD3; B = 8'h8F; #100;
A = 8'hD3; B = 8'h90; #100;
A = 8'hD3; B = 8'h91; #100;
A = 8'hD3; B = 8'h92; #100;
A = 8'hD3; B = 8'h93; #100;
A = 8'hD3; B = 8'h94; #100;
A = 8'hD3; B = 8'h95; #100;
A = 8'hD3; B = 8'h96; #100;
A = 8'hD3; B = 8'h97; #100;
A = 8'hD3; B = 8'h98; #100;
A = 8'hD3; B = 8'h99; #100;
A = 8'hD3; B = 8'h9A; #100;
A = 8'hD3; B = 8'h9B; #100;
A = 8'hD3; B = 8'h9C; #100;
A = 8'hD3; B = 8'h9D; #100;
A = 8'hD3; B = 8'h9E; #100;
A = 8'hD3; B = 8'h9F; #100;
A = 8'hD3; B = 8'hA0; #100;
A = 8'hD3; B = 8'hA1; #100;
A = 8'hD3; B = 8'hA2; #100;
A = 8'hD3; B = 8'hA3; #100;
A = 8'hD3; B = 8'hA4; #100;
A = 8'hD3; B = 8'hA5; #100;
A = 8'hD3; B = 8'hA6; #100;
A = 8'hD3; B = 8'hA7; #100;
A = 8'hD3; B = 8'hA8; #100;
A = 8'hD3; B = 8'hA9; #100;
A = 8'hD3; B = 8'hAA; #100;
A = 8'hD3; B = 8'hAB; #100;
A = 8'hD3; B = 8'hAC; #100;
A = 8'hD3; B = 8'hAD; #100;
A = 8'hD3; B = 8'hAE; #100;
A = 8'hD3; B = 8'hAF; #100;
A = 8'hD3; B = 8'hB0; #100;
A = 8'hD3; B = 8'hB1; #100;
A = 8'hD3; B = 8'hB2; #100;
A = 8'hD3; B = 8'hB3; #100;
A = 8'hD3; B = 8'hB4; #100;
A = 8'hD3; B = 8'hB5; #100;
A = 8'hD3; B = 8'hB6; #100;
A = 8'hD3; B = 8'hB7; #100;
A = 8'hD3; B = 8'hB8; #100;
A = 8'hD3; B = 8'hB9; #100;
A = 8'hD3; B = 8'hBA; #100;
A = 8'hD3; B = 8'hBB; #100;
A = 8'hD3; B = 8'hBC; #100;
A = 8'hD3; B = 8'hBD; #100;
A = 8'hD3; B = 8'hBE; #100;
A = 8'hD3; B = 8'hBF; #100;
A = 8'hD3; B = 8'hC0; #100;
A = 8'hD3; B = 8'hC1; #100;
A = 8'hD3; B = 8'hC2; #100;
A = 8'hD3; B = 8'hC3; #100;
A = 8'hD3; B = 8'hC4; #100;
A = 8'hD3; B = 8'hC5; #100;
A = 8'hD3; B = 8'hC6; #100;
A = 8'hD3; B = 8'hC7; #100;
A = 8'hD3; B = 8'hC8; #100;
A = 8'hD3; B = 8'hC9; #100;
A = 8'hD3; B = 8'hCA; #100;
A = 8'hD3; B = 8'hCB; #100;
A = 8'hD3; B = 8'hCC; #100;
A = 8'hD3; B = 8'hCD; #100;
A = 8'hD3; B = 8'hCE; #100;
A = 8'hD3; B = 8'hCF; #100;
A = 8'hD3; B = 8'hD0; #100;
A = 8'hD3; B = 8'hD1; #100;
A = 8'hD3; B = 8'hD2; #100;
A = 8'hD3; B = 8'hD3; #100;
A = 8'hD3; B = 8'hD4; #100;
A = 8'hD3; B = 8'hD5; #100;
A = 8'hD3; B = 8'hD6; #100;
A = 8'hD3; B = 8'hD7; #100;
A = 8'hD3; B = 8'hD8; #100;
A = 8'hD3; B = 8'hD9; #100;
A = 8'hD3; B = 8'hDA; #100;
A = 8'hD3; B = 8'hDB; #100;
A = 8'hD3; B = 8'hDC; #100;
A = 8'hD3; B = 8'hDD; #100;
A = 8'hD3; B = 8'hDE; #100;
A = 8'hD3; B = 8'hDF; #100;
A = 8'hD3; B = 8'hE0; #100;
A = 8'hD3; B = 8'hE1; #100;
A = 8'hD3; B = 8'hE2; #100;
A = 8'hD3; B = 8'hE3; #100;
A = 8'hD3; B = 8'hE4; #100;
A = 8'hD3; B = 8'hE5; #100;
A = 8'hD3; B = 8'hE6; #100;
A = 8'hD3; B = 8'hE7; #100;
A = 8'hD3; B = 8'hE8; #100;
A = 8'hD3; B = 8'hE9; #100;
A = 8'hD3; B = 8'hEA; #100;
A = 8'hD3; B = 8'hEB; #100;
A = 8'hD3; B = 8'hEC; #100;
A = 8'hD3; B = 8'hED; #100;
A = 8'hD3; B = 8'hEE; #100;
A = 8'hD3; B = 8'hEF; #100;
A = 8'hD3; B = 8'hF0; #100;
A = 8'hD3; B = 8'hF1; #100;
A = 8'hD3; B = 8'hF2; #100;
A = 8'hD3; B = 8'hF3; #100;
A = 8'hD3; B = 8'hF4; #100;
A = 8'hD3; B = 8'hF5; #100;
A = 8'hD3; B = 8'hF6; #100;
A = 8'hD3; B = 8'hF7; #100;
A = 8'hD3; B = 8'hF8; #100;
A = 8'hD3; B = 8'hF9; #100;
A = 8'hD3; B = 8'hFA; #100;
A = 8'hD3; B = 8'hFB; #100;
A = 8'hD3; B = 8'hFC; #100;
A = 8'hD3; B = 8'hFD; #100;
A = 8'hD3; B = 8'hFE; #100;
A = 8'hD3; B = 8'hFF; #100;
A = 8'hD4; B = 8'h0; #100;
A = 8'hD4; B = 8'h1; #100;
A = 8'hD4; B = 8'h2; #100;
A = 8'hD4; B = 8'h3; #100;
A = 8'hD4; B = 8'h4; #100;
A = 8'hD4; B = 8'h5; #100;
A = 8'hD4; B = 8'h6; #100;
A = 8'hD4; B = 8'h7; #100;
A = 8'hD4; B = 8'h8; #100;
A = 8'hD4; B = 8'h9; #100;
A = 8'hD4; B = 8'hA; #100;
A = 8'hD4; B = 8'hB; #100;
A = 8'hD4; B = 8'hC; #100;
A = 8'hD4; B = 8'hD; #100;
A = 8'hD4; B = 8'hE; #100;
A = 8'hD4; B = 8'hF; #100;
A = 8'hD4; B = 8'h10; #100;
A = 8'hD4; B = 8'h11; #100;
A = 8'hD4; B = 8'h12; #100;
A = 8'hD4; B = 8'h13; #100;
A = 8'hD4; B = 8'h14; #100;
A = 8'hD4; B = 8'h15; #100;
A = 8'hD4; B = 8'h16; #100;
A = 8'hD4; B = 8'h17; #100;
A = 8'hD4; B = 8'h18; #100;
A = 8'hD4; B = 8'h19; #100;
A = 8'hD4; B = 8'h1A; #100;
A = 8'hD4; B = 8'h1B; #100;
A = 8'hD4; B = 8'h1C; #100;
A = 8'hD4; B = 8'h1D; #100;
A = 8'hD4; B = 8'h1E; #100;
A = 8'hD4; B = 8'h1F; #100;
A = 8'hD4; B = 8'h20; #100;
A = 8'hD4; B = 8'h21; #100;
A = 8'hD4; B = 8'h22; #100;
A = 8'hD4; B = 8'h23; #100;
A = 8'hD4; B = 8'h24; #100;
A = 8'hD4; B = 8'h25; #100;
A = 8'hD4; B = 8'h26; #100;
A = 8'hD4; B = 8'h27; #100;
A = 8'hD4; B = 8'h28; #100;
A = 8'hD4; B = 8'h29; #100;
A = 8'hD4; B = 8'h2A; #100;
A = 8'hD4; B = 8'h2B; #100;
A = 8'hD4; B = 8'h2C; #100;
A = 8'hD4; B = 8'h2D; #100;
A = 8'hD4; B = 8'h2E; #100;
A = 8'hD4; B = 8'h2F; #100;
A = 8'hD4; B = 8'h30; #100;
A = 8'hD4; B = 8'h31; #100;
A = 8'hD4; B = 8'h32; #100;
A = 8'hD4; B = 8'h33; #100;
A = 8'hD4; B = 8'h34; #100;
A = 8'hD4; B = 8'h35; #100;
A = 8'hD4; B = 8'h36; #100;
A = 8'hD4; B = 8'h37; #100;
A = 8'hD4; B = 8'h38; #100;
A = 8'hD4; B = 8'h39; #100;
A = 8'hD4; B = 8'h3A; #100;
A = 8'hD4; B = 8'h3B; #100;
A = 8'hD4; B = 8'h3C; #100;
A = 8'hD4; B = 8'h3D; #100;
A = 8'hD4; B = 8'h3E; #100;
A = 8'hD4; B = 8'h3F; #100;
A = 8'hD4; B = 8'h40; #100;
A = 8'hD4; B = 8'h41; #100;
A = 8'hD4; B = 8'h42; #100;
A = 8'hD4; B = 8'h43; #100;
A = 8'hD4; B = 8'h44; #100;
A = 8'hD4; B = 8'h45; #100;
A = 8'hD4; B = 8'h46; #100;
A = 8'hD4; B = 8'h47; #100;
A = 8'hD4; B = 8'h48; #100;
A = 8'hD4; B = 8'h49; #100;
A = 8'hD4; B = 8'h4A; #100;
A = 8'hD4; B = 8'h4B; #100;
A = 8'hD4; B = 8'h4C; #100;
A = 8'hD4; B = 8'h4D; #100;
A = 8'hD4; B = 8'h4E; #100;
A = 8'hD4; B = 8'h4F; #100;
A = 8'hD4; B = 8'h50; #100;
A = 8'hD4; B = 8'h51; #100;
A = 8'hD4; B = 8'h52; #100;
A = 8'hD4; B = 8'h53; #100;
A = 8'hD4; B = 8'h54; #100;
A = 8'hD4; B = 8'h55; #100;
A = 8'hD4; B = 8'h56; #100;
A = 8'hD4; B = 8'h57; #100;
A = 8'hD4; B = 8'h58; #100;
A = 8'hD4; B = 8'h59; #100;
A = 8'hD4; B = 8'h5A; #100;
A = 8'hD4; B = 8'h5B; #100;
A = 8'hD4; B = 8'h5C; #100;
A = 8'hD4; B = 8'h5D; #100;
A = 8'hD4; B = 8'h5E; #100;
A = 8'hD4; B = 8'h5F; #100;
A = 8'hD4; B = 8'h60; #100;
A = 8'hD4; B = 8'h61; #100;
A = 8'hD4; B = 8'h62; #100;
A = 8'hD4; B = 8'h63; #100;
A = 8'hD4; B = 8'h64; #100;
A = 8'hD4; B = 8'h65; #100;
A = 8'hD4; B = 8'h66; #100;
A = 8'hD4; B = 8'h67; #100;
A = 8'hD4; B = 8'h68; #100;
A = 8'hD4; B = 8'h69; #100;
A = 8'hD4; B = 8'h6A; #100;
A = 8'hD4; B = 8'h6B; #100;
A = 8'hD4; B = 8'h6C; #100;
A = 8'hD4; B = 8'h6D; #100;
A = 8'hD4; B = 8'h6E; #100;
A = 8'hD4; B = 8'h6F; #100;
A = 8'hD4; B = 8'h70; #100;
A = 8'hD4; B = 8'h71; #100;
A = 8'hD4; B = 8'h72; #100;
A = 8'hD4; B = 8'h73; #100;
A = 8'hD4; B = 8'h74; #100;
A = 8'hD4; B = 8'h75; #100;
A = 8'hD4; B = 8'h76; #100;
A = 8'hD4; B = 8'h77; #100;
A = 8'hD4; B = 8'h78; #100;
A = 8'hD4; B = 8'h79; #100;
A = 8'hD4; B = 8'h7A; #100;
A = 8'hD4; B = 8'h7B; #100;
A = 8'hD4; B = 8'h7C; #100;
A = 8'hD4; B = 8'h7D; #100;
A = 8'hD4; B = 8'h7E; #100;
A = 8'hD4; B = 8'h7F; #100;
A = 8'hD4; B = 8'h80; #100;
A = 8'hD4; B = 8'h81; #100;
A = 8'hD4; B = 8'h82; #100;
A = 8'hD4; B = 8'h83; #100;
A = 8'hD4; B = 8'h84; #100;
A = 8'hD4; B = 8'h85; #100;
A = 8'hD4; B = 8'h86; #100;
A = 8'hD4; B = 8'h87; #100;
A = 8'hD4; B = 8'h88; #100;
A = 8'hD4; B = 8'h89; #100;
A = 8'hD4; B = 8'h8A; #100;
A = 8'hD4; B = 8'h8B; #100;
A = 8'hD4; B = 8'h8C; #100;
A = 8'hD4; B = 8'h8D; #100;
A = 8'hD4; B = 8'h8E; #100;
A = 8'hD4; B = 8'h8F; #100;
A = 8'hD4; B = 8'h90; #100;
A = 8'hD4; B = 8'h91; #100;
A = 8'hD4; B = 8'h92; #100;
A = 8'hD4; B = 8'h93; #100;
A = 8'hD4; B = 8'h94; #100;
A = 8'hD4; B = 8'h95; #100;
A = 8'hD4; B = 8'h96; #100;
A = 8'hD4; B = 8'h97; #100;
A = 8'hD4; B = 8'h98; #100;
A = 8'hD4; B = 8'h99; #100;
A = 8'hD4; B = 8'h9A; #100;
A = 8'hD4; B = 8'h9B; #100;
A = 8'hD4; B = 8'h9C; #100;
A = 8'hD4; B = 8'h9D; #100;
A = 8'hD4; B = 8'h9E; #100;
A = 8'hD4; B = 8'h9F; #100;
A = 8'hD4; B = 8'hA0; #100;
A = 8'hD4; B = 8'hA1; #100;
A = 8'hD4; B = 8'hA2; #100;
A = 8'hD4; B = 8'hA3; #100;
A = 8'hD4; B = 8'hA4; #100;
A = 8'hD4; B = 8'hA5; #100;
A = 8'hD4; B = 8'hA6; #100;
A = 8'hD4; B = 8'hA7; #100;
A = 8'hD4; B = 8'hA8; #100;
A = 8'hD4; B = 8'hA9; #100;
A = 8'hD4; B = 8'hAA; #100;
A = 8'hD4; B = 8'hAB; #100;
A = 8'hD4; B = 8'hAC; #100;
A = 8'hD4; B = 8'hAD; #100;
A = 8'hD4; B = 8'hAE; #100;
A = 8'hD4; B = 8'hAF; #100;
A = 8'hD4; B = 8'hB0; #100;
A = 8'hD4; B = 8'hB1; #100;
A = 8'hD4; B = 8'hB2; #100;
A = 8'hD4; B = 8'hB3; #100;
A = 8'hD4; B = 8'hB4; #100;
A = 8'hD4; B = 8'hB5; #100;
A = 8'hD4; B = 8'hB6; #100;
A = 8'hD4; B = 8'hB7; #100;
A = 8'hD4; B = 8'hB8; #100;
A = 8'hD4; B = 8'hB9; #100;
A = 8'hD4; B = 8'hBA; #100;
A = 8'hD4; B = 8'hBB; #100;
A = 8'hD4; B = 8'hBC; #100;
A = 8'hD4; B = 8'hBD; #100;
A = 8'hD4; B = 8'hBE; #100;
A = 8'hD4; B = 8'hBF; #100;
A = 8'hD4; B = 8'hC0; #100;
A = 8'hD4; B = 8'hC1; #100;
A = 8'hD4; B = 8'hC2; #100;
A = 8'hD4; B = 8'hC3; #100;
A = 8'hD4; B = 8'hC4; #100;
A = 8'hD4; B = 8'hC5; #100;
A = 8'hD4; B = 8'hC6; #100;
A = 8'hD4; B = 8'hC7; #100;
A = 8'hD4; B = 8'hC8; #100;
A = 8'hD4; B = 8'hC9; #100;
A = 8'hD4; B = 8'hCA; #100;
A = 8'hD4; B = 8'hCB; #100;
A = 8'hD4; B = 8'hCC; #100;
A = 8'hD4; B = 8'hCD; #100;
A = 8'hD4; B = 8'hCE; #100;
A = 8'hD4; B = 8'hCF; #100;
A = 8'hD4; B = 8'hD0; #100;
A = 8'hD4; B = 8'hD1; #100;
A = 8'hD4; B = 8'hD2; #100;
A = 8'hD4; B = 8'hD3; #100;
A = 8'hD4; B = 8'hD4; #100;
A = 8'hD4; B = 8'hD5; #100;
A = 8'hD4; B = 8'hD6; #100;
A = 8'hD4; B = 8'hD7; #100;
A = 8'hD4; B = 8'hD8; #100;
A = 8'hD4; B = 8'hD9; #100;
A = 8'hD4; B = 8'hDA; #100;
A = 8'hD4; B = 8'hDB; #100;
A = 8'hD4; B = 8'hDC; #100;
A = 8'hD4; B = 8'hDD; #100;
A = 8'hD4; B = 8'hDE; #100;
A = 8'hD4; B = 8'hDF; #100;
A = 8'hD4; B = 8'hE0; #100;
A = 8'hD4; B = 8'hE1; #100;
A = 8'hD4; B = 8'hE2; #100;
A = 8'hD4; B = 8'hE3; #100;
A = 8'hD4; B = 8'hE4; #100;
A = 8'hD4; B = 8'hE5; #100;
A = 8'hD4; B = 8'hE6; #100;
A = 8'hD4; B = 8'hE7; #100;
A = 8'hD4; B = 8'hE8; #100;
A = 8'hD4; B = 8'hE9; #100;
A = 8'hD4; B = 8'hEA; #100;
A = 8'hD4; B = 8'hEB; #100;
A = 8'hD4; B = 8'hEC; #100;
A = 8'hD4; B = 8'hED; #100;
A = 8'hD4; B = 8'hEE; #100;
A = 8'hD4; B = 8'hEF; #100;
A = 8'hD4; B = 8'hF0; #100;
A = 8'hD4; B = 8'hF1; #100;
A = 8'hD4; B = 8'hF2; #100;
A = 8'hD4; B = 8'hF3; #100;
A = 8'hD4; B = 8'hF4; #100;
A = 8'hD4; B = 8'hF5; #100;
A = 8'hD4; B = 8'hF6; #100;
A = 8'hD4; B = 8'hF7; #100;
A = 8'hD4; B = 8'hF8; #100;
A = 8'hD4; B = 8'hF9; #100;
A = 8'hD4; B = 8'hFA; #100;
A = 8'hD4; B = 8'hFB; #100;
A = 8'hD4; B = 8'hFC; #100;
A = 8'hD4; B = 8'hFD; #100;
A = 8'hD4; B = 8'hFE; #100;
A = 8'hD4; B = 8'hFF; #100;
A = 8'hD5; B = 8'h0; #100;
A = 8'hD5; B = 8'h1; #100;
A = 8'hD5; B = 8'h2; #100;
A = 8'hD5; B = 8'h3; #100;
A = 8'hD5; B = 8'h4; #100;
A = 8'hD5; B = 8'h5; #100;
A = 8'hD5; B = 8'h6; #100;
A = 8'hD5; B = 8'h7; #100;
A = 8'hD5; B = 8'h8; #100;
A = 8'hD5; B = 8'h9; #100;
A = 8'hD5; B = 8'hA; #100;
A = 8'hD5; B = 8'hB; #100;
A = 8'hD5; B = 8'hC; #100;
A = 8'hD5; B = 8'hD; #100;
A = 8'hD5; B = 8'hE; #100;
A = 8'hD5; B = 8'hF; #100;
A = 8'hD5; B = 8'h10; #100;
A = 8'hD5; B = 8'h11; #100;
A = 8'hD5; B = 8'h12; #100;
A = 8'hD5; B = 8'h13; #100;
A = 8'hD5; B = 8'h14; #100;
A = 8'hD5; B = 8'h15; #100;
A = 8'hD5; B = 8'h16; #100;
A = 8'hD5; B = 8'h17; #100;
A = 8'hD5; B = 8'h18; #100;
A = 8'hD5; B = 8'h19; #100;
A = 8'hD5; B = 8'h1A; #100;
A = 8'hD5; B = 8'h1B; #100;
A = 8'hD5; B = 8'h1C; #100;
A = 8'hD5; B = 8'h1D; #100;
A = 8'hD5; B = 8'h1E; #100;
A = 8'hD5; B = 8'h1F; #100;
A = 8'hD5; B = 8'h20; #100;
A = 8'hD5; B = 8'h21; #100;
A = 8'hD5; B = 8'h22; #100;
A = 8'hD5; B = 8'h23; #100;
A = 8'hD5; B = 8'h24; #100;
A = 8'hD5; B = 8'h25; #100;
A = 8'hD5; B = 8'h26; #100;
A = 8'hD5; B = 8'h27; #100;
A = 8'hD5; B = 8'h28; #100;
A = 8'hD5; B = 8'h29; #100;
A = 8'hD5; B = 8'h2A; #100;
A = 8'hD5; B = 8'h2B; #100;
A = 8'hD5; B = 8'h2C; #100;
A = 8'hD5; B = 8'h2D; #100;
A = 8'hD5; B = 8'h2E; #100;
A = 8'hD5; B = 8'h2F; #100;
A = 8'hD5; B = 8'h30; #100;
A = 8'hD5; B = 8'h31; #100;
A = 8'hD5; B = 8'h32; #100;
A = 8'hD5; B = 8'h33; #100;
A = 8'hD5; B = 8'h34; #100;
A = 8'hD5; B = 8'h35; #100;
A = 8'hD5; B = 8'h36; #100;
A = 8'hD5; B = 8'h37; #100;
A = 8'hD5; B = 8'h38; #100;
A = 8'hD5; B = 8'h39; #100;
A = 8'hD5; B = 8'h3A; #100;
A = 8'hD5; B = 8'h3B; #100;
A = 8'hD5; B = 8'h3C; #100;
A = 8'hD5; B = 8'h3D; #100;
A = 8'hD5; B = 8'h3E; #100;
A = 8'hD5; B = 8'h3F; #100;
A = 8'hD5; B = 8'h40; #100;
A = 8'hD5; B = 8'h41; #100;
A = 8'hD5; B = 8'h42; #100;
A = 8'hD5; B = 8'h43; #100;
A = 8'hD5; B = 8'h44; #100;
A = 8'hD5; B = 8'h45; #100;
A = 8'hD5; B = 8'h46; #100;
A = 8'hD5; B = 8'h47; #100;
A = 8'hD5; B = 8'h48; #100;
A = 8'hD5; B = 8'h49; #100;
A = 8'hD5; B = 8'h4A; #100;
A = 8'hD5; B = 8'h4B; #100;
A = 8'hD5; B = 8'h4C; #100;
A = 8'hD5; B = 8'h4D; #100;
A = 8'hD5; B = 8'h4E; #100;
A = 8'hD5; B = 8'h4F; #100;
A = 8'hD5; B = 8'h50; #100;
A = 8'hD5; B = 8'h51; #100;
A = 8'hD5; B = 8'h52; #100;
A = 8'hD5; B = 8'h53; #100;
A = 8'hD5; B = 8'h54; #100;
A = 8'hD5; B = 8'h55; #100;
A = 8'hD5; B = 8'h56; #100;
A = 8'hD5; B = 8'h57; #100;
A = 8'hD5; B = 8'h58; #100;
A = 8'hD5; B = 8'h59; #100;
A = 8'hD5; B = 8'h5A; #100;
A = 8'hD5; B = 8'h5B; #100;
A = 8'hD5; B = 8'h5C; #100;
A = 8'hD5; B = 8'h5D; #100;
A = 8'hD5; B = 8'h5E; #100;
A = 8'hD5; B = 8'h5F; #100;
A = 8'hD5; B = 8'h60; #100;
A = 8'hD5; B = 8'h61; #100;
A = 8'hD5; B = 8'h62; #100;
A = 8'hD5; B = 8'h63; #100;
A = 8'hD5; B = 8'h64; #100;
A = 8'hD5; B = 8'h65; #100;
A = 8'hD5; B = 8'h66; #100;
A = 8'hD5; B = 8'h67; #100;
A = 8'hD5; B = 8'h68; #100;
A = 8'hD5; B = 8'h69; #100;
A = 8'hD5; B = 8'h6A; #100;
A = 8'hD5; B = 8'h6B; #100;
A = 8'hD5; B = 8'h6C; #100;
A = 8'hD5; B = 8'h6D; #100;
A = 8'hD5; B = 8'h6E; #100;
A = 8'hD5; B = 8'h6F; #100;
A = 8'hD5; B = 8'h70; #100;
A = 8'hD5; B = 8'h71; #100;
A = 8'hD5; B = 8'h72; #100;
A = 8'hD5; B = 8'h73; #100;
A = 8'hD5; B = 8'h74; #100;
A = 8'hD5; B = 8'h75; #100;
A = 8'hD5; B = 8'h76; #100;
A = 8'hD5; B = 8'h77; #100;
A = 8'hD5; B = 8'h78; #100;
A = 8'hD5; B = 8'h79; #100;
A = 8'hD5; B = 8'h7A; #100;
A = 8'hD5; B = 8'h7B; #100;
A = 8'hD5; B = 8'h7C; #100;
A = 8'hD5; B = 8'h7D; #100;
A = 8'hD5; B = 8'h7E; #100;
A = 8'hD5; B = 8'h7F; #100;
A = 8'hD5; B = 8'h80; #100;
A = 8'hD5; B = 8'h81; #100;
A = 8'hD5; B = 8'h82; #100;
A = 8'hD5; B = 8'h83; #100;
A = 8'hD5; B = 8'h84; #100;
A = 8'hD5; B = 8'h85; #100;
A = 8'hD5; B = 8'h86; #100;
A = 8'hD5; B = 8'h87; #100;
A = 8'hD5; B = 8'h88; #100;
A = 8'hD5; B = 8'h89; #100;
A = 8'hD5; B = 8'h8A; #100;
A = 8'hD5; B = 8'h8B; #100;
A = 8'hD5; B = 8'h8C; #100;
A = 8'hD5; B = 8'h8D; #100;
A = 8'hD5; B = 8'h8E; #100;
A = 8'hD5; B = 8'h8F; #100;
A = 8'hD5; B = 8'h90; #100;
A = 8'hD5; B = 8'h91; #100;
A = 8'hD5; B = 8'h92; #100;
A = 8'hD5; B = 8'h93; #100;
A = 8'hD5; B = 8'h94; #100;
A = 8'hD5; B = 8'h95; #100;
A = 8'hD5; B = 8'h96; #100;
A = 8'hD5; B = 8'h97; #100;
A = 8'hD5; B = 8'h98; #100;
A = 8'hD5; B = 8'h99; #100;
A = 8'hD5; B = 8'h9A; #100;
A = 8'hD5; B = 8'h9B; #100;
A = 8'hD5; B = 8'h9C; #100;
A = 8'hD5; B = 8'h9D; #100;
A = 8'hD5; B = 8'h9E; #100;
A = 8'hD5; B = 8'h9F; #100;
A = 8'hD5; B = 8'hA0; #100;
A = 8'hD5; B = 8'hA1; #100;
A = 8'hD5; B = 8'hA2; #100;
A = 8'hD5; B = 8'hA3; #100;
A = 8'hD5; B = 8'hA4; #100;
A = 8'hD5; B = 8'hA5; #100;
A = 8'hD5; B = 8'hA6; #100;
A = 8'hD5; B = 8'hA7; #100;
A = 8'hD5; B = 8'hA8; #100;
A = 8'hD5; B = 8'hA9; #100;
A = 8'hD5; B = 8'hAA; #100;
A = 8'hD5; B = 8'hAB; #100;
A = 8'hD5; B = 8'hAC; #100;
A = 8'hD5; B = 8'hAD; #100;
A = 8'hD5; B = 8'hAE; #100;
A = 8'hD5; B = 8'hAF; #100;
A = 8'hD5; B = 8'hB0; #100;
A = 8'hD5; B = 8'hB1; #100;
A = 8'hD5; B = 8'hB2; #100;
A = 8'hD5; B = 8'hB3; #100;
A = 8'hD5; B = 8'hB4; #100;
A = 8'hD5; B = 8'hB5; #100;
A = 8'hD5; B = 8'hB6; #100;
A = 8'hD5; B = 8'hB7; #100;
A = 8'hD5; B = 8'hB8; #100;
A = 8'hD5; B = 8'hB9; #100;
A = 8'hD5; B = 8'hBA; #100;
A = 8'hD5; B = 8'hBB; #100;
A = 8'hD5; B = 8'hBC; #100;
A = 8'hD5; B = 8'hBD; #100;
A = 8'hD5; B = 8'hBE; #100;
A = 8'hD5; B = 8'hBF; #100;
A = 8'hD5; B = 8'hC0; #100;
A = 8'hD5; B = 8'hC1; #100;
A = 8'hD5; B = 8'hC2; #100;
A = 8'hD5; B = 8'hC3; #100;
A = 8'hD5; B = 8'hC4; #100;
A = 8'hD5; B = 8'hC5; #100;
A = 8'hD5; B = 8'hC6; #100;
A = 8'hD5; B = 8'hC7; #100;
A = 8'hD5; B = 8'hC8; #100;
A = 8'hD5; B = 8'hC9; #100;
A = 8'hD5; B = 8'hCA; #100;
A = 8'hD5; B = 8'hCB; #100;
A = 8'hD5; B = 8'hCC; #100;
A = 8'hD5; B = 8'hCD; #100;
A = 8'hD5; B = 8'hCE; #100;
A = 8'hD5; B = 8'hCF; #100;
A = 8'hD5; B = 8'hD0; #100;
A = 8'hD5; B = 8'hD1; #100;
A = 8'hD5; B = 8'hD2; #100;
A = 8'hD5; B = 8'hD3; #100;
A = 8'hD5; B = 8'hD4; #100;
A = 8'hD5; B = 8'hD5; #100;
A = 8'hD5; B = 8'hD6; #100;
A = 8'hD5; B = 8'hD7; #100;
A = 8'hD5; B = 8'hD8; #100;
A = 8'hD5; B = 8'hD9; #100;
A = 8'hD5; B = 8'hDA; #100;
A = 8'hD5; B = 8'hDB; #100;
A = 8'hD5; B = 8'hDC; #100;
A = 8'hD5; B = 8'hDD; #100;
A = 8'hD5; B = 8'hDE; #100;
A = 8'hD5; B = 8'hDF; #100;
A = 8'hD5; B = 8'hE0; #100;
A = 8'hD5; B = 8'hE1; #100;
A = 8'hD5; B = 8'hE2; #100;
A = 8'hD5; B = 8'hE3; #100;
A = 8'hD5; B = 8'hE4; #100;
A = 8'hD5; B = 8'hE5; #100;
A = 8'hD5; B = 8'hE6; #100;
A = 8'hD5; B = 8'hE7; #100;
A = 8'hD5; B = 8'hE8; #100;
A = 8'hD5; B = 8'hE9; #100;
A = 8'hD5; B = 8'hEA; #100;
A = 8'hD5; B = 8'hEB; #100;
A = 8'hD5; B = 8'hEC; #100;
A = 8'hD5; B = 8'hED; #100;
A = 8'hD5; B = 8'hEE; #100;
A = 8'hD5; B = 8'hEF; #100;
A = 8'hD5; B = 8'hF0; #100;
A = 8'hD5; B = 8'hF1; #100;
A = 8'hD5; B = 8'hF2; #100;
A = 8'hD5; B = 8'hF3; #100;
A = 8'hD5; B = 8'hF4; #100;
A = 8'hD5; B = 8'hF5; #100;
A = 8'hD5; B = 8'hF6; #100;
A = 8'hD5; B = 8'hF7; #100;
A = 8'hD5; B = 8'hF8; #100;
A = 8'hD5; B = 8'hF9; #100;
A = 8'hD5; B = 8'hFA; #100;
A = 8'hD5; B = 8'hFB; #100;
A = 8'hD5; B = 8'hFC; #100;
A = 8'hD5; B = 8'hFD; #100;
A = 8'hD5; B = 8'hFE; #100;
A = 8'hD5; B = 8'hFF; #100;
A = 8'hD6; B = 8'h0; #100;
A = 8'hD6; B = 8'h1; #100;
A = 8'hD6; B = 8'h2; #100;
A = 8'hD6; B = 8'h3; #100;
A = 8'hD6; B = 8'h4; #100;
A = 8'hD6; B = 8'h5; #100;
A = 8'hD6; B = 8'h6; #100;
A = 8'hD6; B = 8'h7; #100;
A = 8'hD6; B = 8'h8; #100;
A = 8'hD6; B = 8'h9; #100;
A = 8'hD6; B = 8'hA; #100;
A = 8'hD6; B = 8'hB; #100;
A = 8'hD6; B = 8'hC; #100;
A = 8'hD6; B = 8'hD; #100;
A = 8'hD6; B = 8'hE; #100;
A = 8'hD6; B = 8'hF; #100;
A = 8'hD6; B = 8'h10; #100;
A = 8'hD6; B = 8'h11; #100;
A = 8'hD6; B = 8'h12; #100;
A = 8'hD6; B = 8'h13; #100;
A = 8'hD6; B = 8'h14; #100;
A = 8'hD6; B = 8'h15; #100;
A = 8'hD6; B = 8'h16; #100;
A = 8'hD6; B = 8'h17; #100;
A = 8'hD6; B = 8'h18; #100;
A = 8'hD6; B = 8'h19; #100;
A = 8'hD6; B = 8'h1A; #100;
A = 8'hD6; B = 8'h1B; #100;
A = 8'hD6; B = 8'h1C; #100;
A = 8'hD6; B = 8'h1D; #100;
A = 8'hD6; B = 8'h1E; #100;
A = 8'hD6; B = 8'h1F; #100;
A = 8'hD6; B = 8'h20; #100;
A = 8'hD6; B = 8'h21; #100;
A = 8'hD6; B = 8'h22; #100;
A = 8'hD6; B = 8'h23; #100;
A = 8'hD6; B = 8'h24; #100;
A = 8'hD6; B = 8'h25; #100;
A = 8'hD6; B = 8'h26; #100;
A = 8'hD6; B = 8'h27; #100;
A = 8'hD6; B = 8'h28; #100;
A = 8'hD6; B = 8'h29; #100;
A = 8'hD6; B = 8'h2A; #100;
A = 8'hD6; B = 8'h2B; #100;
A = 8'hD6; B = 8'h2C; #100;
A = 8'hD6; B = 8'h2D; #100;
A = 8'hD6; B = 8'h2E; #100;
A = 8'hD6; B = 8'h2F; #100;
A = 8'hD6; B = 8'h30; #100;
A = 8'hD6; B = 8'h31; #100;
A = 8'hD6; B = 8'h32; #100;
A = 8'hD6; B = 8'h33; #100;
A = 8'hD6; B = 8'h34; #100;
A = 8'hD6; B = 8'h35; #100;
A = 8'hD6; B = 8'h36; #100;
A = 8'hD6; B = 8'h37; #100;
A = 8'hD6; B = 8'h38; #100;
A = 8'hD6; B = 8'h39; #100;
A = 8'hD6; B = 8'h3A; #100;
A = 8'hD6; B = 8'h3B; #100;
A = 8'hD6; B = 8'h3C; #100;
A = 8'hD6; B = 8'h3D; #100;
A = 8'hD6; B = 8'h3E; #100;
A = 8'hD6; B = 8'h3F; #100;
A = 8'hD6; B = 8'h40; #100;
A = 8'hD6; B = 8'h41; #100;
A = 8'hD6; B = 8'h42; #100;
A = 8'hD6; B = 8'h43; #100;
A = 8'hD6; B = 8'h44; #100;
A = 8'hD6; B = 8'h45; #100;
A = 8'hD6; B = 8'h46; #100;
A = 8'hD6; B = 8'h47; #100;
A = 8'hD6; B = 8'h48; #100;
A = 8'hD6; B = 8'h49; #100;
A = 8'hD6; B = 8'h4A; #100;
A = 8'hD6; B = 8'h4B; #100;
A = 8'hD6; B = 8'h4C; #100;
A = 8'hD6; B = 8'h4D; #100;
A = 8'hD6; B = 8'h4E; #100;
A = 8'hD6; B = 8'h4F; #100;
A = 8'hD6; B = 8'h50; #100;
A = 8'hD6; B = 8'h51; #100;
A = 8'hD6; B = 8'h52; #100;
A = 8'hD6; B = 8'h53; #100;
A = 8'hD6; B = 8'h54; #100;
A = 8'hD6; B = 8'h55; #100;
A = 8'hD6; B = 8'h56; #100;
A = 8'hD6; B = 8'h57; #100;
A = 8'hD6; B = 8'h58; #100;
A = 8'hD6; B = 8'h59; #100;
A = 8'hD6; B = 8'h5A; #100;
A = 8'hD6; B = 8'h5B; #100;
A = 8'hD6; B = 8'h5C; #100;
A = 8'hD6; B = 8'h5D; #100;
A = 8'hD6; B = 8'h5E; #100;
A = 8'hD6; B = 8'h5F; #100;
A = 8'hD6; B = 8'h60; #100;
A = 8'hD6; B = 8'h61; #100;
A = 8'hD6; B = 8'h62; #100;
A = 8'hD6; B = 8'h63; #100;
A = 8'hD6; B = 8'h64; #100;
A = 8'hD6; B = 8'h65; #100;
A = 8'hD6; B = 8'h66; #100;
A = 8'hD6; B = 8'h67; #100;
A = 8'hD6; B = 8'h68; #100;
A = 8'hD6; B = 8'h69; #100;
A = 8'hD6; B = 8'h6A; #100;
A = 8'hD6; B = 8'h6B; #100;
A = 8'hD6; B = 8'h6C; #100;
A = 8'hD6; B = 8'h6D; #100;
A = 8'hD6; B = 8'h6E; #100;
A = 8'hD6; B = 8'h6F; #100;
A = 8'hD6; B = 8'h70; #100;
A = 8'hD6; B = 8'h71; #100;
A = 8'hD6; B = 8'h72; #100;
A = 8'hD6; B = 8'h73; #100;
A = 8'hD6; B = 8'h74; #100;
A = 8'hD6; B = 8'h75; #100;
A = 8'hD6; B = 8'h76; #100;
A = 8'hD6; B = 8'h77; #100;
A = 8'hD6; B = 8'h78; #100;
A = 8'hD6; B = 8'h79; #100;
A = 8'hD6; B = 8'h7A; #100;
A = 8'hD6; B = 8'h7B; #100;
A = 8'hD6; B = 8'h7C; #100;
A = 8'hD6; B = 8'h7D; #100;
A = 8'hD6; B = 8'h7E; #100;
A = 8'hD6; B = 8'h7F; #100;
A = 8'hD6; B = 8'h80; #100;
A = 8'hD6; B = 8'h81; #100;
A = 8'hD6; B = 8'h82; #100;
A = 8'hD6; B = 8'h83; #100;
A = 8'hD6; B = 8'h84; #100;
A = 8'hD6; B = 8'h85; #100;
A = 8'hD6; B = 8'h86; #100;
A = 8'hD6; B = 8'h87; #100;
A = 8'hD6; B = 8'h88; #100;
A = 8'hD6; B = 8'h89; #100;
A = 8'hD6; B = 8'h8A; #100;
A = 8'hD6; B = 8'h8B; #100;
A = 8'hD6; B = 8'h8C; #100;
A = 8'hD6; B = 8'h8D; #100;
A = 8'hD6; B = 8'h8E; #100;
A = 8'hD6; B = 8'h8F; #100;
A = 8'hD6; B = 8'h90; #100;
A = 8'hD6; B = 8'h91; #100;
A = 8'hD6; B = 8'h92; #100;
A = 8'hD6; B = 8'h93; #100;
A = 8'hD6; B = 8'h94; #100;
A = 8'hD6; B = 8'h95; #100;
A = 8'hD6; B = 8'h96; #100;
A = 8'hD6; B = 8'h97; #100;
A = 8'hD6; B = 8'h98; #100;
A = 8'hD6; B = 8'h99; #100;
A = 8'hD6; B = 8'h9A; #100;
A = 8'hD6; B = 8'h9B; #100;
A = 8'hD6; B = 8'h9C; #100;
A = 8'hD6; B = 8'h9D; #100;
A = 8'hD6; B = 8'h9E; #100;
A = 8'hD6; B = 8'h9F; #100;
A = 8'hD6; B = 8'hA0; #100;
A = 8'hD6; B = 8'hA1; #100;
A = 8'hD6; B = 8'hA2; #100;
A = 8'hD6; B = 8'hA3; #100;
A = 8'hD6; B = 8'hA4; #100;
A = 8'hD6; B = 8'hA5; #100;
A = 8'hD6; B = 8'hA6; #100;
A = 8'hD6; B = 8'hA7; #100;
A = 8'hD6; B = 8'hA8; #100;
A = 8'hD6; B = 8'hA9; #100;
A = 8'hD6; B = 8'hAA; #100;
A = 8'hD6; B = 8'hAB; #100;
A = 8'hD6; B = 8'hAC; #100;
A = 8'hD6; B = 8'hAD; #100;
A = 8'hD6; B = 8'hAE; #100;
A = 8'hD6; B = 8'hAF; #100;
A = 8'hD6; B = 8'hB0; #100;
A = 8'hD6; B = 8'hB1; #100;
A = 8'hD6; B = 8'hB2; #100;
A = 8'hD6; B = 8'hB3; #100;
A = 8'hD6; B = 8'hB4; #100;
A = 8'hD6; B = 8'hB5; #100;
A = 8'hD6; B = 8'hB6; #100;
A = 8'hD6; B = 8'hB7; #100;
A = 8'hD6; B = 8'hB8; #100;
A = 8'hD6; B = 8'hB9; #100;
A = 8'hD6; B = 8'hBA; #100;
A = 8'hD6; B = 8'hBB; #100;
A = 8'hD6; B = 8'hBC; #100;
A = 8'hD6; B = 8'hBD; #100;
A = 8'hD6; B = 8'hBE; #100;
A = 8'hD6; B = 8'hBF; #100;
A = 8'hD6; B = 8'hC0; #100;
A = 8'hD6; B = 8'hC1; #100;
A = 8'hD6; B = 8'hC2; #100;
A = 8'hD6; B = 8'hC3; #100;
A = 8'hD6; B = 8'hC4; #100;
A = 8'hD6; B = 8'hC5; #100;
A = 8'hD6; B = 8'hC6; #100;
A = 8'hD6; B = 8'hC7; #100;
A = 8'hD6; B = 8'hC8; #100;
A = 8'hD6; B = 8'hC9; #100;
A = 8'hD6; B = 8'hCA; #100;
A = 8'hD6; B = 8'hCB; #100;
A = 8'hD6; B = 8'hCC; #100;
A = 8'hD6; B = 8'hCD; #100;
A = 8'hD6; B = 8'hCE; #100;
A = 8'hD6; B = 8'hCF; #100;
A = 8'hD6; B = 8'hD0; #100;
A = 8'hD6; B = 8'hD1; #100;
A = 8'hD6; B = 8'hD2; #100;
A = 8'hD6; B = 8'hD3; #100;
A = 8'hD6; B = 8'hD4; #100;
A = 8'hD6; B = 8'hD5; #100;
A = 8'hD6; B = 8'hD6; #100;
A = 8'hD6; B = 8'hD7; #100;
A = 8'hD6; B = 8'hD8; #100;
A = 8'hD6; B = 8'hD9; #100;
A = 8'hD6; B = 8'hDA; #100;
A = 8'hD6; B = 8'hDB; #100;
A = 8'hD6; B = 8'hDC; #100;
A = 8'hD6; B = 8'hDD; #100;
A = 8'hD6; B = 8'hDE; #100;
A = 8'hD6; B = 8'hDF; #100;
A = 8'hD6; B = 8'hE0; #100;
A = 8'hD6; B = 8'hE1; #100;
A = 8'hD6; B = 8'hE2; #100;
A = 8'hD6; B = 8'hE3; #100;
A = 8'hD6; B = 8'hE4; #100;
A = 8'hD6; B = 8'hE5; #100;
A = 8'hD6; B = 8'hE6; #100;
A = 8'hD6; B = 8'hE7; #100;
A = 8'hD6; B = 8'hE8; #100;
A = 8'hD6; B = 8'hE9; #100;
A = 8'hD6; B = 8'hEA; #100;
A = 8'hD6; B = 8'hEB; #100;
A = 8'hD6; B = 8'hEC; #100;
A = 8'hD6; B = 8'hED; #100;
A = 8'hD6; B = 8'hEE; #100;
A = 8'hD6; B = 8'hEF; #100;
A = 8'hD6; B = 8'hF0; #100;
A = 8'hD6; B = 8'hF1; #100;
A = 8'hD6; B = 8'hF2; #100;
A = 8'hD6; B = 8'hF3; #100;
A = 8'hD6; B = 8'hF4; #100;
A = 8'hD6; B = 8'hF5; #100;
A = 8'hD6; B = 8'hF6; #100;
A = 8'hD6; B = 8'hF7; #100;
A = 8'hD6; B = 8'hF8; #100;
A = 8'hD6; B = 8'hF9; #100;
A = 8'hD6; B = 8'hFA; #100;
A = 8'hD6; B = 8'hFB; #100;
A = 8'hD6; B = 8'hFC; #100;
A = 8'hD6; B = 8'hFD; #100;
A = 8'hD6; B = 8'hFE; #100;
A = 8'hD6; B = 8'hFF; #100;
A = 8'hD7; B = 8'h0; #100;
A = 8'hD7; B = 8'h1; #100;
A = 8'hD7; B = 8'h2; #100;
A = 8'hD7; B = 8'h3; #100;
A = 8'hD7; B = 8'h4; #100;
A = 8'hD7; B = 8'h5; #100;
A = 8'hD7; B = 8'h6; #100;
A = 8'hD7; B = 8'h7; #100;
A = 8'hD7; B = 8'h8; #100;
A = 8'hD7; B = 8'h9; #100;
A = 8'hD7; B = 8'hA; #100;
A = 8'hD7; B = 8'hB; #100;
A = 8'hD7; B = 8'hC; #100;
A = 8'hD7; B = 8'hD; #100;
A = 8'hD7; B = 8'hE; #100;
A = 8'hD7; B = 8'hF; #100;
A = 8'hD7; B = 8'h10; #100;
A = 8'hD7; B = 8'h11; #100;
A = 8'hD7; B = 8'h12; #100;
A = 8'hD7; B = 8'h13; #100;
A = 8'hD7; B = 8'h14; #100;
A = 8'hD7; B = 8'h15; #100;
A = 8'hD7; B = 8'h16; #100;
A = 8'hD7; B = 8'h17; #100;
A = 8'hD7; B = 8'h18; #100;
A = 8'hD7; B = 8'h19; #100;
A = 8'hD7; B = 8'h1A; #100;
A = 8'hD7; B = 8'h1B; #100;
A = 8'hD7; B = 8'h1C; #100;
A = 8'hD7; B = 8'h1D; #100;
A = 8'hD7; B = 8'h1E; #100;
A = 8'hD7; B = 8'h1F; #100;
A = 8'hD7; B = 8'h20; #100;
A = 8'hD7; B = 8'h21; #100;
A = 8'hD7; B = 8'h22; #100;
A = 8'hD7; B = 8'h23; #100;
A = 8'hD7; B = 8'h24; #100;
A = 8'hD7; B = 8'h25; #100;
A = 8'hD7; B = 8'h26; #100;
A = 8'hD7; B = 8'h27; #100;
A = 8'hD7; B = 8'h28; #100;
A = 8'hD7; B = 8'h29; #100;
A = 8'hD7; B = 8'h2A; #100;
A = 8'hD7; B = 8'h2B; #100;
A = 8'hD7; B = 8'h2C; #100;
A = 8'hD7; B = 8'h2D; #100;
A = 8'hD7; B = 8'h2E; #100;
A = 8'hD7; B = 8'h2F; #100;
A = 8'hD7; B = 8'h30; #100;
A = 8'hD7; B = 8'h31; #100;
A = 8'hD7; B = 8'h32; #100;
A = 8'hD7; B = 8'h33; #100;
A = 8'hD7; B = 8'h34; #100;
A = 8'hD7; B = 8'h35; #100;
A = 8'hD7; B = 8'h36; #100;
A = 8'hD7; B = 8'h37; #100;
A = 8'hD7; B = 8'h38; #100;
A = 8'hD7; B = 8'h39; #100;
A = 8'hD7; B = 8'h3A; #100;
A = 8'hD7; B = 8'h3B; #100;
A = 8'hD7; B = 8'h3C; #100;
A = 8'hD7; B = 8'h3D; #100;
A = 8'hD7; B = 8'h3E; #100;
A = 8'hD7; B = 8'h3F; #100;
A = 8'hD7; B = 8'h40; #100;
A = 8'hD7; B = 8'h41; #100;
A = 8'hD7; B = 8'h42; #100;
A = 8'hD7; B = 8'h43; #100;
A = 8'hD7; B = 8'h44; #100;
A = 8'hD7; B = 8'h45; #100;
A = 8'hD7; B = 8'h46; #100;
A = 8'hD7; B = 8'h47; #100;
A = 8'hD7; B = 8'h48; #100;
A = 8'hD7; B = 8'h49; #100;
A = 8'hD7; B = 8'h4A; #100;
A = 8'hD7; B = 8'h4B; #100;
A = 8'hD7; B = 8'h4C; #100;
A = 8'hD7; B = 8'h4D; #100;
A = 8'hD7; B = 8'h4E; #100;
A = 8'hD7; B = 8'h4F; #100;
A = 8'hD7; B = 8'h50; #100;
A = 8'hD7; B = 8'h51; #100;
A = 8'hD7; B = 8'h52; #100;
A = 8'hD7; B = 8'h53; #100;
A = 8'hD7; B = 8'h54; #100;
A = 8'hD7; B = 8'h55; #100;
A = 8'hD7; B = 8'h56; #100;
A = 8'hD7; B = 8'h57; #100;
A = 8'hD7; B = 8'h58; #100;
A = 8'hD7; B = 8'h59; #100;
A = 8'hD7; B = 8'h5A; #100;
A = 8'hD7; B = 8'h5B; #100;
A = 8'hD7; B = 8'h5C; #100;
A = 8'hD7; B = 8'h5D; #100;
A = 8'hD7; B = 8'h5E; #100;
A = 8'hD7; B = 8'h5F; #100;
A = 8'hD7; B = 8'h60; #100;
A = 8'hD7; B = 8'h61; #100;
A = 8'hD7; B = 8'h62; #100;
A = 8'hD7; B = 8'h63; #100;
A = 8'hD7; B = 8'h64; #100;
A = 8'hD7; B = 8'h65; #100;
A = 8'hD7; B = 8'h66; #100;
A = 8'hD7; B = 8'h67; #100;
A = 8'hD7; B = 8'h68; #100;
A = 8'hD7; B = 8'h69; #100;
A = 8'hD7; B = 8'h6A; #100;
A = 8'hD7; B = 8'h6B; #100;
A = 8'hD7; B = 8'h6C; #100;
A = 8'hD7; B = 8'h6D; #100;
A = 8'hD7; B = 8'h6E; #100;
A = 8'hD7; B = 8'h6F; #100;
A = 8'hD7; B = 8'h70; #100;
A = 8'hD7; B = 8'h71; #100;
A = 8'hD7; B = 8'h72; #100;
A = 8'hD7; B = 8'h73; #100;
A = 8'hD7; B = 8'h74; #100;
A = 8'hD7; B = 8'h75; #100;
A = 8'hD7; B = 8'h76; #100;
A = 8'hD7; B = 8'h77; #100;
A = 8'hD7; B = 8'h78; #100;
A = 8'hD7; B = 8'h79; #100;
A = 8'hD7; B = 8'h7A; #100;
A = 8'hD7; B = 8'h7B; #100;
A = 8'hD7; B = 8'h7C; #100;
A = 8'hD7; B = 8'h7D; #100;
A = 8'hD7; B = 8'h7E; #100;
A = 8'hD7; B = 8'h7F; #100;
A = 8'hD7; B = 8'h80; #100;
A = 8'hD7; B = 8'h81; #100;
A = 8'hD7; B = 8'h82; #100;
A = 8'hD7; B = 8'h83; #100;
A = 8'hD7; B = 8'h84; #100;
A = 8'hD7; B = 8'h85; #100;
A = 8'hD7; B = 8'h86; #100;
A = 8'hD7; B = 8'h87; #100;
A = 8'hD7; B = 8'h88; #100;
A = 8'hD7; B = 8'h89; #100;
A = 8'hD7; B = 8'h8A; #100;
A = 8'hD7; B = 8'h8B; #100;
A = 8'hD7; B = 8'h8C; #100;
A = 8'hD7; B = 8'h8D; #100;
A = 8'hD7; B = 8'h8E; #100;
A = 8'hD7; B = 8'h8F; #100;
A = 8'hD7; B = 8'h90; #100;
A = 8'hD7; B = 8'h91; #100;
A = 8'hD7; B = 8'h92; #100;
A = 8'hD7; B = 8'h93; #100;
A = 8'hD7; B = 8'h94; #100;
A = 8'hD7; B = 8'h95; #100;
A = 8'hD7; B = 8'h96; #100;
A = 8'hD7; B = 8'h97; #100;
A = 8'hD7; B = 8'h98; #100;
A = 8'hD7; B = 8'h99; #100;
A = 8'hD7; B = 8'h9A; #100;
A = 8'hD7; B = 8'h9B; #100;
A = 8'hD7; B = 8'h9C; #100;
A = 8'hD7; B = 8'h9D; #100;
A = 8'hD7; B = 8'h9E; #100;
A = 8'hD7; B = 8'h9F; #100;
A = 8'hD7; B = 8'hA0; #100;
A = 8'hD7; B = 8'hA1; #100;
A = 8'hD7; B = 8'hA2; #100;
A = 8'hD7; B = 8'hA3; #100;
A = 8'hD7; B = 8'hA4; #100;
A = 8'hD7; B = 8'hA5; #100;
A = 8'hD7; B = 8'hA6; #100;
A = 8'hD7; B = 8'hA7; #100;
A = 8'hD7; B = 8'hA8; #100;
A = 8'hD7; B = 8'hA9; #100;
A = 8'hD7; B = 8'hAA; #100;
A = 8'hD7; B = 8'hAB; #100;
A = 8'hD7; B = 8'hAC; #100;
A = 8'hD7; B = 8'hAD; #100;
A = 8'hD7; B = 8'hAE; #100;
A = 8'hD7; B = 8'hAF; #100;
A = 8'hD7; B = 8'hB0; #100;
A = 8'hD7; B = 8'hB1; #100;
A = 8'hD7; B = 8'hB2; #100;
A = 8'hD7; B = 8'hB3; #100;
A = 8'hD7; B = 8'hB4; #100;
A = 8'hD7; B = 8'hB5; #100;
A = 8'hD7; B = 8'hB6; #100;
A = 8'hD7; B = 8'hB7; #100;
A = 8'hD7; B = 8'hB8; #100;
A = 8'hD7; B = 8'hB9; #100;
A = 8'hD7; B = 8'hBA; #100;
A = 8'hD7; B = 8'hBB; #100;
A = 8'hD7; B = 8'hBC; #100;
A = 8'hD7; B = 8'hBD; #100;
A = 8'hD7; B = 8'hBE; #100;
A = 8'hD7; B = 8'hBF; #100;
A = 8'hD7; B = 8'hC0; #100;
A = 8'hD7; B = 8'hC1; #100;
A = 8'hD7; B = 8'hC2; #100;
A = 8'hD7; B = 8'hC3; #100;
A = 8'hD7; B = 8'hC4; #100;
A = 8'hD7; B = 8'hC5; #100;
A = 8'hD7; B = 8'hC6; #100;
A = 8'hD7; B = 8'hC7; #100;
A = 8'hD7; B = 8'hC8; #100;
A = 8'hD7; B = 8'hC9; #100;
A = 8'hD7; B = 8'hCA; #100;
A = 8'hD7; B = 8'hCB; #100;
A = 8'hD7; B = 8'hCC; #100;
A = 8'hD7; B = 8'hCD; #100;
A = 8'hD7; B = 8'hCE; #100;
A = 8'hD7; B = 8'hCF; #100;
A = 8'hD7; B = 8'hD0; #100;
A = 8'hD7; B = 8'hD1; #100;
A = 8'hD7; B = 8'hD2; #100;
A = 8'hD7; B = 8'hD3; #100;
A = 8'hD7; B = 8'hD4; #100;
A = 8'hD7; B = 8'hD5; #100;
A = 8'hD7; B = 8'hD6; #100;
A = 8'hD7; B = 8'hD7; #100;
A = 8'hD7; B = 8'hD8; #100;
A = 8'hD7; B = 8'hD9; #100;
A = 8'hD7; B = 8'hDA; #100;
A = 8'hD7; B = 8'hDB; #100;
A = 8'hD7; B = 8'hDC; #100;
A = 8'hD7; B = 8'hDD; #100;
A = 8'hD7; B = 8'hDE; #100;
A = 8'hD7; B = 8'hDF; #100;
A = 8'hD7; B = 8'hE0; #100;
A = 8'hD7; B = 8'hE1; #100;
A = 8'hD7; B = 8'hE2; #100;
A = 8'hD7; B = 8'hE3; #100;
A = 8'hD7; B = 8'hE4; #100;
A = 8'hD7; B = 8'hE5; #100;
A = 8'hD7; B = 8'hE6; #100;
A = 8'hD7; B = 8'hE7; #100;
A = 8'hD7; B = 8'hE8; #100;
A = 8'hD7; B = 8'hE9; #100;
A = 8'hD7; B = 8'hEA; #100;
A = 8'hD7; B = 8'hEB; #100;
A = 8'hD7; B = 8'hEC; #100;
A = 8'hD7; B = 8'hED; #100;
A = 8'hD7; B = 8'hEE; #100;
A = 8'hD7; B = 8'hEF; #100;
A = 8'hD7; B = 8'hF0; #100;
A = 8'hD7; B = 8'hF1; #100;
A = 8'hD7; B = 8'hF2; #100;
A = 8'hD7; B = 8'hF3; #100;
A = 8'hD7; B = 8'hF4; #100;
A = 8'hD7; B = 8'hF5; #100;
A = 8'hD7; B = 8'hF6; #100;
A = 8'hD7; B = 8'hF7; #100;
A = 8'hD7; B = 8'hF8; #100;
A = 8'hD7; B = 8'hF9; #100;
A = 8'hD7; B = 8'hFA; #100;
A = 8'hD7; B = 8'hFB; #100;
A = 8'hD7; B = 8'hFC; #100;
A = 8'hD7; B = 8'hFD; #100;
A = 8'hD7; B = 8'hFE; #100;
A = 8'hD7; B = 8'hFF; #100;
A = 8'hD8; B = 8'h0; #100;
A = 8'hD8; B = 8'h1; #100;
A = 8'hD8; B = 8'h2; #100;
A = 8'hD8; B = 8'h3; #100;
A = 8'hD8; B = 8'h4; #100;
A = 8'hD8; B = 8'h5; #100;
A = 8'hD8; B = 8'h6; #100;
A = 8'hD8; B = 8'h7; #100;
A = 8'hD8; B = 8'h8; #100;
A = 8'hD8; B = 8'h9; #100;
A = 8'hD8; B = 8'hA; #100;
A = 8'hD8; B = 8'hB; #100;
A = 8'hD8; B = 8'hC; #100;
A = 8'hD8; B = 8'hD; #100;
A = 8'hD8; B = 8'hE; #100;
A = 8'hD8; B = 8'hF; #100;
A = 8'hD8; B = 8'h10; #100;
A = 8'hD8; B = 8'h11; #100;
A = 8'hD8; B = 8'h12; #100;
A = 8'hD8; B = 8'h13; #100;
A = 8'hD8; B = 8'h14; #100;
A = 8'hD8; B = 8'h15; #100;
A = 8'hD8; B = 8'h16; #100;
A = 8'hD8; B = 8'h17; #100;
A = 8'hD8; B = 8'h18; #100;
A = 8'hD8; B = 8'h19; #100;
A = 8'hD8; B = 8'h1A; #100;
A = 8'hD8; B = 8'h1B; #100;
A = 8'hD8; B = 8'h1C; #100;
A = 8'hD8; B = 8'h1D; #100;
A = 8'hD8; B = 8'h1E; #100;
A = 8'hD8; B = 8'h1F; #100;
A = 8'hD8; B = 8'h20; #100;
A = 8'hD8; B = 8'h21; #100;
A = 8'hD8; B = 8'h22; #100;
A = 8'hD8; B = 8'h23; #100;
A = 8'hD8; B = 8'h24; #100;
A = 8'hD8; B = 8'h25; #100;
A = 8'hD8; B = 8'h26; #100;
A = 8'hD8; B = 8'h27; #100;
A = 8'hD8; B = 8'h28; #100;
A = 8'hD8; B = 8'h29; #100;
A = 8'hD8; B = 8'h2A; #100;
A = 8'hD8; B = 8'h2B; #100;
A = 8'hD8; B = 8'h2C; #100;
A = 8'hD8; B = 8'h2D; #100;
A = 8'hD8; B = 8'h2E; #100;
A = 8'hD8; B = 8'h2F; #100;
A = 8'hD8; B = 8'h30; #100;
A = 8'hD8; B = 8'h31; #100;
A = 8'hD8; B = 8'h32; #100;
A = 8'hD8; B = 8'h33; #100;
A = 8'hD8; B = 8'h34; #100;
A = 8'hD8; B = 8'h35; #100;
A = 8'hD8; B = 8'h36; #100;
A = 8'hD8; B = 8'h37; #100;
A = 8'hD8; B = 8'h38; #100;
A = 8'hD8; B = 8'h39; #100;
A = 8'hD8; B = 8'h3A; #100;
A = 8'hD8; B = 8'h3B; #100;
A = 8'hD8; B = 8'h3C; #100;
A = 8'hD8; B = 8'h3D; #100;
A = 8'hD8; B = 8'h3E; #100;
A = 8'hD8; B = 8'h3F; #100;
A = 8'hD8; B = 8'h40; #100;
A = 8'hD8; B = 8'h41; #100;
A = 8'hD8; B = 8'h42; #100;
A = 8'hD8; B = 8'h43; #100;
A = 8'hD8; B = 8'h44; #100;
A = 8'hD8; B = 8'h45; #100;
A = 8'hD8; B = 8'h46; #100;
A = 8'hD8; B = 8'h47; #100;
A = 8'hD8; B = 8'h48; #100;
A = 8'hD8; B = 8'h49; #100;
A = 8'hD8; B = 8'h4A; #100;
A = 8'hD8; B = 8'h4B; #100;
A = 8'hD8; B = 8'h4C; #100;
A = 8'hD8; B = 8'h4D; #100;
A = 8'hD8; B = 8'h4E; #100;
A = 8'hD8; B = 8'h4F; #100;
A = 8'hD8; B = 8'h50; #100;
A = 8'hD8; B = 8'h51; #100;
A = 8'hD8; B = 8'h52; #100;
A = 8'hD8; B = 8'h53; #100;
A = 8'hD8; B = 8'h54; #100;
A = 8'hD8; B = 8'h55; #100;
A = 8'hD8; B = 8'h56; #100;
A = 8'hD8; B = 8'h57; #100;
A = 8'hD8; B = 8'h58; #100;
A = 8'hD8; B = 8'h59; #100;
A = 8'hD8; B = 8'h5A; #100;
A = 8'hD8; B = 8'h5B; #100;
A = 8'hD8; B = 8'h5C; #100;
A = 8'hD8; B = 8'h5D; #100;
A = 8'hD8; B = 8'h5E; #100;
A = 8'hD8; B = 8'h5F; #100;
A = 8'hD8; B = 8'h60; #100;
A = 8'hD8; B = 8'h61; #100;
A = 8'hD8; B = 8'h62; #100;
A = 8'hD8; B = 8'h63; #100;
A = 8'hD8; B = 8'h64; #100;
A = 8'hD8; B = 8'h65; #100;
A = 8'hD8; B = 8'h66; #100;
A = 8'hD8; B = 8'h67; #100;
A = 8'hD8; B = 8'h68; #100;
A = 8'hD8; B = 8'h69; #100;
A = 8'hD8; B = 8'h6A; #100;
A = 8'hD8; B = 8'h6B; #100;
A = 8'hD8; B = 8'h6C; #100;
A = 8'hD8; B = 8'h6D; #100;
A = 8'hD8; B = 8'h6E; #100;
A = 8'hD8; B = 8'h6F; #100;
A = 8'hD8; B = 8'h70; #100;
A = 8'hD8; B = 8'h71; #100;
A = 8'hD8; B = 8'h72; #100;
A = 8'hD8; B = 8'h73; #100;
A = 8'hD8; B = 8'h74; #100;
A = 8'hD8; B = 8'h75; #100;
A = 8'hD8; B = 8'h76; #100;
A = 8'hD8; B = 8'h77; #100;
A = 8'hD8; B = 8'h78; #100;
A = 8'hD8; B = 8'h79; #100;
A = 8'hD8; B = 8'h7A; #100;
A = 8'hD8; B = 8'h7B; #100;
A = 8'hD8; B = 8'h7C; #100;
A = 8'hD8; B = 8'h7D; #100;
A = 8'hD8; B = 8'h7E; #100;
A = 8'hD8; B = 8'h7F; #100;
A = 8'hD8; B = 8'h80; #100;
A = 8'hD8; B = 8'h81; #100;
A = 8'hD8; B = 8'h82; #100;
A = 8'hD8; B = 8'h83; #100;
A = 8'hD8; B = 8'h84; #100;
A = 8'hD8; B = 8'h85; #100;
A = 8'hD8; B = 8'h86; #100;
A = 8'hD8; B = 8'h87; #100;
A = 8'hD8; B = 8'h88; #100;
A = 8'hD8; B = 8'h89; #100;
A = 8'hD8; B = 8'h8A; #100;
A = 8'hD8; B = 8'h8B; #100;
A = 8'hD8; B = 8'h8C; #100;
A = 8'hD8; B = 8'h8D; #100;
A = 8'hD8; B = 8'h8E; #100;
A = 8'hD8; B = 8'h8F; #100;
A = 8'hD8; B = 8'h90; #100;
A = 8'hD8; B = 8'h91; #100;
A = 8'hD8; B = 8'h92; #100;
A = 8'hD8; B = 8'h93; #100;
A = 8'hD8; B = 8'h94; #100;
A = 8'hD8; B = 8'h95; #100;
A = 8'hD8; B = 8'h96; #100;
A = 8'hD8; B = 8'h97; #100;
A = 8'hD8; B = 8'h98; #100;
A = 8'hD8; B = 8'h99; #100;
A = 8'hD8; B = 8'h9A; #100;
A = 8'hD8; B = 8'h9B; #100;
A = 8'hD8; B = 8'h9C; #100;
A = 8'hD8; B = 8'h9D; #100;
A = 8'hD8; B = 8'h9E; #100;
A = 8'hD8; B = 8'h9F; #100;
A = 8'hD8; B = 8'hA0; #100;
A = 8'hD8; B = 8'hA1; #100;
A = 8'hD8; B = 8'hA2; #100;
A = 8'hD8; B = 8'hA3; #100;
A = 8'hD8; B = 8'hA4; #100;
A = 8'hD8; B = 8'hA5; #100;
A = 8'hD8; B = 8'hA6; #100;
A = 8'hD8; B = 8'hA7; #100;
A = 8'hD8; B = 8'hA8; #100;
A = 8'hD8; B = 8'hA9; #100;
A = 8'hD8; B = 8'hAA; #100;
A = 8'hD8; B = 8'hAB; #100;
A = 8'hD8; B = 8'hAC; #100;
A = 8'hD8; B = 8'hAD; #100;
A = 8'hD8; B = 8'hAE; #100;
A = 8'hD8; B = 8'hAF; #100;
A = 8'hD8; B = 8'hB0; #100;
A = 8'hD8; B = 8'hB1; #100;
A = 8'hD8; B = 8'hB2; #100;
A = 8'hD8; B = 8'hB3; #100;
A = 8'hD8; B = 8'hB4; #100;
A = 8'hD8; B = 8'hB5; #100;
A = 8'hD8; B = 8'hB6; #100;
A = 8'hD8; B = 8'hB7; #100;
A = 8'hD8; B = 8'hB8; #100;
A = 8'hD8; B = 8'hB9; #100;
A = 8'hD8; B = 8'hBA; #100;
A = 8'hD8; B = 8'hBB; #100;
A = 8'hD8; B = 8'hBC; #100;
A = 8'hD8; B = 8'hBD; #100;
A = 8'hD8; B = 8'hBE; #100;
A = 8'hD8; B = 8'hBF; #100;
A = 8'hD8; B = 8'hC0; #100;
A = 8'hD8; B = 8'hC1; #100;
A = 8'hD8; B = 8'hC2; #100;
A = 8'hD8; B = 8'hC3; #100;
A = 8'hD8; B = 8'hC4; #100;
A = 8'hD8; B = 8'hC5; #100;
A = 8'hD8; B = 8'hC6; #100;
A = 8'hD8; B = 8'hC7; #100;
A = 8'hD8; B = 8'hC8; #100;
A = 8'hD8; B = 8'hC9; #100;
A = 8'hD8; B = 8'hCA; #100;
A = 8'hD8; B = 8'hCB; #100;
A = 8'hD8; B = 8'hCC; #100;
A = 8'hD8; B = 8'hCD; #100;
A = 8'hD8; B = 8'hCE; #100;
A = 8'hD8; B = 8'hCF; #100;
A = 8'hD8; B = 8'hD0; #100;
A = 8'hD8; B = 8'hD1; #100;
A = 8'hD8; B = 8'hD2; #100;
A = 8'hD8; B = 8'hD3; #100;
A = 8'hD8; B = 8'hD4; #100;
A = 8'hD8; B = 8'hD5; #100;
A = 8'hD8; B = 8'hD6; #100;
A = 8'hD8; B = 8'hD7; #100;
A = 8'hD8; B = 8'hD8; #100;
A = 8'hD8; B = 8'hD9; #100;
A = 8'hD8; B = 8'hDA; #100;
A = 8'hD8; B = 8'hDB; #100;
A = 8'hD8; B = 8'hDC; #100;
A = 8'hD8; B = 8'hDD; #100;
A = 8'hD8; B = 8'hDE; #100;
A = 8'hD8; B = 8'hDF; #100;
A = 8'hD8; B = 8'hE0; #100;
A = 8'hD8; B = 8'hE1; #100;
A = 8'hD8; B = 8'hE2; #100;
A = 8'hD8; B = 8'hE3; #100;
A = 8'hD8; B = 8'hE4; #100;
A = 8'hD8; B = 8'hE5; #100;
A = 8'hD8; B = 8'hE6; #100;
A = 8'hD8; B = 8'hE7; #100;
A = 8'hD8; B = 8'hE8; #100;
A = 8'hD8; B = 8'hE9; #100;
A = 8'hD8; B = 8'hEA; #100;
A = 8'hD8; B = 8'hEB; #100;
A = 8'hD8; B = 8'hEC; #100;
A = 8'hD8; B = 8'hED; #100;
A = 8'hD8; B = 8'hEE; #100;
A = 8'hD8; B = 8'hEF; #100;
A = 8'hD8; B = 8'hF0; #100;
A = 8'hD8; B = 8'hF1; #100;
A = 8'hD8; B = 8'hF2; #100;
A = 8'hD8; B = 8'hF3; #100;
A = 8'hD8; B = 8'hF4; #100;
A = 8'hD8; B = 8'hF5; #100;
A = 8'hD8; B = 8'hF6; #100;
A = 8'hD8; B = 8'hF7; #100;
A = 8'hD8; B = 8'hF8; #100;
A = 8'hD8; B = 8'hF9; #100;
A = 8'hD8; B = 8'hFA; #100;
A = 8'hD8; B = 8'hFB; #100;
A = 8'hD8; B = 8'hFC; #100;
A = 8'hD8; B = 8'hFD; #100;
A = 8'hD8; B = 8'hFE; #100;
A = 8'hD8; B = 8'hFF; #100;
A = 8'hD9; B = 8'h0; #100;
A = 8'hD9; B = 8'h1; #100;
A = 8'hD9; B = 8'h2; #100;
A = 8'hD9; B = 8'h3; #100;
A = 8'hD9; B = 8'h4; #100;
A = 8'hD9; B = 8'h5; #100;
A = 8'hD9; B = 8'h6; #100;
A = 8'hD9; B = 8'h7; #100;
A = 8'hD9; B = 8'h8; #100;
A = 8'hD9; B = 8'h9; #100;
A = 8'hD9; B = 8'hA; #100;
A = 8'hD9; B = 8'hB; #100;
A = 8'hD9; B = 8'hC; #100;
A = 8'hD9; B = 8'hD; #100;
A = 8'hD9; B = 8'hE; #100;
A = 8'hD9; B = 8'hF; #100;
A = 8'hD9; B = 8'h10; #100;
A = 8'hD9; B = 8'h11; #100;
A = 8'hD9; B = 8'h12; #100;
A = 8'hD9; B = 8'h13; #100;
A = 8'hD9; B = 8'h14; #100;
A = 8'hD9; B = 8'h15; #100;
A = 8'hD9; B = 8'h16; #100;
A = 8'hD9; B = 8'h17; #100;
A = 8'hD9; B = 8'h18; #100;
A = 8'hD9; B = 8'h19; #100;
A = 8'hD9; B = 8'h1A; #100;
A = 8'hD9; B = 8'h1B; #100;
A = 8'hD9; B = 8'h1C; #100;
A = 8'hD9; B = 8'h1D; #100;
A = 8'hD9; B = 8'h1E; #100;
A = 8'hD9; B = 8'h1F; #100;
A = 8'hD9; B = 8'h20; #100;
A = 8'hD9; B = 8'h21; #100;
A = 8'hD9; B = 8'h22; #100;
A = 8'hD9; B = 8'h23; #100;
A = 8'hD9; B = 8'h24; #100;
A = 8'hD9; B = 8'h25; #100;
A = 8'hD9; B = 8'h26; #100;
A = 8'hD9; B = 8'h27; #100;
A = 8'hD9; B = 8'h28; #100;
A = 8'hD9; B = 8'h29; #100;
A = 8'hD9; B = 8'h2A; #100;
A = 8'hD9; B = 8'h2B; #100;
A = 8'hD9; B = 8'h2C; #100;
A = 8'hD9; B = 8'h2D; #100;
A = 8'hD9; B = 8'h2E; #100;
A = 8'hD9; B = 8'h2F; #100;
A = 8'hD9; B = 8'h30; #100;
A = 8'hD9; B = 8'h31; #100;
A = 8'hD9; B = 8'h32; #100;
A = 8'hD9; B = 8'h33; #100;
A = 8'hD9; B = 8'h34; #100;
A = 8'hD9; B = 8'h35; #100;
A = 8'hD9; B = 8'h36; #100;
A = 8'hD9; B = 8'h37; #100;
A = 8'hD9; B = 8'h38; #100;
A = 8'hD9; B = 8'h39; #100;
A = 8'hD9; B = 8'h3A; #100;
A = 8'hD9; B = 8'h3B; #100;
A = 8'hD9; B = 8'h3C; #100;
A = 8'hD9; B = 8'h3D; #100;
A = 8'hD9; B = 8'h3E; #100;
A = 8'hD9; B = 8'h3F; #100;
A = 8'hD9; B = 8'h40; #100;
A = 8'hD9; B = 8'h41; #100;
A = 8'hD9; B = 8'h42; #100;
A = 8'hD9; B = 8'h43; #100;
A = 8'hD9; B = 8'h44; #100;
A = 8'hD9; B = 8'h45; #100;
A = 8'hD9; B = 8'h46; #100;
A = 8'hD9; B = 8'h47; #100;
A = 8'hD9; B = 8'h48; #100;
A = 8'hD9; B = 8'h49; #100;
A = 8'hD9; B = 8'h4A; #100;
A = 8'hD9; B = 8'h4B; #100;
A = 8'hD9; B = 8'h4C; #100;
A = 8'hD9; B = 8'h4D; #100;
A = 8'hD9; B = 8'h4E; #100;
A = 8'hD9; B = 8'h4F; #100;
A = 8'hD9; B = 8'h50; #100;
A = 8'hD9; B = 8'h51; #100;
A = 8'hD9; B = 8'h52; #100;
A = 8'hD9; B = 8'h53; #100;
A = 8'hD9; B = 8'h54; #100;
A = 8'hD9; B = 8'h55; #100;
A = 8'hD9; B = 8'h56; #100;
A = 8'hD9; B = 8'h57; #100;
A = 8'hD9; B = 8'h58; #100;
A = 8'hD9; B = 8'h59; #100;
A = 8'hD9; B = 8'h5A; #100;
A = 8'hD9; B = 8'h5B; #100;
A = 8'hD9; B = 8'h5C; #100;
A = 8'hD9; B = 8'h5D; #100;
A = 8'hD9; B = 8'h5E; #100;
A = 8'hD9; B = 8'h5F; #100;
A = 8'hD9; B = 8'h60; #100;
A = 8'hD9; B = 8'h61; #100;
A = 8'hD9; B = 8'h62; #100;
A = 8'hD9; B = 8'h63; #100;
A = 8'hD9; B = 8'h64; #100;
A = 8'hD9; B = 8'h65; #100;
A = 8'hD9; B = 8'h66; #100;
A = 8'hD9; B = 8'h67; #100;
A = 8'hD9; B = 8'h68; #100;
A = 8'hD9; B = 8'h69; #100;
A = 8'hD9; B = 8'h6A; #100;
A = 8'hD9; B = 8'h6B; #100;
A = 8'hD9; B = 8'h6C; #100;
A = 8'hD9; B = 8'h6D; #100;
A = 8'hD9; B = 8'h6E; #100;
A = 8'hD9; B = 8'h6F; #100;
A = 8'hD9; B = 8'h70; #100;
A = 8'hD9; B = 8'h71; #100;
A = 8'hD9; B = 8'h72; #100;
A = 8'hD9; B = 8'h73; #100;
A = 8'hD9; B = 8'h74; #100;
A = 8'hD9; B = 8'h75; #100;
A = 8'hD9; B = 8'h76; #100;
A = 8'hD9; B = 8'h77; #100;
A = 8'hD9; B = 8'h78; #100;
A = 8'hD9; B = 8'h79; #100;
A = 8'hD9; B = 8'h7A; #100;
A = 8'hD9; B = 8'h7B; #100;
A = 8'hD9; B = 8'h7C; #100;
A = 8'hD9; B = 8'h7D; #100;
A = 8'hD9; B = 8'h7E; #100;
A = 8'hD9; B = 8'h7F; #100;
A = 8'hD9; B = 8'h80; #100;
A = 8'hD9; B = 8'h81; #100;
A = 8'hD9; B = 8'h82; #100;
A = 8'hD9; B = 8'h83; #100;
A = 8'hD9; B = 8'h84; #100;
A = 8'hD9; B = 8'h85; #100;
A = 8'hD9; B = 8'h86; #100;
A = 8'hD9; B = 8'h87; #100;
A = 8'hD9; B = 8'h88; #100;
A = 8'hD9; B = 8'h89; #100;
A = 8'hD9; B = 8'h8A; #100;
A = 8'hD9; B = 8'h8B; #100;
A = 8'hD9; B = 8'h8C; #100;
A = 8'hD9; B = 8'h8D; #100;
A = 8'hD9; B = 8'h8E; #100;
A = 8'hD9; B = 8'h8F; #100;
A = 8'hD9; B = 8'h90; #100;
A = 8'hD9; B = 8'h91; #100;
A = 8'hD9; B = 8'h92; #100;
A = 8'hD9; B = 8'h93; #100;
A = 8'hD9; B = 8'h94; #100;
A = 8'hD9; B = 8'h95; #100;
A = 8'hD9; B = 8'h96; #100;
A = 8'hD9; B = 8'h97; #100;
A = 8'hD9; B = 8'h98; #100;
A = 8'hD9; B = 8'h99; #100;
A = 8'hD9; B = 8'h9A; #100;
A = 8'hD9; B = 8'h9B; #100;
A = 8'hD9; B = 8'h9C; #100;
A = 8'hD9; B = 8'h9D; #100;
A = 8'hD9; B = 8'h9E; #100;
A = 8'hD9; B = 8'h9F; #100;
A = 8'hD9; B = 8'hA0; #100;
A = 8'hD9; B = 8'hA1; #100;
A = 8'hD9; B = 8'hA2; #100;
A = 8'hD9; B = 8'hA3; #100;
A = 8'hD9; B = 8'hA4; #100;
A = 8'hD9; B = 8'hA5; #100;
A = 8'hD9; B = 8'hA6; #100;
A = 8'hD9; B = 8'hA7; #100;
A = 8'hD9; B = 8'hA8; #100;
A = 8'hD9; B = 8'hA9; #100;
A = 8'hD9; B = 8'hAA; #100;
A = 8'hD9; B = 8'hAB; #100;
A = 8'hD9; B = 8'hAC; #100;
A = 8'hD9; B = 8'hAD; #100;
A = 8'hD9; B = 8'hAE; #100;
A = 8'hD9; B = 8'hAF; #100;
A = 8'hD9; B = 8'hB0; #100;
A = 8'hD9; B = 8'hB1; #100;
A = 8'hD9; B = 8'hB2; #100;
A = 8'hD9; B = 8'hB3; #100;
A = 8'hD9; B = 8'hB4; #100;
A = 8'hD9; B = 8'hB5; #100;
A = 8'hD9; B = 8'hB6; #100;
A = 8'hD9; B = 8'hB7; #100;
A = 8'hD9; B = 8'hB8; #100;
A = 8'hD9; B = 8'hB9; #100;
A = 8'hD9; B = 8'hBA; #100;
A = 8'hD9; B = 8'hBB; #100;
A = 8'hD9; B = 8'hBC; #100;
A = 8'hD9; B = 8'hBD; #100;
A = 8'hD9; B = 8'hBE; #100;
A = 8'hD9; B = 8'hBF; #100;
A = 8'hD9; B = 8'hC0; #100;
A = 8'hD9; B = 8'hC1; #100;
A = 8'hD9; B = 8'hC2; #100;
A = 8'hD9; B = 8'hC3; #100;
A = 8'hD9; B = 8'hC4; #100;
A = 8'hD9; B = 8'hC5; #100;
A = 8'hD9; B = 8'hC6; #100;
A = 8'hD9; B = 8'hC7; #100;
A = 8'hD9; B = 8'hC8; #100;
A = 8'hD9; B = 8'hC9; #100;
A = 8'hD9; B = 8'hCA; #100;
A = 8'hD9; B = 8'hCB; #100;
A = 8'hD9; B = 8'hCC; #100;
A = 8'hD9; B = 8'hCD; #100;
A = 8'hD9; B = 8'hCE; #100;
A = 8'hD9; B = 8'hCF; #100;
A = 8'hD9; B = 8'hD0; #100;
A = 8'hD9; B = 8'hD1; #100;
A = 8'hD9; B = 8'hD2; #100;
A = 8'hD9; B = 8'hD3; #100;
A = 8'hD9; B = 8'hD4; #100;
A = 8'hD9; B = 8'hD5; #100;
A = 8'hD9; B = 8'hD6; #100;
A = 8'hD9; B = 8'hD7; #100;
A = 8'hD9; B = 8'hD8; #100;
A = 8'hD9; B = 8'hD9; #100;
A = 8'hD9; B = 8'hDA; #100;
A = 8'hD9; B = 8'hDB; #100;
A = 8'hD9; B = 8'hDC; #100;
A = 8'hD9; B = 8'hDD; #100;
A = 8'hD9; B = 8'hDE; #100;
A = 8'hD9; B = 8'hDF; #100;
A = 8'hD9; B = 8'hE0; #100;
A = 8'hD9; B = 8'hE1; #100;
A = 8'hD9; B = 8'hE2; #100;
A = 8'hD9; B = 8'hE3; #100;
A = 8'hD9; B = 8'hE4; #100;
A = 8'hD9; B = 8'hE5; #100;
A = 8'hD9; B = 8'hE6; #100;
A = 8'hD9; B = 8'hE7; #100;
A = 8'hD9; B = 8'hE8; #100;
A = 8'hD9; B = 8'hE9; #100;
A = 8'hD9; B = 8'hEA; #100;
A = 8'hD9; B = 8'hEB; #100;
A = 8'hD9; B = 8'hEC; #100;
A = 8'hD9; B = 8'hED; #100;
A = 8'hD9; B = 8'hEE; #100;
A = 8'hD9; B = 8'hEF; #100;
A = 8'hD9; B = 8'hF0; #100;
A = 8'hD9; B = 8'hF1; #100;
A = 8'hD9; B = 8'hF2; #100;
A = 8'hD9; B = 8'hF3; #100;
A = 8'hD9; B = 8'hF4; #100;
A = 8'hD9; B = 8'hF5; #100;
A = 8'hD9; B = 8'hF6; #100;
A = 8'hD9; B = 8'hF7; #100;
A = 8'hD9; B = 8'hF8; #100;
A = 8'hD9; B = 8'hF9; #100;
A = 8'hD9; B = 8'hFA; #100;
A = 8'hD9; B = 8'hFB; #100;
A = 8'hD9; B = 8'hFC; #100;
A = 8'hD9; B = 8'hFD; #100;
A = 8'hD9; B = 8'hFE; #100;
A = 8'hD9; B = 8'hFF; #100;
A = 8'hDA; B = 8'h0; #100;
A = 8'hDA; B = 8'h1; #100;
A = 8'hDA; B = 8'h2; #100;
A = 8'hDA; B = 8'h3; #100;
A = 8'hDA; B = 8'h4; #100;
A = 8'hDA; B = 8'h5; #100;
A = 8'hDA; B = 8'h6; #100;
A = 8'hDA; B = 8'h7; #100;
A = 8'hDA; B = 8'h8; #100;
A = 8'hDA; B = 8'h9; #100;
A = 8'hDA; B = 8'hA; #100;
A = 8'hDA; B = 8'hB; #100;
A = 8'hDA; B = 8'hC; #100;
A = 8'hDA; B = 8'hD; #100;
A = 8'hDA; B = 8'hE; #100;
A = 8'hDA; B = 8'hF; #100;
A = 8'hDA; B = 8'h10; #100;
A = 8'hDA; B = 8'h11; #100;
A = 8'hDA; B = 8'h12; #100;
A = 8'hDA; B = 8'h13; #100;
A = 8'hDA; B = 8'h14; #100;
A = 8'hDA; B = 8'h15; #100;
A = 8'hDA; B = 8'h16; #100;
A = 8'hDA; B = 8'h17; #100;
A = 8'hDA; B = 8'h18; #100;
A = 8'hDA; B = 8'h19; #100;
A = 8'hDA; B = 8'h1A; #100;
A = 8'hDA; B = 8'h1B; #100;
A = 8'hDA; B = 8'h1C; #100;
A = 8'hDA; B = 8'h1D; #100;
A = 8'hDA; B = 8'h1E; #100;
A = 8'hDA; B = 8'h1F; #100;
A = 8'hDA; B = 8'h20; #100;
A = 8'hDA; B = 8'h21; #100;
A = 8'hDA; B = 8'h22; #100;
A = 8'hDA; B = 8'h23; #100;
A = 8'hDA; B = 8'h24; #100;
A = 8'hDA; B = 8'h25; #100;
A = 8'hDA; B = 8'h26; #100;
A = 8'hDA; B = 8'h27; #100;
A = 8'hDA; B = 8'h28; #100;
A = 8'hDA; B = 8'h29; #100;
A = 8'hDA; B = 8'h2A; #100;
A = 8'hDA; B = 8'h2B; #100;
A = 8'hDA; B = 8'h2C; #100;
A = 8'hDA; B = 8'h2D; #100;
A = 8'hDA; B = 8'h2E; #100;
A = 8'hDA; B = 8'h2F; #100;
A = 8'hDA; B = 8'h30; #100;
A = 8'hDA; B = 8'h31; #100;
A = 8'hDA; B = 8'h32; #100;
A = 8'hDA; B = 8'h33; #100;
A = 8'hDA; B = 8'h34; #100;
A = 8'hDA; B = 8'h35; #100;
A = 8'hDA; B = 8'h36; #100;
A = 8'hDA; B = 8'h37; #100;
A = 8'hDA; B = 8'h38; #100;
A = 8'hDA; B = 8'h39; #100;
A = 8'hDA; B = 8'h3A; #100;
A = 8'hDA; B = 8'h3B; #100;
A = 8'hDA; B = 8'h3C; #100;
A = 8'hDA; B = 8'h3D; #100;
A = 8'hDA; B = 8'h3E; #100;
A = 8'hDA; B = 8'h3F; #100;
A = 8'hDA; B = 8'h40; #100;
A = 8'hDA; B = 8'h41; #100;
A = 8'hDA; B = 8'h42; #100;
A = 8'hDA; B = 8'h43; #100;
A = 8'hDA; B = 8'h44; #100;
A = 8'hDA; B = 8'h45; #100;
A = 8'hDA; B = 8'h46; #100;
A = 8'hDA; B = 8'h47; #100;
A = 8'hDA; B = 8'h48; #100;
A = 8'hDA; B = 8'h49; #100;
A = 8'hDA; B = 8'h4A; #100;
A = 8'hDA; B = 8'h4B; #100;
A = 8'hDA; B = 8'h4C; #100;
A = 8'hDA; B = 8'h4D; #100;
A = 8'hDA; B = 8'h4E; #100;
A = 8'hDA; B = 8'h4F; #100;
A = 8'hDA; B = 8'h50; #100;
A = 8'hDA; B = 8'h51; #100;
A = 8'hDA; B = 8'h52; #100;
A = 8'hDA; B = 8'h53; #100;
A = 8'hDA; B = 8'h54; #100;
A = 8'hDA; B = 8'h55; #100;
A = 8'hDA; B = 8'h56; #100;
A = 8'hDA; B = 8'h57; #100;
A = 8'hDA; B = 8'h58; #100;
A = 8'hDA; B = 8'h59; #100;
A = 8'hDA; B = 8'h5A; #100;
A = 8'hDA; B = 8'h5B; #100;
A = 8'hDA; B = 8'h5C; #100;
A = 8'hDA; B = 8'h5D; #100;
A = 8'hDA; B = 8'h5E; #100;
A = 8'hDA; B = 8'h5F; #100;
A = 8'hDA; B = 8'h60; #100;
A = 8'hDA; B = 8'h61; #100;
A = 8'hDA; B = 8'h62; #100;
A = 8'hDA; B = 8'h63; #100;
A = 8'hDA; B = 8'h64; #100;
A = 8'hDA; B = 8'h65; #100;
A = 8'hDA; B = 8'h66; #100;
A = 8'hDA; B = 8'h67; #100;
A = 8'hDA; B = 8'h68; #100;
A = 8'hDA; B = 8'h69; #100;
A = 8'hDA; B = 8'h6A; #100;
A = 8'hDA; B = 8'h6B; #100;
A = 8'hDA; B = 8'h6C; #100;
A = 8'hDA; B = 8'h6D; #100;
A = 8'hDA; B = 8'h6E; #100;
A = 8'hDA; B = 8'h6F; #100;
A = 8'hDA; B = 8'h70; #100;
A = 8'hDA; B = 8'h71; #100;
A = 8'hDA; B = 8'h72; #100;
A = 8'hDA; B = 8'h73; #100;
A = 8'hDA; B = 8'h74; #100;
A = 8'hDA; B = 8'h75; #100;
A = 8'hDA; B = 8'h76; #100;
A = 8'hDA; B = 8'h77; #100;
A = 8'hDA; B = 8'h78; #100;
A = 8'hDA; B = 8'h79; #100;
A = 8'hDA; B = 8'h7A; #100;
A = 8'hDA; B = 8'h7B; #100;
A = 8'hDA; B = 8'h7C; #100;
A = 8'hDA; B = 8'h7D; #100;
A = 8'hDA; B = 8'h7E; #100;
A = 8'hDA; B = 8'h7F; #100;
A = 8'hDA; B = 8'h80; #100;
A = 8'hDA; B = 8'h81; #100;
A = 8'hDA; B = 8'h82; #100;
A = 8'hDA; B = 8'h83; #100;
A = 8'hDA; B = 8'h84; #100;
A = 8'hDA; B = 8'h85; #100;
A = 8'hDA; B = 8'h86; #100;
A = 8'hDA; B = 8'h87; #100;
A = 8'hDA; B = 8'h88; #100;
A = 8'hDA; B = 8'h89; #100;
A = 8'hDA; B = 8'h8A; #100;
A = 8'hDA; B = 8'h8B; #100;
A = 8'hDA; B = 8'h8C; #100;
A = 8'hDA; B = 8'h8D; #100;
A = 8'hDA; B = 8'h8E; #100;
A = 8'hDA; B = 8'h8F; #100;
A = 8'hDA; B = 8'h90; #100;
A = 8'hDA; B = 8'h91; #100;
A = 8'hDA; B = 8'h92; #100;
A = 8'hDA; B = 8'h93; #100;
A = 8'hDA; B = 8'h94; #100;
A = 8'hDA; B = 8'h95; #100;
A = 8'hDA; B = 8'h96; #100;
A = 8'hDA; B = 8'h97; #100;
A = 8'hDA; B = 8'h98; #100;
A = 8'hDA; B = 8'h99; #100;
A = 8'hDA; B = 8'h9A; #100;
A = 8'hDA; B = 8'h9B; #100;
A = 8'hDA; B = 8'h9C; #100;
A = 8'hDA; B = 8'h9D; #100;
A = 8'hDA; B = 8'h9E; #100;
A = 8'hDA; B = 8'h9F; #100;
A = 8'hDA; B = 8'hA0; #100;
A = 8'hDA; B = 8'hA1; #100;
A = 8'hDA; B = 8'hA2; #100;
A = 8'hDA; B = 8'hA3; #100;
A = 8'hDA; B = 8'hA4; #100;
A = 8'hDA; B = 8'hA5; #100;
A = 8'hDA; B = 8'hA6; #100;
A = 8'hDA; B = 8'hA7; #100;
A = 8'hDA; B = 8'hA8; #100;
A = 8'hDA; B = 8'hA9; #100;
A = 8'hDA; B = 8'hAA; #100;
A = 8'hDA; B = 8'hAB; #100;
A = 8'hDA; B = 8'hAC; #100;
A = 8'hDA; B = 8'hAD; #100;
A = 8'hDA; B = 8'hAE; #100;
A = 8'hDA; B = 8'hAF; #100;
A = 8'hDA; B = 8'hB0; #100;
A = 8'hDA; B = 8'hB1; #100;
A = 8'hDA; B = 8'hB2; #100;
A = 8'hDA; B = 8'hB3; #100;
A = 8'hDA; B = 8'hB4; #100;
A = 8'hDA; B = 8'hB5; #100;
A = 8'hDA; B = 8'hB6; #100;
A = 8'hDA; B = 8'hB7; #100;
A = 8'hDA; B = 8'hB8; #100;
A = 8'hDA; B = 8'hB9; #100;
A = 8'hDA; B = 8'hBA; #100;
A = 8'hDA; B = 8'hBB; #100;
A = 8'hDA; B = 8'hBC; #100;
A = 8'hDA; B = 8'hBD; #100;
A = 8'hDA; B = 8'hBE; #100;
A = 8'hDA; B = 8'hBF; #100;
A = 8'hDA; B = 8'hC0; #100;
A = 8'hDA; B = 8'hC1; #100;
A = 8'hDA; B = 8'hC2; #100;
A = 8'hDA; B = 8'hC3; #100;
A = 8'hDA; B = 8'hC4; #100;
A = 8'hDA; B = 8'hC5; #100;
A = 8'hDA; B = 8'hC6; #100;
A = 8'hDA; B = 8'hC7; #100;
A = 8'hDA; B = 8'hC8; #100;
A = 8'hDA; B = 8'hC9; #100;
A = 8'hDA; B = 8'hCA; #100;
A = 8'hDA; B = 8'hCB; #100;
A = 8'hDA; B = 8'hCC; #100;
A = 8'hDA; B = 8'hCD; #100;
A = 8'hDA; B = 8'hCE; #100;
A = 8'hDA; B = 8'hCF; #100;
A = 8'hDA; B = 8'hD0; #100;
A = 8'hDA; B = 8'hD1; #100;
A = 8'hDA; B = 8'hD2; #100;
A = 8'hDA; B = 8'hD3; #100;
A = 8'hDA; B = 8'hD4; #100;
A = 8'hDA; B = 8'hD5; #100;
A = 8'hDA; B = 8'hD6; #100;
A = 8'hDA; B = 8'hD7; #100;
A = 8'hDA; B = 8'hD8; #100;
A = 8'hDA; B = 8'hD9; #100;
A = 8'hDA; B = 8'hDA; #100;
A = 8'hDA; B = 8'hDB; #100;
A = 8'hDA; B = 8'hDC; #100;
A = 8'hDA; B = 8'hDD; #100;
A = 8'hDA; B = 8'hDE; #100;
A = 8'hDA; B = 8'hDF; #100;
A = 8'hDA; B = 8'hE0; #100;
A = 8'hDA; B = 8'hE1; #100;
A = 8'hDA; B = 8'hE2; #100;
A = 8'hDA; B = 8'hE3; #100;
A = 8'hDA; B = 8'hE4; #100;
A = 8'hDA; B = 8'hE5; #100;
A = 8'hDA; B = 8'hE6; #100;
A = 8'hDA; B = 8'hE7; #100;
A = 8'hDA; B = 8'hE8; #100;
A = 8'hDA; B = 8'hE9; #100;
A = 8'hDA; B = 8'hEA; #100;
A = 8'hDA; B = 8'hEB; #100;
A = 8'hDA; B = 8'hEC; #100;
A = 8'hDA; B = 8'hED; #100;
A = 8'hDA; B = 8'hEE; #100;
A = 8'hDA; B = 8'hEF; #100;
A = 8'hDA; B = 8'hF0; #100;
A = 8'hDA; B = 8'hF1; #100;
A = 8'hDA; B = 8'hF2; #100;
A = 8'hDA; B = 8'hF3; #100;
A = 8'hDA; B = 8'hF4; #100;
A = 8'hDA; B = 8'hF5; #100;
A = 8'hDA; B = 8'hF6; #100;
A = 8'hDA; B = 8'hF7; #100;
A = 8'hDA; B = 8'hF8; #100;
A = 8'hDA; B = 8'hF9; #100;
A = 8'hDA; B = 8'hFA; #100;
A = 8'hDA; B = 8'hFB; #100;
A = 8'hDA; B = 8'hFC; #100;
A = 8'hDA; B = 8'hFD; #100;
A = 8'hDA; B = 8'hFE; #100;
A = 8'hDA; B = 8'hFF; #100;
A = 8'hDB; B = 8'h0; #100;
A = 8'hDB; B = 8'h1; #100;
A = 8'hDB; B = 8'h2; #100;
A = 8'hDB; B = 8'h3; #100;
A = 8'hDB; B = 8'h4; #100;
A = 8'hDB; B = 8'h5; #100;
A = 8'hDB; B = 8'h6; #100;
A = 8'hDB; B = 8'h7; #100;
A = 8'hDB; B = 8'h8; #100;
A = 8'hDB; B = 8'h9; #100;
A = 8'hDB; B = 8'hA; #100;
A = 8'hDB; B = 8'hB; #100;
A = 8'hDB; B = 8'hC; #100;
A = 8'hDB; B = 8'hD; #100;
A = 8'hDB; B = 8'hE; #100;
A = 8'hDB; B = 8'hF; #100;
A = 8'hDB; B = 8'h10; #100;
A = 8'hDB; B = 8'h11; #100;
A = 8'hDB; B = 8'h12; #100;
A = 8'hDB; B = 8'h13; #100;
A = 8'hDB; B = 8'h14; #100;
A = 8'hDB; B = 8'h15; #100;
A = 8'hDB; B = 8'h16; #100;
A = 8'hDB; B = 8'h17; #100;
A = 8'hDB; B = 8'h18; #100;
A = 8'hDB; B = 8'h19; #100;
A = 8'hDB; B = 8'h1A; #100;
A = 8'hDB; B = 8'h1B; #100;
A = 8'hDB; B = 8'h1C; #100;
A = 8'hDB; B = 8'h1D; #100;
A = 8'hDB; B = 8'h1E; #100;
A = 8'hDB; B = 8'h1F; #100;
A = 8'hDB; B = 8'h20; #100;
A = 8'hDB; B = 8'h21; #100;
A = 8'hDB; B = 8'h22; #100;
A = 8'hDB; B = 8'h23; #100;
A = 8'hDB; B = 8'h24; #100;
A = 8'hDB; B = 8'h25; #100;
A = 8'hDB; B = 8'h26; #100;
A = 8'hDB; B = 8'h27; #100;
A = 8'hDB; B = 8'h28; #100;
A = 8'hDB; B = 8'h29; #100;
A = 8'hDB; B = 8'h2A; #100;
A = 8'hDB; B = 8'h2B; #100;
A = 8'hDB; B = 8'h2C; #100;
A = 8'hDB; B = 8'h2D; #100;
A = 8'hDB; B = 8'h2E; #100;
A = 8'hDB; B = 8'h2F; #100;
A = 8'hDB; B = 8'h30; #100;
A = 8'hDB; B = 8'h31; #100;
A = 8'hDB; B = 8'h32; #100;
A = 8'hDB; B = 8'h33; #100;
A = 8'hDB; B = 8'h34; #100;
A = 8'hDB; B = 8'h35; #100;
A = 8'hDB; B = 8'h36; #100;
A = 8'hDB; B = 8'h37; #100;
A = 8'hDB; B = 8'h38; #100;
A = 8'hDB; B = 8'h39; #100;
A = 8'hDB; B = 8'h3A; #100;
A = 8'hDB; B = 8'h3B; #100;
A = 8'hDB; B = 8'h3C; #100;
A = 8'hDB; B = 8'h3D; #100;
A = 8'hDB; B = 8'h3E; #100;
A = 8'hDB; B = 8'h3F; #100;
A = 8'hDB; B = 8'h40; #100;
A = 8'hDB; B = 8'h41; #100;
A = 8'hDB; B = 8'h42; #100;
A = 8'hDB; B = 8'h43; #100;
A = 8'hDB; B = 8'h44; #100;
A = 8'hDB; B = 8'h45; #100;
A = 8'hDB; B = 8'h46; #100;
A = 8'hDB; B = 8'h47; #100;
A = 8'hDB; B = 8'h48; #100;
A = 8'hDB; B = 8'h49; #100;
A = 8'hDB; B = 8'h4A; #100;
A = 8'hDB; B = 8'h4B; #100;
A = 8'hDB; B = 8'h4C; #100;
A = 8'hDB; B = 8'h4D; #100;
A = 8'hDB; B = 8'h4E; #100;
A = 8'hDB; B = 8'h4F; #100;
A = 8'hDB; B = 8'h50; #100;
A = 8'hDB; B = 8'h51; #100;
A = 8'hDB; B = 8'h52; #100;
A = 8'hDB; B = 8'h53; #100;
A = 8'hDB; B = 8'h54; #100;
A = 8'hDB; B = 8'h55; #100;
A = 8'hDB; B = 8'h56; #100;
A = 8'hDB; B = 8'h57; #100;
A = 8'hDB; B = 8'h58; #100;
A = 8'hDB; B = 8'h59; #100;
A = 8'hDB; B = 8'h5A; #100;
A = 8'hDB; B = 8'h5B; #100;
A = 8'hDB; B = 8'h5C; #100;
A = 8'hDB; B = 8'h5D; #100;
A = 8'hDB; B = 8'h5E; #100;
A = 8'hDB; B = 8'h5F; #100;
A = 8'hDB; B = 8'h60; #100;
A = 8'hDB; B = 8'h61; #100;
A = 8'hDB; B = 8'h62; #100;
A = 8'hDB; B = 8'h63; #100;
A = 8'hDB; B = 8'h64; #100;
A = 8'hDB; B = 8'h65; #100;
A = 8'hDB; B = 8'h66; #100;
A = 8'hDB; B = 8'h67; #100;
A = 8'hDB; B = 8'h68; #100;
A = 8'hDB; B = 8'h69; #100;
A = 8'hDB; B = 8'h6A; #100;
A = 8'hDB; B = 8'h6B; #100;
A = 8'hDB; B = 8'h6C; #100;
A = 8'hDB; B = 8'h6D; #100;
A = 8'hDB; B = 8'h6E; #100;
A = 8'hDB; B = 8'h6F; #100;
A = 8'hDB; B = 8'h70; #100;
A = 8'hDB; B = 8'h71; #100;
A = 8'hDB; B = 8'h72; #100;
A = 8'hDB; B = 8'h73; #100;
A = 8'hDB; B = 8'h74; #100;
A = 8'hDB; B = 8'h75; #100;
A = 8'hDB; B = 8'h76; #100;
A = 8'hDB; B = 8'h77; #100;
A = 8'hDB; B = 8'h78; #100;
A = 8'hDB; B = 8'h79; #100;
A = 8'hDB; B = 8'h7A; #100;
A = 8'hDB; B = 8'h7B; #100;
A = 8'hDB; B = 8'h7C; #100;
A = 8'hDB; B = 8'h7D; #100;
A = 8'hDB; B = 8'h7E; #100;
A = 8'hDB; B = 8'h7F; #100;
A = 8'hDB; B = 8'h80; #100;
A = 8'hDB; B = 8'h81; #100;
A = 8'hDB; B = 8'h82; #100;
A = 8'hDB; B = 8'h83; #100;
A = 8'hDB; B = 8'h84; #100;
A = 8'hDB; B = 8'h85; #100;
A = 8'hDB; B = 8'h86; #100;
A = 8'hDB; B = 8'h87; #100;
A = 8'hDB; B = 8'h88; #100;
A = 8'hDB; B = 8'h89; #100;
A = 8'hDB; B = 8'h8A; #100;
A = 8'hDB; B = 8'h8B; #100;
A = 8'hDB; B = 8'h8C; #100;
A = 8'hDB; B = 8'h8D; #100;
A = 8'hDB; B = 8'h8E; #100;
A = 8'hDB; B = 8'h8F; #100;
A = 8'hDB; B = 8'h90; #100;
A = 8'hDB; B = 8'h91; #100;
A = 8'hDB; B = 8'h92; #100;
A = 8'hDB; B = 8'h93; #100;
A = 8'hDB; B = 8'h94; #100;
A = 8'hDB; B = 8'h95; #100;
A = 8'hDB; B = 8'h96; #100;
A = 8'hDB; B = 8'h97; #100;
A = 8'hDB; B = 8'h98; #100;
A = 8'hDB; B = 8'h99; #100;
A = 8'hDB; B = 8'h9A; #100;
A = 8'hDB; B = 8'h9B; #100;
A = 8'hDB; B = 8'h9C; #100;
A = 8'hDB; B = 8'h9D; #100;
A = 8'hDB; B = 8'h9E; #100;
A = 8'hDB; B = 8'h9F; #100;
A = 8'hDB; B = 8'hA0; #100;
A = 8'hDB; B = 8'hA1; #100;
A = 8'hDB; B = 8'hA2; #100;
A = 8'hDB; B = 8'hA3; #100;
A = 8'hDB; B = 8'hA4; #100;
A = 8'hDB; B = 8'hA5; #100;
A = 8'hDB; B = 8'hA6; #100;
A = 8'hDB; B = 8'hA7; #100;
A = 8'hDB; B = 8'hA8; #100;
A = 8'hDB; B = 8'hA9; #100;
A = 8'hDB; B = 8'hAA; #100;
A = 8'hDB; B = 8'hAB; #100;
A = 8'hDB; B = 8'hAC; #100;
A = 8'hDB; B = 8'hAD; #100;
A = 8'hDB; B = 8'hAE; #100;
A = 8'hDB; B = 8'hAF; #100;
A = 8'hDB; B = 8'hB0; #100;
A = 8'hDB; B = 8'hB1; #100;
A = 8'hDB; B = 8'hB2; #100;
A = 8'hDB; B = 8'hB3; #100;
A = 8'hDB; B = 8'hB4; #100;
A = 8'hDB; B = 8'hB5; #100;
A = 8'hDB; B = 8'hB6; #100;
A = 8'hDB; B = 8'hB7; #100;
A = 8'hDB; B = 8'hB8; #100;
A = 8'hDB; B = 8'hB9; #100;
A = 8'hDB; B = 8'hBA; #100;
A = 8'hDB; B = 8'hBB; #100;
A = 8'hDB; B = 8'hBC; #100;
A = 8'hDB; B = 8'hBD; #100;
A = 8'hDB; B = 8'hBE; #100;
A = 8'hDB; B = 8'hBF; #100;
A = 8'hDB; B = 8'hC0; #100;
A = 8'hDB; B = 8'hC1; #100;
A = 8'hDB; B = 8'hC2; #100;
A = 8'hDB; B = 8'hC3; #100;
A = 8'hDB; B = 8'hC4; #100;
A = 8'hDB; B = 8'hC5; #100;
A = 8'hDB; B = 8'hC6; #100;
A = 8'hDB; B = 8'hC7; #100;
A = 8'hDB; B = 8'hC8; #100;
A = 8'hDB; B = 8'hC9; #100;
A = 8'hDB; B = 8'hCA; #100;
A = 8'hDB; B = 8'hCB; #100;
A = 8'hDB; B = 8'hCC; #100;
A = 8'hDB; B = 8'hCD; #100;
A = 8'hDB; B = 8'hCE; #100;
A = 8'hDB; B = 8'hCF; #100;
A = 8'hDB; B = 8'hD0; #100;
A = 8'hDB; B = 8'hD1; #100;
A = 8'hDB; B = 8'hD2; #100;
A = 8'hDB; B = 8'hD3; #100;
A = 8'hDB; B = 8'hD4; #100;
A = 8'hDB; B = 8'hD5; #100;
A = 8'hDB; B = 8'hD6; #100;
A = 8'hDB; B = 8'hD7; #100;
A = 8'hDB; B = 8'hD8; #100;
A = 8'hDB; B = 8'hD9; #100;
A = 8'hDB; B = 8'hDA; #100;
A = 8'hDB; B = 8'hDB; #100;
A = 8'hDB; B = 8'hDC; #100;
A = 8'hDB; B = 8'hDD; #100;
A = 8'hDB; B = 8'hDE; #100;
A = 8'hDB; B = 8'hDF; #100;
A = 8'hDB; B = 8'hE0; #100;
A = 8'hDB; B = 8'hE1; #100;
A = 8'hDB; B = 8'hE2; #100;
A = 8'hDB; B = 8'hE3; #100;
A = 8'hDB; B = 8'hE4; #100;
A = 8'hDB; B = 8'hE5; #100;
A = 8'hDB; B = 8'hE6; #100;
A = 8'hDB; B = 8'hE7; #100;
A = 8'hDB; B = 8'hE8; #100;
A = 8'hDB; B = 8'hE9; #100;
A = 8'hDB; B = 8'hEA; #100;
A = 8'hDB; B = 8'hEB; #100;
A = 8'hDB; B = 8'hEC; #100;
A = 8'hDB; B = 8'hED; #100;
A = 8'hDB; B = 8'hEE; #100;
A = 8'hDB; B = 8'hEF; #100;
A = 8'hDB; B = 8'hF0; #100;
A = 8'hDB; B = 8'hF1; #100;
A = 8'hDB; B = 8'hF2; #100;
A = 8'hDB; B = 8'hF3; #100;
A = 8'hDB; B = 8'hF4; #100;
A = 8'hDB; B = 8'hF5; #100;
A = 8'hDB; B = 8'hF6; #100;
A = 8'hDB; B = 8'hF7; #100;
A = 8'hDB; B = 8'hF8; #100;
A = 8'hDB; B = 8'hF9; #100;
A = 8'hDB; B = 8'hFA; #100;
A = 8'hDB; B = 8'hFB; #100;
A = 8'hDB; B = 8'hFC; #100;
A = 8'hDB; B = 8'hFD; #100;
A = 8'hDB; B = 8'hFE; #100;
A = 8'hDB; B = 8'hFF; #100;
A = 8'hDC; B = 8'h0; #100;
A = 8'hDC; B = 8'h1; #100;
A = 8'hDC; B = 8'h2; #100;
A = 8'hDC; B = 8'h3; #100;
A = 8'hDC; B = 8'h4; #100;
A = 8'hDC; B = 8'h5; #100;
A = 8'hDC; B = 8'h6; #100;
A = 8'hDC; B = 8'h7; #100;
A = 8'hDC; B = 8'h8; #100;
A = 8'hDC; B = 8'h9; #100;
A = 8'hDC; B = 8'hA; #100;
A = 8'hDC; B = 8'hB; #100;
A = 8'hDC; B = 8'hC; #100;
A = 8'hDC; B = 8'hD; #100;
A = 8'hDC; B = 8'hE; #100;
A = 8'hDC; B = 8'hF; #100;
A = 8'hDC; B = 8'h10; #100;
A = 8'hDC; B = 8'h11; #100;
A = 8'hDC; B = 8'h12; #100;
A = 8'hDC; B = 8'h13; #100;
A = 8'hDC; B = 8'h14; #100;
A = 8'hDC; B = 8'h15; #100;
A = 8'hDC; B = 8'h16; #100;
A = 8'hDC; B = 8'h17; #100;
A = 8'hDC; B = 8'h18; #100;
A = 8'hDC; B = 8'h19; #100;
A = 8'hDC; B = 8'h1A; #100;
A = 8'hDC; B = 8'h1B; #100;
A = 8'hDC; B = 8'h1C; #100;
A = 8'hDC; B = 8'h1D; #100;
A = 8'hDC; B = 8'h1E; #100;
A = 8'hDC; B = 8'h1F; #100;
A = 8'hDC; B = 8'h20; #100;
A = 8'hDC; B = 8'h21; #100;
A = 8'hDC; B = 8'h22; #100;
A = 8'hDC; B = 8'h23; #100;
A = 8'hDC; B = 8'h24; #100;
A = 8'hDC; B = 8'h25; #100;
A = 8'hDC; B = 8'h26; #100;
A = 8'hDC; B = 8'h27; #100;
A = 8'hDC; B = 8'h28; #100;
A = 8'hDC; B = 8'h29; #100;
A = 8'hDC; B = 8'h2A; #100;
A = 8'hDC; B = 8'h2B; #100;
A = 8'hDC; B = 8'h2C; #100;
A = 8'hDC; B = 8'h2D; #100;
A = 8'hDC; B = 8'h2E; #100;
A = 8'hDC; B = 8'h2F; #100;
A = 8'hDC; B = 8'h30; #100;
A = 8'hDC; B = 8'h31; #100;
A = 8'hDC; B = 8'h32; #100;
A = 8'hDC; B = 8'h33; #100;
A = 8'hDC; B = 8'h34; #100;
A = 8'hDC; B = 8'h35; #100;
A = 8'hDC; B = 8'h36; #100;
A = 8'hDC; B = 8'h37; #100;
A = 8'hDC; B = 8'h38; #100;
A = 8'hDC; B = 8'h39; #100;
A = 8'hDC; B = 8'h3A; #100;
A = 8'hDC; B = 8'h3B; #100;
A = 8'hDC; B = 8'h3C; #100;
A = 8'hDC; B = 8'h3D; #100;
A = 8'hDC; B = 8'h3E; #100;
A = 8'hDC; B = 8'h3F; #100;
A = 8'hDC; B = 8'h40; #100;
A = 8'hDC; B = 8'h41; #100;
A = 8'hDC; B = 8'h42; #100;
A = 8'hDC; B = 8'h43; #100;
A = 8'hDC; B = 8'h44; #100;
A = 8'hDC; B = 8'h45; #100;
A = 8'hDC; B = 8'h46; #100;
A = 8'hDC; B = 8'h47; #100;
A = 8'hDC; B = 8'h48; #100;
A = 8'hDC; B = 8'h49; #100;
A = 8'hDC; B = 8'h4A; #100;
A = 8'hDC; B = 8'h4B; #100;
A = 8'hDC; B = 8'h4C; #100;
A = 8'hDC; B = 8'h4D; #100;
A = 8'hDC; B = 8'h4E; #100;
A = 8'hDC; B = 8'h4F; #100;
A = 8'hDC; B = 8'h50; #100;
A = 8'hDC; B = 8'h51; #100;
A = 8'hDC; B = 8'h52; #100;
A = 8'hDC; B = 8'h53; #100;
A = 8'hDC; B = 8'h54; #100;
A = 8'hDC; B = 8'h55; #100;
A = 8'hDC; B = 8'h56; #100;
A = 8'hDC; B = 8'h57; #100;
A = 8'hDC; B = 8'h58; #100;
A = 8'hDC; B = 8'h59; #100;
A = 8'hDC; B = 8'h5A; #100;
A = 8'hDC; B = 8'h5B; #100;
A = 8'hDC; B = 8'h5C; #100;
A = 8'hDC; B = 8'h5D; #100;
A = 8'hDC; B = 8'h5E; #100;
A = 8'hDC; B = 8'h5F; #100;
A = 8'hDC; B = 8'h60; #100;
A = 8'hDC; B = 8'h61; #100;
A = 8'hDC; B = 8'h62; #100;
A = 8'hDC; B = 8'h63; #100;
A = 8'hDC; B = 8'h64; #100;
A = 8'hDC; B = 8'h65; #100;
A = 8'hDC; B = 8'h66; #100;
A = 8'hDC; B = 8'h67; #100;
A = 8'hDC; B = 8'h68; #100;
A = 8'hDC; B = 8'h69; #100;
A = 8'hDC; B = 8'h6A; #100;
A = 8'hDC; B = 8'h6B; #100;
A = 8'hDC; B = 8'h6C; #100;
A = 8'hDC; B = 8'h6D; #100;
A = 8'hDC; B = 8'h6E; #100;
A = 8'hDC; B = 8'h6F; #100;
A = 8'hDC; B = 8'h70; #100;
A = 8'hDC; B = 8'h71; #100;
A = 8'hDC; B = 8'h72; #100;
A = 8'hDC; B = 8'h73; #100;
A = 8'hDC; B = 8'h74; #100;
A = 8'hDC; B = 8'h75; #100;
A = 8'hDC; B = 8'h76; #100;
A = 8'hDC; B = 8'h77; #100;
A = 8'hDC; B = 8'h78; #100;
A = 8'hDC; B = 8'h79; #100;
A = 8'hDC; B = 8'h7A; #100;
A = 8'hDC; B = 8'h7B; #100;
A = 8'hDC; B = 8'h7C; #100;
A = 8'hDC; B = 8'h7D; #100;
A = 8'hDC; B = 8'h7E; #100;
A = 8'hDC; B = 8'h7F; #100;
A = 8'hDC; B = 8'h80; #100;
A = 8'hDC; B = 8'h81; #100;
A = 8'hDC; B = 8'h82; #100;
A = 8'hDC; B = 8'h83; #100;
A = 8'hDC; B = 8'h84; #100;
A = 8'hDC; B = 8'h85; #100;
A = 8'hDC; B = 8'h86; #100;
A = 8'hDC; B = 8'h87; #100;
A = 8'hDC; B = 8'h88; #100;
A = 8'hDC; B = 8'h89; #100;
A = 8'hDC; B = 8'h8A; #100;
A = 8'hDC; B = 8'h8B; #100;
A = 8'hDC; B = 8'h8C; #100;
A = 8'hDC; B = 8'h8D; #100;
A = 8'hDC; B = 8'h8E; #100;
A = 8'hDC; B = 8'h8F; #100;
A = 8'hDC; B = 8'h90; #100;
A = 8'hDC; B = 8'h91; #100;
A = 8'hDC; B = 8'h92; #100;
A = 8'hDC; B = 8'h93; #100;
A = 8'hDC; B = 8'h94; #100;
A = 8'hDC; B = 8'h95; #100;
A = 8'hDC; B = 8'h96; #100;
A = 8'hDC; B = 8'h97; #100;
A = 8'hDC; B = 8'h98; #100;
A = 8'hDC; B = 8'h99; #100;
A = 8'hDC; B = 8'h9A; #100;
A = 8'hDC; B = 8'h9B; #100;
A = 8'hDC; B = 8'h9C; #100;
A = 8'hDC; B = 8'h9D; #100;
A = 8'hDC; B = 8'h9E; #100;
A = 8'hDC; B = 8'h9F; #100;
A = 8'hDC; B = 8'hA0; #100;
A = 8'hDC; B = 8'hA1; #100;
A = 8'hDC; B = 8'hA2; #100;
A = 8'hDC; B = 8'hA3; #100;
A = 8'hDC; B = 8'hA4; #100;
A = 8'hDC; B = 8'hA5; #100;
A = 8'hDC; B = 8'hA6; #100;
A = 8'hDC; B = 8'hA7; #100;
A = 8'hDC; B = 8'hA8; #100;
A = 8'hDC; B = 8'hA9; #100;
A = 8'hDC; B = 8'hAA; #100;
A = 8'hDC; B = 8'hAB; #100;
A = 8'hDC; B = 8'hAC; #100;
A = 8'hDC; B = 8'hAD; #100;
A = 8'hDC; B = 8'hAE; #100;
A = 8'hDC; B = 8'hAF; #100;
A = 8'hDC; B = 8'hB0; #100;
A = 8'hDC; B = 8'hB1; #100;
A = 8'hDC; B = 8'hB2; #100;
A = 8'hDC; B = 8'hB3; #100;
A = 8'hDC; B = 8'hB4; #100;
A = 8'hDC; B = 8'hB5; #100;
A = 8'hDC; B = 8'hB6; #100;
A = 8'hDC; B = 8'hB7; #100;
A = 8'hDC; B = 8'hB8; #100;
A = 8'hDC; B = 8'hB9; #100;
A = 8'hDC; B = 8'hBA; #100;
A = 8'hDC; B = 8'hBB; #100;
A = 8'hDC; B = 8'hBC; #100;
A = 8'hDC; B = 8'hBD; #100;
A = 8'hDC; B = 8'hBE; #100;
A = 8'hDC; B = 8'hBF; #100;
A = 8'hDC; B = 8'hC0; #100;
A = 8'hDC; B = 8'hC1; #100;
A = 8'hDC; B = 8'hC2; #100;
A = 8'hDC; B = 8'hC3; #100;
A = 8'hDC; B = 8'hC4; #100;
A = 8'hDC; B = 8'hC5; #100;
A = 8'hDC; B = 8'hC6; #100;
A = 8'hDC; B = 8'hC7; #100;
A = 8'hDC; B = 8'hC8; #100;
A = 8'hDC; B = 8'hC9; #100;
A = 8'hDC; B = 8'hCA; #100;
A = 8'hDC; B = 8'hCB; #100;
A = 8'hDC; B = 8'hCC; #100;
A = 8'hDC; B = 8'hCD; #100;
A = 8'hDC; B = 8'hCE; #100;
A = 8'hDC; B = 8'hCF; #100;
A = 8'hDC; B = 8'hD0; #100;
A = 8'hDC; B = 8'hD1; #100;
A = 8'hDC; B = 8'hD2; #100;
A = 8'hDC; B = 8'hD3; #100;
A = 8'hDC; B = 8'hD4; #100;
A = 8'hDC; B = 8'hD5; #100;
A = 8'hDC; B = 8'hD6; #100;
A = 8'hDC; B = 8'hD7; #100;
A = 8'hDC; B = 8'hD8; #100;
A = 8'hDC; B = 8'hD9; #100;
A = 8'hDC; B = 8'hDA; #100;
A = 8'hDC; B = 8'hDB; #100;
A = 8'hDC; B = 8'hDC; #100;
A = 8'hDC; B = 8'hDD; #100;
A = 8'hDC; B = 8'hDE; #100;
A = 8'hDC; B = 8'hDF; #100;
A = 8'hDC; B = 8'hE0; #100;
A = 8'hDC; B = 8'hE1; #100;
A = 8'hDC; B = 8'hE2; #100;
A = 8'hDC; B = 8'hE3; #100;
A = 8'hDC; B = 8'hE4; #100;
A = 8'hDC; B = 8'hE5; #100;
A = 8'hDC; B = 8'hE6; #100;
A = 8'hDC; B = 8'hE7; #100;
A = 8'hDC; B = 8'hE8; #100;
A = 8'hDC; B = 8'hE9; #100;
A = 8'hDC; B = 8'hEA; #100;
A = 8'hDC; B = 8'hEB; #100;
A = 8'hDC; B = 8'hEC; #100;
A = 8'hDC; B = 8'hED; #100;
A = 8'hDC; B = 8'hEE; #100;
A = 8'hDC; B = 8'hEF; #100;
A = 8'hDC; B = 8'hF0; #100;
A = 8'hDC; B = 8'hF1; #100;
A = 8'hDC; B = 8'hF2; #100;
A = 8'hDC; B = 8'hF3; #100;
A = 8'hDC; B = 8'hF4; #100;
A = 8'hDC; B = 8'hF5; #100;
A = 8'hDC; B = 8'hF6; #100;
A = 8'hDC; B = 8'hF7; #100;
A = 8'hDC; B = 8'hF8; #100;
A = 8'hDC; B = 8'hF9; #100;
A = 8'hDC; B = 8'hFA; #100;
A = 8'hDC; B = 8'hFB; #100;
A = 8'hDC; B = 8'hFC; #100;
A = 8'hDC; B = 8'hFD; #100;
A = 8'hDC; B = 8'hFE; #100;
A = 8'hDC; B = 8'hFF; #100;
A = 8'hDD; B = 8'h0; #100;
A = 8'hDD; B = 8'h1; #100;
A = 8'hDD; B = 8'h2; #100;
A = 8'hDD; B = 8'h3; #100;
A = 8'hDD; B = 8'h4; #100;
A = 8'hDD; B = 8'h5; #100;
A = 8'hDD; B = 8'h6; #100;
A = 8'hDD; B = 8'h7; #100;
A = 8'hDD; B = 8'h8; #100;
A = 8'hDD; B = 8'h9; #100;
A = 8'hDD; B = 8'hA; #100;
A = 8'hDD; B = 8'hB; #100;
A = 8'hDD; B = 8'hC; #100;
A = 8'hDD; B = 8'hD; #100;
A = 8'hDD; B = 8'hE; #100;
A = 8'hDD; B = 8'hF; #100;
A = 8'hDD; B = 8'h10; #100;
A = 8'hDD; B = 8'h11; #100;
A = 8'hDD; B = 8'h12; #100;
A = 8'hDD; B = 8'h13; #100;
A = 8'hDD; B = 8'h14; #100;
A = 8'hDD; B = 8'h15; #100;
A = 8'hDD; B = 8'h16; #100;
A = 8'hDD; B = 8'h17; #100;
A = 8'hDD; B = 8'h18; #100;
A = 8'hDD; B = 8'h19; #100;
A = 8'hDD; B = 8'h1A; #100;
A = 8'hDD; B = 8'h1B; #100;
A = 8'hDD; B = 8'h1C; #100;
A = 8'hDD; B = 8'h1D; #100;
A = 8'hDD; B = 8'h1E; #100;
A = 8'hDD; B = 8'h1F; #100;
A = 8'hDD; B = 8'h20; #100;
A = 8'hDD; B = 8'h21; #100;
A = 8'hDD; B = 8'h22; #100;
A = 8'hDD; B = 8'h23; #100;
A = 8'hDD; B = 8'h24; #100;
A = 8'hDD; B = 8'h25; #100;
A = 8'hDD; B = 8'h26; #100;
A = 8'hDD; B = 8'h27; #100;
A = 8'hDD; B = 8'h28; #100;
A = 8'hDD; B = 8'h29; #100;
A = 8'hDD; B = 8'h2A; #100;
A = 8'hDD; B = 8'h2B; #100;
A = 8'hDD; B = 8'h2C; #100;
A = 8'hDD; B = 8'h2D; #100;
A = 8'hDD; B = 8'h2E; #100;
A = 8'hDD; B = 8'h2F; #100;
A = 8'hDD; B = 8'h30; #100;
A = 8'hDD; B = 8'h31; #100;
A = 8'hDD; B = 8'h32; #100;
A = 8'hDD; B = 8'h33; #100;
A = 8'hDD; B = 8'h34; #100;
A = 8'hDD; B = 8'h35; #100;
A = 8'hDD; B = 8'h36; #100;
A = 8'hDD; B = 8'h37; #100;
A = 8'hDD; B = 8'h38; #100;
A = 8'hDD; B = 8'h39; #100;
A = 8'hDD; B = 8'h3A; #100;
A = 8'hDD; B = 8'h3B; #100;
A = 8'hDD; B = 8'h3C; #100;
A = 8'hDD; B = 8'h3D; #100;
A = 8'hDD; B = 8'h3E; #100;
A = 8'hDD; B = 8'h3F; #100;
A = 8'hDD; B = 8'h40; #100;
A = 8'hDD; B = 8'h41; #100;
A = 8'hDD; B = 8'h42; #100;
A = 8'hDD; B = 8'h43; #100;
A = 8'hDD; B = 8'h44; #100;
A = 8'hDD; B = 8'h45; #100;
A = 8'hDD; B = 8'h46; #100;
A = 8'hDD; B = 8'h47; #100;
A = 8'hDD; B = 8'h48; #100;
A = 8'hDD; B = 8'h49; #100;
A = 8'hDD; B = 8'h4A; #100;
A = 8'hDD; B = 8'h4B; #100;
A = 8'hDD; B = 8'h4C; #100;
A = 8'hDD; B = 8'h4D; #100;
A = 8'hDD; B = 8'h4E; #100;
A = 8'hDD; B = 8'h4F; #100;
A = 8'hDD; B = 8'h50; #100;
A = 8'hDD; B = 8'h51; #100;
A = 8'hDD; B = 8'h52; #100;
A = 8'hDD; B = 8'h53; #100;
A = 8'hDD; B = 8'h54; #100;
A = 8'hDD; B = 8'h55; #100;
A = 8'hDD; B = 8'h56; #100;
A = 8'hDD; B = 8'h57; #100;
A = 8'hDD; B = 8'h58; #100;
A = 8'hDD; B = 8'h59; #100;
A = 8'hDD; B = 8'h5A; #100;
A = 8'hDD; B = 8'h5B; #100;
A = 8'hDD; B = 8'h5C; #100;
A = 8'hDD; B = 8'h5D; #100;
A = 8'hDD; B = 8'h5E; #100;
A = 8'hDD; B = 8'h5F; #100;
A = 8'hDD; B = 8'h60; #100;
A = 8'hDD; B = 8'h61; #100;
A = 8'hDD; B = 8'h62; #100;
A = 8'hDD; B = 8'h63; #100;
A = 8'hDD; B = 8'h64; #100;
A = 8'hDD; B = 8'h65; #100;
A = 8'hDD; B = 8'h66; #100;
A = 8'hDD; B = 8'h67; #100;
A = 8'hDD; B = 8'h68; #100;
A = 8'hDD; B = 8'h69; #100;
A = 8'hDD; B = 8'h6A; #100;
A = 8'hDD; B = 8'h6B; #100;
A = 8'hDD; B = 8'h6C; #100;
A = 8'hDD; B = 8'h6D; #100;
A = 8'hDD; B = 8'h6E; #100;
A = 8'hDD; B = 8'h6F; #100;
A = 8'hDD; B = 8'h70; #100;
A = 8'hDD; B = 8'h71; #100;
A = 8'hDD; B = 8'h72; #100;
A = 8'hDD; B = 8'h73; #100;
A = 8'hDD; B = 8'h74; #100;
A = 8'hDD; B = 8'h75; #100;
A = 8'hDD; B = 8'h76; #100;
A = 8'hDD; B = 8'h77; #100;
A = 8'hDD; B = 8'h78; #100;
A = 8'hDD; B = 8'h79; #100;
A = 8'hDD; B = 8'h7A; #100;
A = 8'hDD; B = 8'h7B; #100;
A = 8'hDD; B = 8'h7C; #100;
A = 8'hDD; B = 8'h7D; #100;
A = 8'hDD; B = 8'h7E; #100;
A = 8'hDD; B = 8'h7F; #100;
A = 8'hDD; B = 8'h80; #100;
A = 8'hDD; B = 8'h81; #100;
A = 8'hDD; B = 8'h82; #100;
A = 8'hDD; B = 8'h83; #100;
A = 8'hDD; B = 8'h84; #100;
A = 8'hDD; B = 8'h85; #100;
A = 8'hDD; B = 8'h86; #100;
A = 8'hDD; B = 8'h87; #100;
A = 8'hDD; B = 8'h88; #100;
A = 8'hDD; B = 8'h89; #100;
A = 8'hDD; B = 8'h8A; #100;
A = 8'hDD; B = 8'h8B; #100;
A = 8'hDD; B = 8'h8C; #100;
A = 8'hDD; B = 8'h8D; #100;
A = 8'hDD; B = 8'h8E; #100;
A = 8'hDD; B = 8'h8F; #100;
A = 8'hDD; B = 8'h90; #100;
A = 8'hDD; B = 8'h91; #100;
A = 8'hDD; B = 8'h92; #100;
A = 8'hDD; B = 8'h93; #100;
A = 8'hDD; B = 8'h94; #100;
A = 8'hDD; B = 8'h95; #100;
A = 8'hDD; B = 8'h96; #100;
A = 8'hDD; B = 8'h97; #100;
A = 8'hDD; B = 8'h98; #100;
A = 8'hDD; B = 8'h99; #100;
A = 8'hDD; B = 8'h9A; #100;
A = 8'hDD; B = 8'h9B; #100;
A = 8'hDD; B = 8'h9C; #100;
A = 8'hDD; B = 8'h9D; #100;
A = 8'hDD; B = 8'h9E; #100;
A = 8'hDD; B = 8'h9F; #100;
A = 8'hDD; B = 8'hA0; #100;
A = 8'hDD; B = 8'hA1; #100;
A = 8'hDD; B = 8'hA2; #100;
A = 8'hDD; B = 8'hA3; #100;
A = 8'hDD; B = 8'hA4; #100;
A = 8'hDD; B = 8'hA5; #100;
A = 8'hDD; B = 8'hA6; #100;
A = 8'hDD; B = 8'hA7; #100;
A = 8'hDD; B = 8'hA8; #100;
A = 8'hDD; B = 8'hA9; #100;
A = 8'hDD; B = 8'hAA; #100;
A = 8'hDD; B = 8'hAB; #100;
A = 8'hDD; B = 8'hAC; #100;
A = 8'hDD; B = 8'hAD; #100;
A = 8'hDD; B = 8'hAE; #100;
A = 8'hDD; B = 8'hAF; #100;
A = 8'hDD; B = 8'hB0; #100;
A = 8'hDD; B = 8'hB1; #100;
A = 8'hDD; B = 8'hB2; #100;
A = 8'hDD; B = 8'hB3; #100;
A = 8'hDD; B = 8'hB4; #100;
A = 8'hDD; B = 8'hB5; #100;
A = 8'hDD; B = 8'hB6; #100;
A = 8'hDD; B = 8'hB7; #100;
A = 8'hDD; B = 8'hB8; #100;
A = 8'hDD; B = 8'hB9; #100;
A = 8'hDD; B = 8'hBA; #100;
A = 8'hDD; B = 8'hBB; #100;
A = 8'hDD; B = 8'hBC; #100;
A = 8'hDD; B = 8'hBD; #100;
A = 8'hDD; B = 8'hBE; #100;
A = 8'hDD; B = 8'hBF; #100;
A = 8'hDD; B = 8'hC0; #100;
A = 8'hDD; B = 8'hC1; #100;
A = 8'hDD; B = 8'hC2; #100;
A = 8'hDD; B = 8'hC3; #100;
A = 8'hDD; B = 8'hC4; #100;
A = 8'hDD; B = 8'hC5; #100;
A = 8'hDD; B = 8'hC6; #100;
A = 8'hDD; B = 8'hC7; #100;
A = 8'hDD; B = 8'hC8; #100;
A = 8'hDD; B = 8'hC9; #100;
A = 8'hDD; B = 8'hCA; #100;
A = 8'hDD; B = 8'hCB; #100;
A = 8'hDD; B = 8'hCC; #100;
A = 8'hDD; B = 8'hCD; #100;
A = 8'hDD; B = 8'hCE; #100;
A = 8'hDD; B = 8'hCF; #100;
A = 8'hDD; B = 8'hD0; #100;
A = 8'hDD; B = 8'hD1; #100;
A = 8'hDD; B = 8'hD2; #100;
A = 8'hDD; B = 8'hD3; #100;
A = 8'hDD; B = 8'hD4; #100;
A = 8'hDD; B = 8'hD5; #100;
A = 8'hDD; B = 8'hD6; #100;
A = 8'hDD; B = 8'hD7; #100;
A = 8'hDD; B = 8'hD8; #100;
A = 8'hDD; B = 8'hD9; #100;
A = 8'hDD; B = 8'hDA; #100;
A = 8'hDD; B = 8'hDB; #100;
A = 8'hDD; B = 8'hDC; #100;
A = 8'hDD; B = 8'hDD; #100;
A = 8'hDD; B = 8'hDE; #100;
A = 8'hDD; B = 8'hDF; #100;
A = 8'hDD; B = 8'hE0; #100;
A = 8'hDD; B = 8'hE1; #100;
A = 8'hDD; B = 8'hE2; #100;
A = 8'hDD; B = 8'hE3; #100;
A = 8'hDD; B = 8'hE4; #100;
A = 8'hDD; B = 8'hE5; #100;
A = 8'hDD; B = 8'hE6; #100;
A = 8'hDD; B = 8'hE7; #100;
A = 8'hDD; B = 8'hE8; #100;
A = 8'hDD; B = 8'hE9; #100;
A = 8'hDD; B = 8'hEA; #100;
A = 8'hDD; B = 8'hEB; #100;
A = 8'hDD; B = 8'hEC; #100;
A = 8'hDD; B = 8'hED; #100;
A = 8'hDD; B = 8'hEE; #100;
A = 8'hDD; B = 8'hEF; #100;
A = 8'hDD; B = 8'hF0; #100;
A = 8'hDD; B = 8'hF1; #100;
A = 8'hDD; B = 8'hF2; #100;
A = 8'hDD; B = 8'hF3; #100;
A = 8'hDD; B = 8'hF4; #100;
A = 8'hDD; B = 8'hF5; #100;
A = 8'hDD; B = 8'hF6; #100;
A = 8'hDD; B = 8'hF7; #100;
A = 8'hDD; B = 8'hF8; #100;
A = 8'hDD; B = 8'hF9; #100;
A = 8'hDD; B = 8'hFA; #100;
A = 8'hDD; B = 8'hFB; #100;
A = 8'hDD; B = 8'hFC; #100;
A = 8'hDD; B = 8'hFD; #100;
A = 8'hDD; B = 8'hFE; #100;
A = 8'hDD; B = 8'hFF; #100;
A = 8'hDE; B = 8'h0; #100;
A = 8'hDE; B = 8'h1; #100;
A = 8'hDE; B = 8'h2; #100;
A = 8'hDE; B = 8'h3; #100;
A = 8'hDE; B = 8'h4; #100;
A = 8'hDE; B = 8'h5; #100;
A = 8'hDE; B = 8'h6; #100;
A = 8'hDE; B = 8'h7; #100;
A = 8'hDE; B = 8'h8; #100;
A = 8'hDE; B = 8'h9; #100;
A = 8'hDE; B = 8'hA; #100;
A = 8'hDE; B = 8'hB; #100;
A = 8'hDE; B = 8'hC; #100;
A = 8'hDE; B = 8'hD; #100;
A = 8'hDE; B = 8'hE; #100;
A = 8'hDE; B = 8'hF; #100;
A = 8'hDE; B = 8'h10; #100;
A = 8'hDE; B = 8'h11; #100;
A = 8'hDE; B = 8'h12; #100;
A = 8'hDE; B = 8'h13; #100;
A = 8'hDE; B = 8'h14; #100;
A = 8'hDE; B = 8'h15; #100;
A = 8'hDE; B = 8'h16; #100;
A = 8'hDE; B = 8'h17; #100;
A = 8'hDE; B = 8'h18; #100;
A = 8'hDE; B = 8'h19; #100;
A = 8'hDE; B = 8'h1A; #100;
A = 8'hDE; B = 8'h1B; #100;
A = 8'hDE; B = 8'h1C; #100;
A = 8'hDE; B = 8'h1D; #100;
A = 8'hDE; B = 8'h1E; #100;
A = 8'hDE; B = 8'h1F; #100;
A = 8'hDE; B = 8'h20; #100;
A = 8'hDE; B = 8'h21; #100;
A = 8'hDE; B = 8'h22; #100;
A = 8'hDE; B = 8'h23; #100;
A = 8'hDE; B = 8'h24; #100;
A = 8'hDE; B = 8'h25; #100;
A = 8'hDE; B = 8'h26; #100;
A = 8'hDE; B = 8'h27; #100;
A = 8'hDE; B = 8'h28; #100;
A = 8'hDE; B = 8'h29; #100;
A = 8'hDE; B = 8'h2A; #100;
A = 8'hDE; B = 8'h2B; #100;
A = 8'hDE; B = 8'h2C; #100;
A = 8'hDE; B = 8'h2D; #100;
A = 8'hDE; B = 8'h2E; #100;
A = 8'hDE; B = 8'h2F; #100;
A = 8'hDE; B = 8'h30; #100;
A = 8'hDE; B = 8'h31; #100;
A = 8'hDE; B = 8'h32; #100;
A = 8'hDE; B = 8'h33; #100;
A = 8'hDE; B = 8'h34; #100;
A = 8'hDE; B = 8'h35; #100;
A = 8'hDE; B = 8'h36; #100;
A = 8'hDE; B = 8'h37; #100;
A = 8'hDE; B = 8'h38; #100;
A = 8'hDE; B = 8'h39; #100;
A = 8'hDE; B = 8'h3A; #100;
A = 8'hDE; B = 8'h3B; #100;
A = 8'hDE; B = 8'h3C; #100;
A = 8'hDE; B = 8'h3D; #100;
A = 8'hDE; B = 8'h3E; #100;
A = 8'hDE; B = 8'h3F; #100;
A = 8'hDE; B = 8'h40; #100;
A = 8'hDE; B = 8'h41; #100;
A = 8'hDE; B = 8'h42; #100;
A = 8'hDE; B = 8'h43; #100;
A = 8'hDE; B = 8'h44; #100;
A = 8'hDE; B = 8'h45; #100;
A = 8'hDE; B = 8'h46; #100;
A = 8'hDE; B = 8'h47; #100;
A = 8'hDE; B = 8'h48; #100;
A = 8'hDE; B = 8'h49; #100;
A = 8'hDE; B = 8'h4A; #100;
A = 8'hDE; B = 8'h4B; #100;
A = 8'hDE; B = 8'h4C; #100;
A = 8'hDE; B = 8'h4D; #100;
A = 8'hDE; B = 8'h4E; #100;
A = 8'hDE; B = 8'h4F; #100;
A = 8'hDE; B = 8'h50; #100;
A = 8'hDE; B = 8'h51; #100;
A = 8'hDE; B = 8'h52; #100;
A = 8'hDE; B = 8'h53; #100;
A = 8'hDE; B = 8'h54; #100;
A = 8'hDE; B = 8'h55; #100;
A = 8'hDE; B = 8'h56; #100;
A = 8'hDE; B = 8'h57; #100;
A = 8'hDE; B = 8'h58; #100;
A = 8'hDE; B = 8'h59; #100;
A = 8'hDE; B = 8'h5A; #100;
A = 8'hDE; B = 8'h5B; #100;
A = 8'hDE; B = 8'h5C; #100;
A = 8'hDE; B = 8'h5D; #100;
A = 8'hDE; B = 8'h5E; #100;
A = 8'hDE; B = 8'h5F; #100;
A = 8'hDE; B = 8'h60; #100;
A = 8'hDE; B = 8'h61; #100;
A = 8'hDE; B = 8'h62; #100;
A = 8'hDE; B = 8'h63; #100;
A = 8'hDE; B = 8'h64; #100;
A = 8'hDE; B = 8'h65; #100;
A = 8'hDE; B = 8'h66; #100;
A = 8'hDE; B = 8'h67; #100;
A = 8'hDE; B = 8'h68; #100;
A = 8'hDE; B = 8'h69; #100;
A = 8'hDE; B = 8'h6A; #100;
A = 8'hDE; B = 8'h6B; #100;
A = 8'hDE; B = 8'h6C; #100;
A = 8'hDE; B = 8'h6D; #100;
A = 8'hDE; B = 8'h6E; #100;
A = 8'hDE; B = 8'h6F; #100;
A = 8'hDE; B = 8'h70; #100;
A = 8'hDE; B = 8'h71; #100;
A = 8'hDE; B = 8'h72; #100;
A = 8'hDE; B = 8'h73; #100;
A = 8'hDE; B = 8'h74; #100;
A = 8'hDE; B = 8'h75; #100;
A = 8'hDE; B = 8'h76; #100;
A = 8'hDE; B = 8'h77; #100;
A = 8'hDE; B = 8'h78; #100;
A = 8'hDE; B = 8'h79; #100;
A = 8'hDE; B = 8'h7A; #100;
A = 8'hDE; B = 8'h7B; #100;
A = 8'hDE; B = 8'h7C; #100;
A = 8'hDE; B = 8'h7D; #100;
A = 8'hDE; B = 8'h7E; #100;
A = 8'hDE; B = 8'h7F; #100;
A = 8'hDE; B = 8'h80; #100;
A = 8'hDE; B = 8'h81; #100;
A = 8'hDE; B = 8'h82; #100;
A = 8'hDE; B = 8'h83; #100;
A = 8'hDE; B = 8'h84; #100;
A = 8'hDE; B = 8'h85; #100;
A = 8'hDE; B = 8'h86; #100;
A = 8'hDE; B = 8'h87; #100;
A = 8'hDE; B = 8'h88; #100;
A = 8'hDE; B = 8'h89; #100;
A = 8'hDE; B = 8'h8A; #100;
A = 8'hDE; B = 8'h8B; #100;
A = 8'hDE; B = 8'h8C; #100;
A = 8'hDE; B = 8'h8D; #100;
A = 8'hDE; B = 8'h8E; #100;
A = 8'hDE; B = 8'h8F; #100;
A = 8'hDE; B = 8'h90; #100;
A = 8'hDE; B = 8'h91; #100;
A = 8'hDE; B = 8'h92; #100;
A = 8'hDE; B = 8'h93; #100;
A = 8'hDE; B = 8'h94; #100;
A = 8'hDE; B = 8'h95; #100;
A = 8'hDE; B = 8'h96; #100;
A = 8'hDE; B = 8'h97; #100;
A = 8'hDE; B = 8'h98; #100;
A = 8'hDE; B = 8'h99; #100;
A = 8'hDE; B = 8'h9A; #100;
A = 8'hDE; B = 8'h9B; #100;
A = 8'hDE; B = 8'h9C; #100;
A = 8'hDE; B = 8'h9D; #100;
A = 8'hDE; B = 8'h9E; #100;
A = 8'hDE; B = 8'h9F; #100;
A = 8'hDE; B = 8'hA0; #100;
A = 8'hDE; B = 8'hA1; #100;
A = 8'hDE; B = 8'hA2; #100;
A = 8'hDE; B = 8'hA3; #100;
A = 8'hDE; B = 8'hA4; #100;
A = 8'hDE; B = 8'hA5; #100;
A = 8'hDE; B = 8'hA6; #100;
A = 8'hDE; B = 8'hA7; #100;
A = 8'hDE; B = 8'hA8; #100;
A = 8'hDE; B = 8'hA9; #100;
A = 8'hDE; B = 8'hAA; #100;
A = 8'hDE; B = 8'hAB; #100;
A = 8'hDE; B = 8'hAC; #100;
A = 8'hDE; B = 8'hAD; #100;
A = 8'hDE; B = 8'hAE; #100;
A = 8'hDE; B = 8'hAF; #100;
A = 8'hDE; B = 8'hB0; #100;
A = 8'hDE; B = 8'hB1; #100;
A = 8'hDE; B = 8'hB2; #100;
A = 8'hDE; B = 8'hB3; #100;
A = 8'hDE; B = 8'hB4; #100;
A = 8'hDE; B = 8'hB5; #100;
A = 8'hDE; B = 8'hB6; #100;
A = 8'hDE; B = 8'hB7; #100;
A = 8'hDE; B = 8'hB8; #100;
A = 8'hDE; B = 8'hB9; #100;
A = 8'hDE; B = 8'hBA; #100;
A = 8'hDE; B = 8'hBB; #100;
A = 8'hDE; B = 8'hBC; #100;
A = 8'hDE; B = 8'hBD; #100;
A = 8'hDE; B = 8'hBE; #100;
A = 8'hDE; B = 8'hBF; #100;
A = 8'hDE; B = 8'hC0; #100;
A = 8'hDE; B = 8'hC1; #100;
A = 8'hDE; B = 8'hC2; #100;
A = 8'hDE; B = 8'hC3; #100;
A = 8'hDE; B = 8'hC4; #100;
A = 8'hDE; B = 8'hC5; #100;
A = 8'hDE; B = 8'hC6; #100;
A = 8'hDE; B = 8'hC7; #100;
A = 8'hDE; B = 8'hC8; #100;
A = 8'hDE; B = 8'hC9; #100;
A = 8'hDE; B = 8'hCA; #100;
A = 8'hDE; B = 8'hCB; #100;
A = 8'hDE; B = 8'hCC; #100;
A = 8'hDE; B = 8'hCD; #100;
A = 8'hDE; B = 8'hCE; #100;
A = 8'hDE; B = 8'hCF; #100;
A = 8'hDE; B = 8'hD0; #100;
A = 8'hDE; B = 8'hD1; #100;
A = 8'hDE; B = 8'hD2; #100;
A = 8'hDE; B = 8'hD3; #100;
A = 8'hDE; B = 8'hD4; #100;
A = 8'hDE; B = 8'hD5; #100;
A = 8'hDE; B = 8'hD6; #100;
A = 8'hDE; B = 8'hD7; #100;
A = 8'hDE; B = 8'hD8; #100;
A = 8'hDE; B = 8'hD9; #100;
A = 8'hDE; B = 8'hDA; #100;
A = 8'hDE; B = 8'hDB; #100;
A = 8'hDE; B = 8'hDC; #100;
A = 8'hDE; B = 8'hDD; #100;
A = 8'hDE; B = 8'hDE; #100;
A = 8'hDE; B = 8'hDF; #100;
A = 8'hDE; B = 8'hE0; #100;
A = 8'hDE; B = 8'hE1; #100;
A = 8'hDE; B = 8'hE2; #100;
A = 8'hDE; B = 8'hE3; #100;
A = 8'hDE; B = 8'hE4; #100;
A = 8'hDE; B = 8'hE5; #100;
A = 8'hDE; B = 8'hE6; #100;
A = 8'hDE; B = 8'hE7; #100;
A = 8'hDE; B = 8'hE8; #100;
A = 8'hDE; B = 8'hE9; #100;
A = 8'hDE; B = 8'hEA; #100;
A = 8'hDE; B = 8'hEB; #100;
A = 8'hDE; B = 8'hEC; #100;
A = 8'hDE; B = 8'hED; #100;
A = 8'hDE; B = 8'hEE; #100;
A = 8'hDE; B = 8'hEF; #100;
A = 8'hDE; B = 8'hF0; #100;
A = 8'hDE; B = 8'hF1; #100;
A = 8'hDE; B = 8'hF2; #100;
A = 8'hDE; B = 8'hF3; #100;
A = 8'hDE; B = 8'hF4; #100;
A = 8'hDE; B = 8'hF5; #100;
A = 8'hDE; B = 8'hF6; #100;
A = 8'hDE; B = 8'hF7; #100;
A = 8'hDE; B = 8'hF8; #100;
A = 8'hDE; B = 8'hF9; #100;
A = 8'hDE; B = 8'hFA; #100;
A = 8'hDE; B = 8'hFB; #100;
A = 8'hDE; B = 8'hFC; #100;
A = 8'hDE; B = 8'hFD; #100;
A = 8'hDE; B = 8'hFE; #100;
A = 8'hDE; B = 8'hFF; #100;
A = 8'hDF; B = 8'h0; #100;
A = 8'hDF; B = 8'h1; #100;
A = 8'hDF; B = 8'h2; #100;
A = 8'hDF; B = 8'h3; #100;
A = 8'hDF; B = 8'h4; #100;
A = 8'hDF; B = 8'h5; #100;
A = 8'hDF; B = 8'h6; #100;
A = 8'hDF; B = 8'h7; #100;
A = 8'hDF; B = 8'h8; #100;
A = 8'hDF; B = 8'h9; #100;
A = 8'hDF; B = 8'hA; #100;
A = 8'hDF; B = 8'hB; #100;
A = 8'hDF; B = 8'hC; #100;
A = 8'hDF; B = 8'hD; #100;
A = 8'hDF; B = 8'hE; #100;
A = 8'hDF; B = 8'hF; #100;
A = 8'hDF; B = 8'h10; #100;
A = 8'hDF; B = 8'h11; #100;
A = 8'hDF; B = 8'h12; #100;
A = 8'hDF; B = 8'h13; #100;
A = 8'hDF; B = 8'h14; #100;
A = 8'hDF; B = 8'h15; #100;
A = 8'hDF; B = 8'h16; #100;
A = 8'hDF; B = 8'h17; #100;
A = 8'hDF; B = 8'h18; #100;
A = 8'hDF; B = 8'h19; #100;
A = 8'hDF; B = 8'h1A; #100;
A = 8'hDF; B = 8'h1B; #100;
A = 8'hDF; B = 8'h1C; #100;
A = 8'hDF; B = 8'h1D; #100;
A = 8'hDF; B = 8'h1E; #100;
A = 8'hDF; B = 8'h1F; #100;
A = 8'hDF; B = 8'h20; #100;
A = 8'hDF; B = 8'h21; #100;
A = 8'hDF; B = 8'h22; #100;
A = 8'hDF; B = 8'h23; #100;
A = 8'hDF; B = 8'h24; #100;
A = 8'hDF; B = 8'h25; #100;
A = 8'hDF; B = 8'h26; #100;
A = 8'hDF; B = 8'h27; #100;
A = 8'hDF; B = 8'h28; #100;
A = 8'hDF; B = 8'h29; #100;
A = 8'hDF; B = 8'h2A; #100;
A = 8'hDF; B = 8'h2B; #100;
A = 8'hDF; B = 8'h2C; #100;
A = 8'hDF; B = 8'h2D; #100;
A = 8'hDF; B = 8'h2E; #100;
A = 8'hDF; B = 8'h2F; #100;
A = 8'hDF; B = 8'h30; #100;
A = 8'hDF; B = 8'h31; #100;
A = 8'hDF; B = 8'h32; #100;
A = 8'hDF; B = 8'h33; #100;
A = 8'hDF; B = 8'h34; #100;
A = 8'hDF; B = 8'h35; #100;
A = 8'hDF; B = 8'h36; #100;
A = 8'hDF; B = 8'h37; #100;
A = 8'hDF; B = 8'h38; #100;
A = 8'hDF; B = 8'h39; #100;
A = 8'hDF; B = 8'h3A; #100;
A = 8'hDF; B = 8'h3B; #100;
A = 8'hDF; B = 8'h3C; #100;
A = 8'hDF; B = 8'h3D; #100;
A = 8'hDF; B = 8'h3E; #100;
A = 8'hDF; B = 8'h3F; #100;
A = 8'hDF; B = 8'h40; #100;
A = 8'hDF; B = 8'h41; #100;
A = 8'hDF; B = 8'h42; #100;
A = 8'hDF; B = 8'h43; #100;
A = 8'hDF; B = 8'h44; #100;
A = 8'hDF; B = 8'h45; #100;
A = 8'hDF; B = 8'h46; #100;
A = 8'hDF; B = 8'h47; #100;
A = 8'hDF; B = 8'h48; #100;
A = 8'hDF; B = 8'h49; #100;
A = 8'hDF; B = 8'h4A; #100;
A = 8'hDF; B = 8'h4B; #100;
A = 8'hDF; B = 8'h4C; #100;
A = 8'hDF; B = 8'h4D; #100;
A = 8'hDF; B = 8'h4E; #100;
A = 8'hDF; B = 8'h4F; #100;
A = 8'hDF; B = 8'h50; #100;
A = 8'hDF; B = 8'h51; #100;
A = 8'hDF; B = 8'h52; #100;
A = 8'hDF; B = 8'h53; #100;
A = 8'hDF; B = 8'h54; #100;
A = 8'hDF; B = 8'h55; #100;
A = 8'hDF; B = 8'h56; #100;
A = 8'hDF; B = 8'h57; #100;
A = 8'hDF; B = 8'h58; #100;
A = 8'hDF; B = 8'h59; #100;
A = 8'hDF; B = 8'h5A; #100;
A = 8'hDF; B = 8'h5B; #100;
A = 8'hDF; B = 8'h5C; #100;
A = 8'hDF; B = 8'h5D; #100;
A = 8'hDF; B = 8'h5E; #100;
A = 8'hDF; B = 8'h5F; #100;
A = 8'hDF; B = 8'h60; #100;
A = 8'hDF; B = 8'h61; #100;
A = 8'hDF; B = 8'h62; #100;
A = 8'hDF; B = 8'h63; #100;
A = 8'hDF; B = 8'h64; #100;
A = 8'hDF; B = 8'h65; #100;
A = 8'hDF; B = 8'h66; #100;
A = 8'hDF; B = 8'h67; #100;
A = 8'hDF; B = 8'h68; #100;
A = 8'hDF; B = 8'h69; #100;
A = 8'hDF; B = 8'h6A; #100;
A = 8'hDF; B = 8'h6B; #100;
A = 8'hDF; B = 8'h6C; #100;
A = 8'hDF; B = 8'h6D; #100;
A = 8'hDF; B = 8'h6E; #100;
A = 8'hDF; B = 8'h6F; #100;
A = 8'hDF; B = 8'h70; #100;
A = 8'hDF; B = 8'h71; #100;
A = 8'hDF; B = 8'h72; #100;
A = 8'hDF; B = 8'h73; #100;
A = 8'hDF; B = 8'h74; #100;
A = 8'hDF; B = 8'h75; #100;
A = 8'hDF; B = 8'h76; #100;
A = 8'hDF; B = 8'h77; #100;
A = 8'hDF; B = 8'h78; #100;
A = 8'hDF; B = 8'h79; #100;
A = 8'hDF; B = 8'h7A; #100;
A = 8'hDF; B = 8'h7B; #100;
A = 8'hDF; B = 8'h7C; #100;
A = 8'hDF; B = 8'h7D; #100;
A = 8'hDF; B = 8'h7E; #100;
A = 8'hDF; B = 8'h7F; #100;
A = 8'hDF; B = 8'h80; #100;
A = 8'hDF; B = 8'h81; #100;
A = 8'hDF; B = 8'h82; #100;
A = 8'hDF; B = 8'h83; #100;
A = 8'hDF; B = 8'h84; #100;
A = 8'hDF; B = 8'h85; #100;
A = 8'hDF; B = 8'h86; #100;
A = 8'hDF; B = 8'h87; #100;
A = 8'hDF; B = 8'h88; #100;
A = 8'hDF; B = 8'h89; #100;
A = 8'hDF; B = 8'h8A; #100;
A = 8'hDF; B = 8'h8B; #100;
A = 8'hDF; B = 8'h8C; #100;
A = 8'hDF; B = 8'h8D; #100;
A = 8'hDF; B = 8'h8E; #100;
A = 8'hDF; B = 8'h8F; #100;
A = 8'hDF; B = 8'h90; #100;
A = 8'hDF; B = 8'h91; #100;
A = 8'hDF; B = 8'h92; #100;
A = 8'hDF; B = 8'h93; #100;
A = 8'hDF; B = 8'h94; #100;
A = 8'hDF; B = 8'h95; #100;
A = 8'hDF; B = 8'h96; #100;
A = 8'hDF; B = 8'h97; #100;
A = 8'hDF; B = 8'h98; #100;
A = 8'hDF; B = 8'h99; #100;
A = 8'hDF; B = 8'h9A; #100;
A = 8'hDF; B = 8'h9B; #100;
A = 8'hDF; B = 8'h9C; #100;
A = 8'hDF; B = 8'h9D; #100;
A = 8'hDF; B = 8'h9E; #100;
A = 8'hDF; B = 8'h9F; #100;
A = 8'hDF; B = 8'hA0; #100;
A = 8'hDF; B = 8'hA1; #100;
A = 8'hDF; B = 8'hA2; #100;
A = 8'hDF; B = 8'hA3; #100;
A = 8'hDF; B = 8'hA4; #100;
A = 8'hDF; B = 8'hA5; #100;
A = 8'hDF; B = 8'hA6; #100;
A = 8'hDF; B = 8'hA7; #100;
A = 8'hDF; B = 8'hA8; #100;
A = 8'hDF; B = 8'hA9; #100;
A = 8'hDF; B = 8'hAA; #100;
A = 8'hDF; B = 8'hAB; #100;
A = 8'hDF; B = 8'hAC; #100;
A = 8'hDF; B = 8'hAD; #100;
A = 8'hDF; B = 8'hAE; #100;
A = 8'hDF; B = 8'hAF; #100;
A = 8'hDF; B = 8'hB0; #100;
A = 8'hDF; B = 8'hB1; #100;
A = 8'hDF; B = 8'hB2; #100;
A = 8'hDF; B = 8'hB3; #100;
A = 8'hDF; B = 8'hB4; #100;
A = 8'hDF; B = 8'hB5; #100;
A = 8'hDF; B = 8'hB6; #100;
A = 8'hDF; B = 8'hB7; #100;
A = 8'hDF; B = 8'hB8; #100;
A = 8'hDF; B = 8'hB9; #100;
A = 8'hDF; B = 8'hBA; #100;
A = 8'hDF; B = 8'hBB; #100;
A = 8'hDF; B = 8'hBC; #100;
A = 8'hDF; B = 8'hBD; #100;
A = 8'hDF; B = 8'hBE; #100;
A = 8'hDF; B = 8'hBF; #100;
A = 8'hDF; B = 8'hC0; #100;
A = 8'hDF; B = 8'hC1; #100;
A = 8'hDF; B = 8'hC2; #100;
A = 8'hDF; B = 8'hC3; #100;
A = 8'hDF; B = 8'hC4; #100;
A = 8'hDF; B = 8'hC5; #100;
A = 8'hDF; B = 8'hC6; #100;
A = 8'hDF; B = 8'hC7; #100;
A = 8'hDF; B = 8'hC8; #100;
A = 8'hDF; B = 8'hC9; #100;
A = 8'hDF; B = 8'hCA; #100;
A = 8'hDF; B = 8'hCB; #100;
A = 8'hDF; B = 8'hCC; #100;
A = 8'hDF; B = 8'hCD; #100;
A = 8'hDF; B = 8'hCE; #100;
A = 8'hDF; B = 8'hCF; #100;
A = 8'hDF; B = 8'hD0; #100;
A = 8'hDF; B = 8'hD1; #100;
A = 8'hDF; B = 8'hD2; #100;
A = 8'hDF; B = 8'hD3; #100;
A = 8'hDF; B = 8'hD4; #100;
A = 8'hDF; B = 8'hD5; #100;
A = 8'hDF; B = 8'hD6; #100;
A = 8'hDF; B = 8'hD7; #100;
A = 8'hDF; B = 8'hD8; #100;
A = 8'hDF; B = 8'hD9; #100;
A = 8'hDF; B = 8'hDA; #100;
A = 8'hDF; B = 8'hDB; #100;
A = 8'hDF; B = 8'hDC; #100;
A = 8'hDF; B = 8'hDD; #100;
A = 8'hDF; B = 8'hDE; #100;
A = 8'hDF; B = 8'hDF; #100;
A = 8'hDF; B = 8'hE0; #100;
A = 8'hDF; B = 8'hE1; #100;
A = 8'hDF; B = 8'hE2; #100;
A = 8'hDF; B = 8'hE3; #100;
A = 8'hDF; B = 8'hE4; #100;
A = 8'hDF; B = 8'hE5; #100;
A = 8'hDF; B = 8'hE6; #100;
A = 8'hDF; B = 8'hE7; #100;
A = 8'hDF; B = 8'hE8; #100;
A = 8'hDF; B = 8'hE9; #100;
A = 8'hDF; B = 8'hEA; #100;
A = 8'hDF; B = 8'hEB; #100;
A = 8'hDF; B = 8'hEC; #100;
A = 8'hDF; B = 8'hED; #100;
A = 8'hDF; B = 8'hEE; #100;
A = 8'hDF; B = 8'hEF; #100;
A = 8'hDF; B = 8'hF0; #100;
A = 8'hDF; B = 8'hF1; #100;
A = 8'hDF; B = 8'hF2; #100;
A = 8'hDF; B = 8'hF3; #100;
A = 8'hDF; B = 8'hF4; #100;
A = 8'hDF; B = 8'hF5; #100;
A = 8'hDF; B = 8'hF6; #100;
A = 8'hDF; B = 8'hF7; #100;
A = 8'hDF; B = 8'hF8; #100;
A = 8'hDF; B = 8'hF9; #100;
A = 8'hDF; B = 8'hFA; #100;
A = 8'hDF; B = 8'hFB; #100;
A = 8'hDF; B = 8'hFC; #100;
A = 8'hDF; B = 8'hFD; #100;
A = 8'hDF; B = 8'hFE; #100;
A = 8'hDF; B = 8'hFF; #100;
A = 8'hE0; B = 8'h0; #100;
A = 8'hE0; B = 8'h1; #100;
A = 8'hE0; B = 8'h2; #100;
A = 8'hE0; B = 8'h3; #100;
A = 8'hE0; B = 8'h4; #100;
A = 8'hE0; B = 8'h5; #100;
A = 8'hE0; B = 8'h6; #100;
A = 8'hE0; B = 8'h7; #100;
A = 8'hE0; B = 8'h8; #100;
A = 8'hE0; B = 8'h9; #100;
A = 8'hE0; B = 8'hA; #100;
A = 8'hE0; B = 8'hB; #100;
A = 8'hE0; B = 8'hC; #100;
A = 8'hE0; B = 8'hD; #100;
A = 8'hE0; B = 8'hE; #100;
A = 8'hE0; B = 8'hF; #100;
A = 8'hE0; B = 8'h10; #100;
A = 8'hE0; B = 8'h11; #100;
A = 8'hE0; B = 8'h12; #100;
A = 8'hE0; B = 8'h13; #100;
A = 8'hE0; B = 8'h14; #100;
A = 8'hE0; B = 8'h15; #100;
A = 8'hE0; B = 8'h16; #100;
A = 8'hE0; B = 8'h17; #100;
A = 8'hE0; B = 8'h18; #100;
A = 8'hE0; B = 8'h19; #100;
A = 8'hE0; B = 8'h1A; #100;
A = 8'hE0; B = 8'h1B; #100;
A = 8'hE0; B = 8'h1C; #100;
A = 8'hE0; B = 8'h1D; #100;
A = 8'hE0; B = 8'h1E; #100;
A = 8'hE0; B = 8'h1F; #100;
A = 8'hE0; B = 8'h20; #100;
A = 8'hE0; B = 8'h21; #100;
A = 8'hE0; B = 8'h22; #100;
A = 8'hE0; B = 8'h23; #100;
A = 8'hE0; B = 8'h24; #100;
A = 8'hE0; B = 8'h25; #100;
A = 8'hE0; B = 8'h26; #100;
A = 8'hE0; B = 8'h27; #100;
A = 8'hE0; B = 8'h28; #100;
A = 8'hE0; B = 8'h29; #100;
A = 8'hE0; B = 8'h2A; #100;
A = 8'hE0; B = 8'h2B; #100;
A = 8'hE0; B = 8'h2C; #100;
A = 8'hE0; B = 8'h2D; #100;
A = 8'hE0; B = 8'h2E; #100;
A = 8'hE0; B = 8'h2F; #100;
A = 8'hE0; B = 8'h30; #100;
A = 8'hE0; B = 8'h31; #100;
A = 8'hE0; B = 8'h32; #100;
A = 8'hE0; B = 8'h33; #100;
A = 8'hE0; B = 8'h34; #100;
A = 8'hE0; B = 8'h35; #100;
A = 8'hE0; B = 8'h36; #100;
A = 8'hE0; B = 8'h37; #100;
A = 8'hE0; B = 8'h38; #100;
A = 8'hE0; B = 8'h39; #100;
A = 8'hE0; B = 8'h3A; #100;
A = 8'hE0; B = 8'h3B; #100;
A = 8'hE0; B = 8'h3C; #100;
A = 8'hE0; B = 8'h3D; #100;
A = 8'hE0; B = 8'h3E; #100;
A = 8'hE0; B = 8'h3F; #100;
A = 8'hE0; B = 8'h40; #100;
A = 8'hE0; B = 8'h41; #100;
A = 8'hE0; B = 8'h42; #100;
A = 8'hE0; B = 8'h43; #100;
A = 8'hE0; B = 8'h44; #100;
A = 8'hE0; B = 8'h45; #100;
A = 8'hE0; B = 8'h46; #100;
A = 8'hE0; B = 8'h47; #100;
A = 8'hE0; B = 8'h48; #100;
A = 8'hE0; B = 8'h49; #100;
A = 8'hE0; B = 8'h4A; #100;
A = 8'hE0; B = 8'h4B; #100;
A = 8'hE0; B = 8'h4C; #100;
A = 8'hE0; B = 8'h4D; #100;
A = 8'hE0; B = 8'h4E; #100;
A = 8'hE0; B = 8'h4F; #100;
A = 8'hE0; B = 8'h50; #100;
A = 8'hE0; B = 8'h51; #100;
A = 8'hE0; B = 8'h52; #100;
A = 8'hE0; B = 8'h53; #100;
A = 8'hE0; B = 8'h54; #100;
A = 8'hE0; B = 8'h55; #100;
A = 8'hE0; B = 8'h56; #100;
A = 8'hE0; B = 8'h57; #100;
A = 8'hE0; B = 8'h58; #100;
A = 8'hE0; B = 8'h59; #100;
A = 8'hE0; B = 8'h5A; #100;
A = 8'hE0; B = 8'h5B; #100;
A = 8'hE0; B = 8'h5C; #100;
A = 8'hE0; B = 8'h5D; #100;
A = 8'hE0; B = 8'h5E; #100;
A = 8'hE0; B = 8'h5F; #100;
A = 8'hE0; B = 8'h60; #100;
A = 8'hE0; B = 8'h61; #100;
A = 8'hE0; B = 8'h62; #100;
A = 8'hE0; B = 8'h63; #100;
A = 8'hE0; B = 8'h64; #100;
A = 8'hE0; B = 8'h65; #100;
A = 8'hE0; B = 8'h66; #100;
A = 8'hE0; B = 8'h67; #100;
A = 8'hE0; B = 8'h68; #100;
A = 8'hE0; B = 8'h69; #100;
A = 8'hE0; B = 8'h6A; #100;
A = 8'hE0; B = 8'h6B; #100;
A = 8'hE0; B = 8'h6C; #100;
A = 8'hE0; B = 8'h6D; #100;
A = 8'hE0; B = 8'h6E; #100;
A = 8'hE0; B = 8'h6F; #100;
A = 8'hE0; B = 8'h70; #100;
A = 8'hE0; B = 8'h71; #100;
A = 8'hE0; B = 8'h72; #100;
A = 8'hE0; B = 8'h73; #100;
A = 8'hE0; B = 8'h74; #100;
A = 8'hE0; B = 8'h75; #100;
A = 8'hE0; B = 8'h76; #100;
A = 8'hE0; B = 8'h77; #100;
A = 8'hE0; B = 8'h78; #100;
A = 8'hE0; B = 8'h79; #100;
A = 8'hE0; B = 8'h7A; #100;
A = 8'hE0; B = 8'h7B; #100;
A = 8'hE0; B = 8'h7C; #100;
A = 8'hE0; B = 8'h7D; #100;
A = 8'hE0; B = 8'h7E; #100;
A = 8'hE0; B = 8'h7F; #100;
A = 8'hE0; B = 8'h80; #100;
A = 8'hE0; B = 8'h81; #100;
A = 8'hE0; B = 8'h82; #100;
A = 8'hE0; B = 8'h83; #100;
A = 8'hE0; B = 8'h84; #100;
A = 8'hE0; B = 8'h85; #100;
A = 8'hE0; B = 8'h86; #100;
A = 8'hE0; B = 8'h87; #100;
A = 8'hE0; B = 8'h88; #100;
A = 8'hE0; B = 8'h89; #100;
A = 8'hE0; B = 8'h8A; #100;
A = 8'hE0; B = 8'h8B; #100;
A = 8'hE0; B = 8'h8C; #100;
A = 8'hE0; B = 8'h8D; #100;
A = 8'hE0; B = 8'h8E; #100;
A = 8'hE0; B = 8'h8F; #100;
A = 8'hE0; B = 8'h90; #100;
A = 8'hE0; B = 8'h91; #100;
A = 8'hE0; B = 8'h92; #100;
A = 8'hE0; B = 8'h93; #100;
A = 8'hE0; B = 8'h94; #100;
A = 8'hE0; B = 8'h95; #100;
A = 8'hE0; B = 8'h96; #100;
A = 8'hE0; B = 8'h97; #100;
A = 8'hE0; B = 8'h98; #100;
A = 8'hE0; B = 8'h99; #100;
A = 8'hE0; B = 8'h9A; #100;
A = 8'hE0; B = 8'h9B; #100;
A = 8'hE0; B = 8'h9C; #100;
A = 8'hE0; B = 8'h9D; #100;
A = 8'hE0; B = 8'h9E; #100;
A = 8'hE0; B = 8'h9F; #100;
A = 8'hE0; B = 8'hA0; #100;
A = 8'hE0; B = 8'hA1; #100;
A = 8'hE0; B = 8'hA2; #100;
A = 8'hE0; B = 8'hA3; #100;
A = 8'hE0; B = 8'hA4; #100;
A = 8'hE0; B = 8'hA5; #100;
A = 8'hE0; B = 8'hA6; #100;
A = 8'hE0; B = 8'hA7; #100;
A = 8'hE0; B = 8'hA8; #100;
A = 8'hE0; B = 8'hA9; #100;
A = 8'hE0; B = 8'hAA; #100;
A = 8'hE0; B = 8'hAB; #100;
A = 8'hE0; B = 8'hAC; #100;
A = 8'hE0; B = 8'hAD; #100;
A = 8'hE0; B = 8'hAE; #100;
A = 8'hE0; B = 8'hAF; #100;
A = 8'hE0; B = 8'hB0; #100;
A = 8'hE0; B = 8'hB1; #100;
A = 8'hE0; B = 8'hB2; #100;
A = 8'hE0; B = 8'hB3; #100;
A = 8'hE0; B = 8'hB4; #100;
A = 8'hE0; B = 8'hB5; #100;
A = 8'hE0; B = 8'hB6; #100;
A = 8'hE0; B = 8'hB7; #100;
A = 8'hE0; B = 8'hB8; #100;
A = 8'hE0; B = 8'hB9; #100;
A = 8'hE0; B = 8'hBA; #100;
A = 8'hE0; B = 8'hBB; #100;
A = 8'hE0; B = 8'hBC; #100;
A = 8'hE0; B = 8'hBD; #100;
A = 8'hE0; B = 8'hBE; #100;
A = 8'hE0; B = 8'hBF; #100;
A = 8'hE0; B = 8'hC0; #100;
A = 8'hE0; B = 8'hC1; #100;
A = 8'hE0; B = 8'hC2; #100;
A = 8'hE0; B = 8'hC3; #100;
A = 8'hE0; B = 8'hC4; #100;
A = 8'hE0; B = 8'hC5; #100;
A = 8'hE0; B = 8'hC6; #100;
A = 8'hE0; B = 8'hC7; #100;
A = 8'hE0; B = 8'hC8; #100;
A = 8'hE0; B = 8'hC9; #100;
A = 8'hE0; B = 8'hCA; #100;
A = 8'hE0; B = 8'hCB; #100;
A = 8'hE0; B = 8'hCC; #100;
A = 8'hE0; B = 8'hCD; #100;
A = 8'hE0; B = 8'hCE; #100;
A = 8'hE0; B = 8'hCF; #100;
A = 8'hE0; B = 8'hD0; #100;
A = 8'hE0; B = 8'hD1; #100;
A = 8'hE0; B = 8'hD2; #100;
A = 8'hE0; B = 8'hD3; #100;
A = 8'hE0; B = 8'hD4; #100;
A = 8'hE0; B = 8'hD5; #100;
A = 8'hE0; B = 8'hD6; #100;
A = 8'hE0; B = 8'hD7; #100;
A = 8'hE0; B = 8'hD8; #100;
A = 8'hE0; B = 8'hD9; #100;
A = 8'hE0; B = 8'hDA; #100;
A = 8'hE0; B = 8'hDB; #100;
A = 8'hE0; B = 8'hDC; #100;
A = 8'hE0; B = 8'hDD; #100;
A = 8'hE0; B = 8'hDE; #100;
A = 8'hE0; B = 8'hDF; #100;
A = 8'hE0; B = 8'hE0; #100;
A = 8'hE0; B = 8'hE1; #100;
A = 8'hE0; B = 8'hE2; #100;
A = 8'hE0; B = 8'hE3; #100;
A = 8'hE0; B = 8'hE4; #100;
A = 8'hE0; B = 8'hE5; #100;
A = 8'hE0; B = 8'hE6; #100;
A = 8'hE0; B = 8'hE7; #100;
A = 8'hE0; B = 8'hE8; #100;
A = 8'hE0; B = 8'hE9; #100;
A = 8'hE0; B = 8'hEA; #100;
A = 8'hE0; B = 8'hEB; #100;
A = 8'hE0; B = 8'hEC; #100;
A = 8'hE0; B = 8'hED; #100;
A = 8'hE0; B = 8'hEE; #100;
A = 8'hE0; B = 8'hEF; #100;
A = 8'hE0; B = 8'hF0; #100;
A = 8'hE0; B = 8'hF1; #100;
A = 8'hE0; B = 8'hF2; #100;
A = 8'hE0; B = 8'hF3; #100;
A = 8'hE0; B = 8'hF4; #100;
A = 8'hE0; B = 8'hF5; #100;
A = 8'hE0; B = 8'hF6; #100;
A = 8'hE0; B = 8'hF7; #100;
A = 8'hE0; B = 8'hF8; #100;
A = 8'hE0; B = 8'hF9; #100;
A = 8'hE0; B = 8'hFA; #100;
A = 8'hE0; B = 8'hFB; #100;
A = 8'hE0; B = 8'hFC; #100;
A = 8'hE0; B = 8'hFD; #100;
A = 8'hE0; B = 8'hFE; #100;
A = 8'hE0; B = 8'hFF; #100;
A = 8'hE1; B = 8'h0; #100;
A = 8'hE1; B = 8'h1; #100;
A = 8'hE1; B = 8'h2; #100;
A = 8'hE1; B = 8'h3; #100;
A = 8'hE1; B = 8'h4; #100;
A = 8'hE1; B = 8'h5; #100;
A = 8'hE1; B = 8'h6; #100;
A = 8'hE1; B = 8'h7; #100;
A = 8'hE1; B = 8'h8; #100;
A = 8'hE1; B = 8'h9; #100;
A = 8'hE1; B = 8'hA; #100;
A = 8'hE1; B = 8'hB; #100;
A = 8'hE1; B = 8'hC; #100;
A = 8'hE1; B = 8'hD; #100;
A = 8'hE1; B = 8'hE; #100;
A = 8'hE1; B = 8'hF; #100;
A = 8'hE1; B = 8'h10; #100;
A = 8'hE1; B = 8'h11; #100;
A = 8'hE1; B = 8'h12; #100;
A = 8'hE1; B = 8'h13; #100;
A = 8'hE1; B = 8'h14; #100;
A = 8'hE1; B = 8'h15; #100;
A = 8'hE1; B = 8'h16; #100;
A = 8'hE1; B = 8'h17; #100;
A = 8'hE1; B = 8'h18; #100;
A = 8'hE1; B = 8'h19; #100;
A = 8'hE1; B = 8'h1A; #100;
A = 8'hE1; B = 8'h1B; #100;
A = 8'hE1; B = 8'h1C; #100;
A = 8'hE1; B = 8'h1D; #100;
A = 8'hE1; B = 8'h1E; #100;
A = 8'hE1; B = 8'h1F; #100;
A = 8'hE1; B = 8'h20; #100;
A = 8'hE1; B = 8'h21; #100;
A = 8'hE1; B = 8'h22; #100;
A = 8'hE1; B = 8'h23; #100;
A = 8'hE1; B = 8'h24; #100;
A = 8'hE1; B = 8'h25; #100;
A = 8'hE1; B = 8'h26; #100;
A = 8'hE1; B = 8'h27; #100;
A = 8'hE1; B = 8'h28; #100;
A = 8'hE1; B = 8'h29; #100;
A = 8'hE1; B = 8'h2A; #100;
A = 8'hE1; B = 8'h2B; #100;
A = 8'hE1; B = 8'h2C; #100;
A = 8'hE1; B = 8'h2D; #100;
A = 8'hE1; B = 8'h2E; #100;
A = 8'hE1; B = 8'h2F; #100;
A = 8'hE1; B = 8'h30; #100;
A = 8'hE1; B = 8'h31; #100;
A = 8'hE1; B = 8'h32; #100;
A = 8'hE1; B = 8'h33; #100;
A = 8'hE1; B = 8'h34; #100;
A = 8'hE1; B = 8'h35; #100;
A = 8'hE1; B = 8'h36; #100;
A = 8'hE1; B = 8'h37; #100;
A = 8'hE1; B = 8'h38; #100;
A = 8'hE1; B = 8'h39; #100;
A = 8'hE1; B = 8'h3A; #100;
A = 8'hE1; B = 8'h3B; #100;
A = 8'hE1; B = 8'h3C; #100;
A = 8'hE1; B = 8'h3D; #100;
A = 8'hE1; B = 8'h3E; #100;
A = 8'hE1; B = 8'h3F; #100;
A = 8'hE1; B = 8'h40; #100;
A = 8'hE1; B = 8'h41; #100;
A = 8'hE1; B = 8'h42; #100;
A = 8'hE1; B = 8'h43; #100;
A = 8'hE1; B = 8'h44; #100;
A = 8'hE1; B = 8'h45; #100;
A = 8'hE1; B = 8'h46; #100;
A = 8'hE1; B = 8'h47; #100;
A = 8'hE1; B = 8'h48; #100;
A = 8'hE1; B = 8'h49; #100;
A = 8'hE1; B = 8'h4A; #100;
A = 8'hE1; B = 8'h4B; #100;
A = 8'hE1; B = 8'h4C; #100;
A = 8'hE1; B = 8'h4D; #100;
A = 8'hE1; B = 8'h4E; #100;
A = 8'hE1; B = 8'h4F; #100;
A = 8'hE1; B = 8'h50; #100;
A = 8'hE1; B = 8'h51; #100;
A = 8'hE1; B = 8'h52; #100;
A = 8'hE1; B = 8'h53; #100;
A = 8'hE1; B = 8'h54; #100;
A = 8'hE1; B = 8'h55; #100;
A = 8'hE1; B = 8'h56; #100;
A = 8'hE1; B = 8'h57; #100;
A = 8'hE1; B = 8'h58; #100;
A = 8'hE1; B = 8'h59; #100;
A = 8'hE1; B = 8'h5A; #100;
A = 8'hE1; B = 8'h5B; #100;
A = 8'hE1; B = 8'h5C; #100;
A = 8'hE1; B = 8'h5D; #100;
A = 8'hE1; B = 8'h5E; #100;
A = 8'hE1; B = 8'h5F; #100;
A = 8'hE1; B = 8'h60; #100;
A = 8'hE1; B = 8'h61; #100;
A = 8'hE1; B = 8'h62; #100;
A = 8'hE1; B = 8'h63; #100;
A = 8'hE1; B = 8'h64; #100;
A = 8'hE1; B = 8'h65; #100;
A = 8'hE1; B = 8'h66; #100;
A = 8'hE1; B = 8'h67; #100;
A = 8'hE1; B = 8'h68; #100;
A = 8'hE1; B = 8'h69; #100;
A = 8'hE1; B = 8'h6A; #100;
A = 8'hE1; B = 8'h6B; #100;
A = 8'hE1; B = 8'h6C; #100;
A = 8'hE1; B = 8'h6D; #100;
A = 8'hE1; B = 8'h6E; #100;
A = 8'hE1; B = 8'h6F; #100;
A = 8'hE1; B = 8'h70; #100;
A = 8'hE1; B = 8'h71; #100;
A = 8'hE1; B = 8'h72; #100;
A = 8'hE1; B = 8'h73; #100;
A = 8'hE1; B = 8'h74; #100;
A = 8'hE1; B = 8'h75; #100;
A = 8'hE1; B = 8'h76; #100;
A = 8'hE1; B = 8'h77; #100;
A = 8'hE1; B = 8'h78; #100;
A = 8'hE1; B = 8'h79; #100;
A = 8'hE1; B = 8'h7A; #100;
A = 8'hE1; B = 8'h7B; #100;
A = 8'hE1; B = 8'h7C; #100;
A = 8'hE1; B = 8'h7D; #100;
A = 8'hE1; B = 8'h7E; #100;
A = 8'hE1; B = 8'h7F; #100;
A = 8'hE1; B = 8'h80; #100;
A = 8'hE1; B = 8'h81; #100;
A = 8'hE1; B = 8'h82; #100;
A = 8'hE1; B = 8'h83; #100;
A = 8'hE1; B = 8'h84; #100;
A = 8'hE1; B = 8'h85; #100;
A = 8'hE1; B = 8'h86; #100;
A = 8'hE1; B = 8'h87; #100;
A = 8'hE1; B = 8'h88; #100;
A = 8'hE1; B = 8'h89; #100;
A = 8'hE1; B = 8'h8A; #100;
A = 8'hE1; B = 8'h8B; #100;
A = 8'hE1; B = 8'h8C; #100;
A = 8'hE1; B = 8'h8D; #100;
A = 8'hE1; B = 8'h8E; #100;
A = 8'hE1; B = 8'h8F; #100;
A = 8'hE1; B = 8'h90; #100;
A = 8'hE1; B = 8'h91; #100;
A = 8'hE1; B = 8'h92; #100;
A = 8'hE1; B = 8'h93; #100;
A = 8'hE1; B = 8'h94; #100;
A = 8'hE1; B = 8'h95; #100;
A = 8'hE1; B = 8'h96; #100;
A = 8'hE1; B = 8'h97; #100;
A = 8'hE1; B = 8'h98; #100;
A = 8'hE1; B = 8'h99; #100;
A = 8'hE1; B = 8'h9A; #100;
A = 8'hE1; B = 8'h9B; #100;
A = 8'hE1; B = 8'h9C; #100;
A = 8'hE1; B = 8'h9D; #100;
A = 8'hE1; B = 8'h9E; #100;
A = 8'hE1; B = 8'h9F; #100;
A = 8'hE1; B = 8'hA0; #100;
A = 8'hE1; B = 8'hA1; #100;
A = 8'hE1; B = 8'hA2; #100;
A = 8'hE1; B = 8'hA3; #100;
A = 8'hE1; B = 8'hA4; #100;
A = 8'hE1; B = 8'hA5; #100;
A = 8'hE1; B = 8'hA6; #100;
A = 8'hE1; B = 8'hA7; #100;
A = 8'hE1; B = 8'hA8; #100;
A = 8'hE1; B = 8'hA9; #100;
A = 8'hE1; B = 8'hAA; #100;
A = 8'hE1; B = 8'hAB; #100;
A = 8'hE1; B = 8'hAC; #100;
A = 8'hE1; B = 8'hAD; #100;
A = 8'hE1; B = 8'hAE; #100;
A = 8'hE1; B = 8'hAF; #100;
A = 8'hE1; B = 8'hB0; #100;
A = 8'hE1; B = 8'hB1; #100;
A = 8'hE1; B = 8'hB2; #100;
A = 8'hE1; B = 8'hB3; #100;
A = 8'hE1; B = 8'hB4; #100;
A = 8'hE1; B = 8'hB5; #100;
A = 8'hE1; B = 8'hB6; #100;
A = 8'hE1; B = 8'hB7; #100;
A = 8'hE1; B = 8'hB8; #100;
A = 8'hE1; B = 8'hB9; #100;
A = 8'hE1; B = 8'hBA; #100;
A = 8'hE1; B = 8'hBB; #100;
A = 8'hE1; B = 8'hBC; #100;
A = 8'hE1; B = 8'hBD; #100;
A = 8'hE1; B = 8'hBE; #100;
A = 8'hE1; B = 8'hBF; #100;
A = 8'hE1; B = 8'hC0; #100;
A = 8'hE1; B = 8'hC1; #100;
A = 8'hE1; B = 8'hC2; #100;
A = 8'hE1; B = 8'hC3; #100;
A = 8'hE1; B = 8'hC4; #100;
A = 8'hE1; B = 8'hC5; #100;
A = 8'hE1; B = 8'hC6; #100;
A = 8'hE1; B = 8'hC7; #100;
A = 8'hE1; B = 8'hC8; #100;
A = 8'hE1; B = 8'hC9; #100;
A = 8'hE1; B = 8'hCA; #100;
A = 8'hE1; B = 8'hCB; #100;
A = 8'hE1; B = 8'hCC; #100;
A = 8'hE1; B = 8'hCD; #100;
A = 8'hE1; B = 8'hCE; #100;
A = 8'hE1; B = 8'hCF; #100;
A = 8'hE1; B = 8'hD0; #100;
A = 8'hE1; B = 8'hD1; #100;
A = 8'hE1; B = 8'hD2; #100;
A = 8'hE1; B = 8'hD3; #100;
A = 8'hE1; B = 8'hD4; #100;
A = 8'hE1; B = 8'hD5; #100;
A = 8'hE1; B = 8'hD6; #100;
A = 8'hE1; B = 8'hD7; #100;
A = 8'hE1; B = 8'hD8; #100;
A = 8'hE1; B = 8'hD9; #100;
A = 8'hE1; B = 8'hDA; #100;
A = 8'hE1; B = 8'hDB; #100;
A = 8'hE1; B = 8'hDC; #100;
A = 8'hE1; B = 8'hDD; #100;
A = 8'hE1; B = 8'hDE; #100;
A = 8'hE1; B = 8'hDF; #100;
A = 8'hE1; B = 8'hE0; #100;
A = 8'hE1; B = 8'hE1; #100;
A = 8'hE1; B = 8'hE2; #100;
A = 8'hE1; B = 8'hE3; #100;
A = 8'hE1; B = 8'hE4; #100;
A = 8'hE1; B = 8'hE5; #100;
A = 8'hE1; B = 8'hE6; #100;
A = 8'hE1; B = 8'hE7; #100;
A = 8'hE1; B = 8'hE8; #100;
A = 8'hE1; B = 8'hE9; #100;
A = 8'hE1; B = 8'hEA; #100;
A = 8'hE1; B = 8'hEB; #100;
A = 8'hE1; B = 8'hEC; #100;
A = 8'hE1; B = 8'hED; #100;
A = 8'hE1; B = 8'hEE; #100;
A = 8'hE1; B = 8'hEF; #100;
A = 8'hE1; B = 8'hF0; #100;
A = 8'hE1; B = 8'hF1; #100;
A = 8'hE1; B = 8'hF2; #100;
A = 8'hE1; B = 8'hF3; #100;
A = 8'hE1; B = 8'hF4; #100;
A = 8'hE1; B = 8'hF5; #100;
A = 8'hE1; B = 8'hF6; #100;
A = 8'hE1; B = 8'hF7; #100;
A = 8'hE1; B = 8'hF8; #100;
A = 8'hE1; B = 8'hF9; #100;
A = 8'hE1; B = 8'hFA; #100;
A = 8'hE1; B = 8'hFB; #100;
A = 8'hE1; B = 8'hFC; #100;
A = 8'hE1; B = 8'hFD; #100;
A = 8'hE1; B = 8'hFE; #100;
A = 8'hE1; B = 8'hFF; #100;
A = 8'hE2; B = 8'h0; #100;
A = 8'hE2; B = 8'h1; #100;
A = 8'hE2; B = 8'h2; #100;
A = 8'hE2; B = 8'h3; #100;
A = 8'hE2; B = 8'h4; #100;
A = 8'hE2; B = 8'h5; #100;
A = 8'hE2; B = 8'h6; #100;
A = 8'hE2; B = 8'h7; #100;
A = 8'hE2; B = 8'h8; #100;
A = 8'hE2; B = 8'h9; #100;
A = 8'hE2; B = 8'hA; #100;
A = 8'hE2; B = 8'hB; #100;
A = 8'hE2; B = 8'hC; #100;
A = 8'hE2; B = 8'hD; #100;
A = 8'hE2; B = 8'hE; #100;
A = 8'hE2; B = 8'hF; #100;
A = 8'hE2; B = 8'h10; #100;
A = 8'hE2; B = 8'h11; #100;
A = 8'hE2; B = 8'h12; #100;
A = 8'hE2; B = 8'h13; #100;
A = 8'hE2; B = 8'h14; #100;
A = 8'hE2; B = 8'h15; #100;
A = 8'hE2; B = 8'h16; #100;
A = 8'hE2; B = 8'h17; #100;
A = 8'hE2; B = 8'h18; #100;
A = 8'hE2; B = 8'h19; #100;
A = 8'hE2; B = 8'h1A; #100;
A = 8'hE2; B = 8'h1B; #100;
A = 8'hE2; B = 8'h1C; #100;
A = 8'hE2; B = 8'h1D; #100;
A = 8'hE2; B = 8'h1E; #100;
A = 8'hE2; B = 8'h1F; #100;
A = 8'hE2; B = 8'h20; #100;
A = 8'hE2; B = 8'h21; #100;
A = 8'hE2; B = 8'h22; #100;
A = 8'hE2; B = 8'h23; #100;
A = 8'hE2; B = 8'h24; #100;
A = 8'hE2; B = 8'h25; #100;
A = 8'hE2; B = 8'h26; #100;
A = 8'hE2; B = 8'h27; #100;
A = 8'hE2; B = 8'h28; #100;
A = 8'hE2; B = 8'h29; #100;
A = 8'hE2; B = 8'h2A; #100;
A = 8'hE2; B = 8'h2B; #100;
A = 8'hE2; B = 8'h2C; #100;
A = 8'hE2; B = 8'h2D; #100;
A = 8'hE2; B = 8'h2E; #100;
A = 8'hE2; B = 8'h2F; #100;
A = 8'hE2; B = 8'h30; #100;
A = 8'hE2; B = 8'h31; #100;
A = 8'hE2; B = 8'h32; #100;
A = 8'hE2; B = 8'h33; #100;
A = 8'hE2; B = 8'h34; #100;
A = 8'hE2; B = 8'h35; #100;
A = 8'hE2; B = 8'h36; #100;
A = 8'hE2; B = 8'h37; #100;
A = 8'hE2; B = 8'h38; #100;
A = 8'hE2; B = 8'h39; #100;
A = 8'hE2; B = 8'h3A; #100;
A = 8'hE2; B = 8'h3B; #100;
A = 8'hE2; B = 8'h3C; #100;
A = 8'hE2; B = 8'h3D; #100;
A = 8'hE2; B = 8'h3E; #100;
A = 8'hE2; B = 8'h3F; #100;
A = 8'hE2; B = 8'h40; #100;
A = 8'hE2; B = 8'h41; #100;
A = 8'hE2; B = 8'h42; #100;
A = 8'hE2; B = 8'h43; #100;
A = 8'hE2; B = 8'h44; #100;
A = 8'hE2; B = 8'h45; #100;
A = 8'hE2; B = 8'h46; #100;
A = 8'hE2; B = 8'h47; #100;
A = 8'hE2; B = 8'h48; #100;
A = 8'hE2; B = 8'h49; #100;
A = 8'hE2; B = 8'h4A; #100;
A = 8'hE2; B = 8'h4B; #100;
A = 8'hE2; B = 8'h4C; #100;
A = 8'hE2; B = 8'h4D; #100;
A = 8'hE2; B = 8'h4E; #100;
A = 8'hE2; B = 8'h4F; #100;
A = 8'hE2; B = 8'h50; #100;
A = 8'hE2; B = 8'h51; #100;
A = 8'hE2; B = 8'h52; #100;
A = 8'hE2; B = 8'h53; #100;
A = 8'hE2; B = 8'h54; #100;
A = 8'hE2; B = 8'h55; #100;
A = 8'hE2; B = 8'h56; #100;
A = 8'hE2; B = 8'h57; #100;
A = 8'hE2; B = 8'h58; #100;
A = 8'hE2; B = 8'h59; #100;
A = 8'hE2; B = 8'h5A; #100;
A = 8'hE2; B = 8'h5B; #100;
A = 8'hE2; B = 8'h5C; #100;
A = 8'hE2; B = 8'h5D; #100;
A = 8'hE2; B = 8'h5E; #100;
A = 8'hE2; B = 8'h5F; #100;
A = 8'hE2; B = 8'h60; #100;
A = 8'hE2; B = 8'h61; #100;
A = 8'hE2; B = 8'h62; #100;
A = 8'hE2; B = 8'h63; #100;
A = 8'hE2; B = 8'h64; #100;
A = 8'hE2; B = 8'h65; #100;
A = 8'hE2; B = 8'h66; #100;
A = 8'hE2; B = 8'h67; #100;
A = 8'hE2; B = 8'h68; #100;
A = 8'hE2; B = 8'h69; #100;
A = 8'hE2; B = 8'h6A; #100;
A = 8'hE2; B = 8'h6B; #100;
A = 8'hE2; B = 8'h6C; #100;
A = 8'hE2; B = 8'h6D; #100;
A = 8'hE2; B = 8'h6E; #100;
A = 8'hE2; B = 8'h6F; #100;
A = 8'hE2; B = 8'h70; #100;
A = 8'hE2; B = 8'h71; #100;
A = 8'hE2; B = 8'h72; #100;
A = 8'hE2; B = 8'h73; #100;
A = 8'hE2; B = 8'h74; #100;
A = 8'hE2; B = 8'h75; #100;
A = 8'hE2; B = 8'h76; #100;
A = 8'hE2; B = 8'h77; #100;
A = 8'hE2; B = 8'h78; #100;
A = 8'hE2; B = 8'h79; #100;
A = 8'hE2; B = 8'h7A; #100;
A = 8'hE2; B = 8'h7B; #100;
A = 8'hE2; B = 8'h7C; #100;
A = 8'hE2; B = 8'h7D; #100;
A = 8'hE2; B = 8'h7E; #100;
A = 8'hE2; B = 8'h7F; #100;
A = 8'hE2; B = 8'h80; #100;
A = 8'hE2; B = 8'h81; #100;
A = 8'hE2; B = 8'h82; #100;
A = 8'hE2; B = 8'h83; #100;
A = 8'hE2; B = 8'h84; #100;
A = 8'hE2; B = 8'h85; #100;
A = 8'hE2; B = 8'h86; #100;
A = 8'hE2; B = 8'h87; #100;
A = 8'hE2; B = 8'h88; #100;
A = 8'hE2; B = 8'h89; #100;
A = 8'hE2; B = 8'h8A; #100;
A = 8'hE2; B = 8'h8B; #100;
A = 8'hE2; B = 8'h8C; #100;
A = 8'hE2; B = 8'h8D; #100;
A = 8'hE2; B = 8'h8E; #100;
A = 8'hE2; B = 8'h8F; #100;
A = 8'hE2; B = 8'h90; #100;
A = 8'hE2; B = 8'h91; #100;
A = 8'hE2; B = 8'h92; #100;
A = 8'hE2; B = 8'h93; #100;
A = 8'hE2; B = 8'h94; #100;
A = 8'hE2; B = 8'h95; #100;
A = 8'hE2; B = 8'h96; #100;
A = 8'hE2; B = 8'h97; #100;
A = 8'hE2; B = 8'h98; #100;
A = 8'hE2; B = 8'h99; #100;
A = 8'hE2; B = 8'h9A; #100;
A = 8'hE2; B = 8'h9B; #100;
A = 8'hE2; B = 8'h9C; #100;
A = 8'hE2; B = 8'h9D; #100;
A = 8'hE2; B = 8'h9E; #100;
A = 8'hE2; B = 8'h9F; #100;
A = 8'hE2; B = 8'hA0; #100;
A = 8'hE2; B = 8'hA1; #100;
A = 8'hE2; B = 8'hA2; #100;
A = 8'hE2; B = 8'hA3; #100;
A = 8'hE2; B = 8'hA4; #100;
A = 8'hE2; B = 8'hA5; #100;
A = 8'hE2; B = 8'hA6; #100;
A = 8'hE2; B = 8'hA7; #100;
A = 8'hE2; B = 8'hA8; #100;
A = 8'hE2; B = 8'hA9; #100;
A = 8'hE2; B = 8'hAA; #100;
A = 8'hE2; B = 8'hAB; #100;
A = 8'hE2; B = 8'hAC; #100;
A = 8'hE2; B = 8'hAD; #100;
A = 8'hE2; B = 8'hAE; #100;
A = 8'hE2; B = 8'hAF; #100;
A = 8'hE2; B = 8'hB0; #100;
A = 8'hE2; B = 8'hB1; #100;
A = 8'hE2; B = 8'hB2; #100;
A = 8'hE2; B = 8'hB3; #100;
A = 8'hE2; B = 8'hB4; #100;
A = 8'hE2; B = 8'hB5; #100;
A = 8'hE2; B = 8'hB6; #100;
A = 8'hE2; B = 8'hB7; #100;
A = 8'hE2; B = 8'hB8; #100;
A = 8'hE2; B = 8'hB9; #100;
A = 8'hE2; B = 8'hBA; #100;
A = 8'hE2; B = 8'hBB; #100;
A = 8'hE2; B = 8'hBC; #100;
A = 8'hE2; B = 8'hBD; #100;
A = 8'hE2; B = 8'hBE; #100;
A = 8'hE2; B = 8'hBF; #100;
A = 8'hE2; B = 8'hC0; #100;
A = 8'hE2; B = 8'hC1; #100;
A = 8'hE2; B = 8'hC2; #100;
A = 8'hE2; B = 8'hC3; #100;
A = 8'hE2; B = 8'hC4; #100;
A = 8'hE2; B = 8'hC5; #100;
A = 8'hE2; B = 8'hC6; #100;
A = 8'hE2; B = 8'hC7; #100;
A = 8'hE2; B = 8'hC8; #100;
A = 8'hE2; B = 8'hC9; #100;
A = 8'hE2; B = 8'hCA; #100;
A = 8'hE2; B = 8'hCB; #100;
A = 8'hE2; B = 8'hCC; #100;
A = 8'hE2; B = 8'hCD; #100;
A = 8'hE2; B = 8'hCE; #100;
A = 8'hE2; B = 8'hCF; #100;
A = 8'hE2; B = 8'hD0; #100;
A = 8'hE2; B = 8'hD1; #100;
A = 8'hE2; B = 8'hD2; #100;
A = 8'hE2; B = 8'hD3; #100;
A = 8'hE2; B = 8'hD4; #100;
A = 8'hE2; B = 8'hD5; #100;
A = 8'hE2; B = 8'hD6; #100;
A = 8'hE2; B = 8'hD7; #100;
A = 8'hE2; B = 8'hD8; #100;
A = 8'hE2; B = 8'hD9; #100;
A = 8'hE2; B = 8'hDA; #100;
A = 8'hE2; B = 8'hDB; #100;
A = 8'hE2; B = 8'hDC; #100;
A = 8'hE2; B = 8'hDD; #100;
A = 8'hE2; B = 8'hDE; #100;
A = 8'hE2; B = 8'hDF; #100;
A = 8'hE2; B = 8'hE0; #100;
A = 8'hE2; B = 8'hE1; #100;
A = 8'hE2; B = 8'hE2; #100;
A = 8'hE2; B = 8'hE3; #100;
A = 8'hE2; B = 8'hE4; #100;
A = 8'hE2; B = 8'hE5; #100;
A = 8'hE2; B = 8'hE6; #100;
A = 8'hE2; B = 8'hE7; #100;
A = 8'hE2; B = 8'hE8; #100;
A = 8'hE2; B = 8'hE9; #100;
A = 8'hE2; B = 8'hEA; #100;
A = 8'hE2; B = 8'hEB; #100;
A = 8'hE2; B = 8'hEC; #100;
A = 8'hE2; B = 8'hED; #100;
A = 8'hE2; B = 8'hEE; #100;
A = 8'hE2; B = 8'hEF; #100;
A = 8'hE2; B = 8'hF0; #100;
A = 8'hE2; B = 8'hF1; #100;
A = 8'hE2; B = 8'hF2; #100;
A = 8'hE2; B = 8'hF3; #100;
A = 8'hE2; B = 8'hF4; #100;
A = 8'hE2; B = 8'hF5; #100;
A = 8'hE2; B = 8'hF6; #100;
A = 8'hE2; B = 8'hF7; #100;
A = 8'hE2; B = 8'hF8; #100;
A = 8'hE2; B = 8'hF9; #100;
A = 8'hE2; B = 8'hFA; #100;
A = 8'hE2; B = 8'hFB; #100;
A = 8'hE2; B = 8'hFC; #100;
A = 8'hE2; B = 8'hFD; #100;
A = 8'hE2; B = 8'hFE; #100;
A = 8'hE2; B = 8'hFF; #100;
A = 8'hE3; B = 8'h0; #100;
A = 8'hE3; B = 8'h1; #100;
A = 8'hE3; B = 8'h2; #100;
A = 8'hE3; B = 8'h3; #100;
A = 8'hE3; B = 8'h4; #100;
A = 8'hE3; B = 8'h5; #100;
A = 8'hE3; B = 8'h6; #100;
A = 8'hE3; B = 8'h7; #100;
A = 8'hE3; B = 8'h8; #100;
A = 8'hE3; B = 8'h9; #100;
A = 8'hE3; B = 8'hA; #100;
A = 8'hE3; B = 8'hB; #100;
A = 8'hE3; B = 8'hC; #100;
A = 8'hE3; B = 8'hD; #100;
A = 8'hE3; B = 8'hE; #100;
A = 8'hE3; B = 8'hF; #100;
A = 8'hE3; B = 8'h10; #100;
A = 8'hE3; B = 8'h11; #100;
A = 8'hE3; B = 8'h12; #100;
A = 8'hE3; B = 8'h13; #100;
A = 8'hE3; B = 8'h14; #100;
A = 8'hE3; B = 8'h15; #100;
A = 8'hE3; B = 8'h16; #100;
A = 8'hE3; B = 8'h17; #100;
A = 8'hE3; B = 8'h18; #100;
A = 8'hE3; B = 8'h19; #100;
A = 8'hE3; B = 8'h1A; #100;
A = 8'hE3; B = 8'h1B; #100;
A = 8'hE3; B = 8'h1C; #100;
A = 8'hE3; B = 8'h1D; #100;
A = 8'hE3; B = 8'h1E; #100;
A = 8'hE3; B = 8'h1F; #100;
A = 8'hE3; B = 8'h20; #100;
A = 8'hE3; B = 8'h21; #100;
A = 8'hE3; B = 8'h22; #100;
A = 8'hE3; B = 8'h23; #100;
A = 8'hE3; B = 8'h24; #100;
A = 8'hE3; B = 8'h25; #100;
A = 8'hE3; B = 8'h26; #100;
A = 8'hE3; B = 8'h27; #100;
A = 8'hE3; B = 8'h28; #100;
A = 8'hE3; B = 8'h29; #100;
A = 8'hE3; B = 8'h2A; #100;
A = 8'hE3; B = 8'h2B; #100;
A = 8'hE3; B = 8'h2C; #100;
A = 8'hE3; B = 8'h2D; #100;
A = 8'hE3; B = 8'h2E; #100;
A = 8'hE3; B = 8'h2F; #100;
A = 8'hE3; B = 8'h30; #100;
A = 8'hE3; B = 8'h31; #100;
A = 8'hE3; B = 8'h32; #100;
A = 8'hE3; B = 8'h33; #100;
A = 8'hE3; B = 8'h34; #100;
A = 8'hE3; B = 8'h35; #100;
A = 8'hE3; B = 8'h36; #100;
A = 8'hE3; B = 8'h37; #100;
A = 8'hE3; B = 8'h38; #100;
A = 8'hE3; B = 8'h39; #100;
A = 8'hE3; B = 8'h3A; #100;
A = 8'hE3; B = 8'h3B; #100;
A = 8'hE3; B = 8'h3C; #100;
A = 8'hE3; B = 8'h3D; #100;
A = 8'hE3; B = 8'h3E; #100;
A = 8'hE3; B = 8'h3F; #100;
A = 8'hE3; B = 8'h40; #100;
A = 8'hE3; B = 8'h41; #100;
A = 8'hE3; B = 8'h42; #100;
A = 8'hE3; B = 8'h43; #100;
A = 8'hE3; B = 8'h44; #100;
A = 8'hE3; B = 8'h45; #100;
A = 8'hE3; B = 8'h46; #100;
A = 8'hE3; B = 8'h47; #100;
A = 8'hE3; B = 8'h48; #100;
A = 8'hE3; B = 8'h49; #100;
A = 8'hE3; B = 8'h4A; #100;
A = 8'hE3; B = 8'h4B; #100;
A = 8'hE3; B = 8'h4C; #100;
A = 8'hE3; B = 8'h4D; #100;
A = 8'hE3; B = 8'h4E; #100;
A = 8'hE3; B = 8'h4F; #100;
A = 8'hE3; B = 8'h50; #100;
A = 8'hE3; B = 8'h51; #100;
A = 8'hE3; B = 8'h52; #100;
A = 8'hE3; B = 8'h53; #100;
A = 8'hE3; B = 8'h54; #100;
A = 8'hE3; B = 8'h55; #100;
A = 8'hE3; B = 8'h56; #100;
A = 8'hE3; B = 8'h57; #100;
A = 8'hE3; B = 8'h58; #100;
A = 8'hE3; B = 8'h59; #100;
A = 8'hE3; B = 8'h5A; #100;
A = 8'hE3; B = 8'h5B; #100;
A = 8'hE3; B = 8'h5C; #100;
A = 8'hE3; B = 8'h5D; #100;
A = 8'hE3; B = 8'h5E; #100;
A = 8'hE3; B = 8'h5F; #100;
A = 8'hE3; B = 8'h60; #100;
A = 8'hE3; B = 8'h61; #100;
A = 8'hE3; B = 8'h62; #100;
A = 8'hE3; B = 8'h63; #100;
A = 8'hE3; B = 8'h64; #100;
A = 8'hE3; B = 8'h65; #100;
A = 8'hE3; B = 8'h66; #100;
A = 8'hE3; B = 8'h67; #100;
A = 8'hE3; B = 8'h68; #100;
A = 8'hE3; B = 8'h69; #100;
A = 8'hE3; B = 8'h6A; #100;
A = 8'hE3; B = 8'h6B; #100;
A = 8'hE3; B = 8'h6C; #100;
A = 8'hE3; B = 8'h6D; #100;
A = 8'hE3; B = 8'h6E; #100;
A = 8'hE3; B = 8'h6F; #100;
A = 8'hE3; B = 8'h70; #100;
A = 8'hE3; B = 8'h71; #100;
A = 8'hE3; B = 8'h72; #100;
A = 8'hE3; B = 8'h73; #100;
A = 8'hE3; B = 8'h74; #100;
A = 8'hE3; B = 8'h75; #100;
A = 8'hE3; B = 8'h76; #100;
A = 8'hE3; B = 8'h77; #100;
A = 8'hE3; B = 8'h78; #100;
A = 8'hE3; B = 8'h79; #100;
A = 8'hE3; B = 8'h7A; #100;
A = 8'hE3; B = 8'h7B; #100;
A = 8'hE3; B = 8'h7C; #100;
A = 8'hE3; B = 8'h7D; #100;
A = 8'hE3; B = 8'h7E; #100;
A = 8'hE3; B = 8'h7F; #100;
A = 8'hE3; B = 8'h80; #100;
A = 8'hE3; B = 8'h81; #100;
A = 8'hE3; B = 8'h82; #100;
A = 8'hE3; B = 8'h83; #100;
A = 8'hE3; B = 8'h84; #100;
A = 8'hE3; B = 8'h85; #100;
A = 8'hE3; B = 8'h86; #100;
A = 8'hE3; B = 8'h87; #100;
A = 8'hE3; B = 8'h88; #100;
A = 8'hE3; B = 8'h89; #100;
A = 8'hE3; B = 8'h8A; #100;
A = 8'hE3; B = 8'h8B; #100;
A = 8'hE3; B = 8'h8C; #100;
A = 8'hE3; B = 8'h8D; #100;
A = 8'hE3; B = 8'h8E; #100;
A = 8'hE3; B = 8'h8F; #100;
A = 8'hE3; B = 8'h90; #100;
A = 8'hE3; B = 8'h91; #100;
A = 8'hE3; B = 8'h92; #100;
A = 8'hE3; B = 8'h93; #100;
A = 8'hE3; B = 8'h94; #100;
A = 8'hE3; B = 8'h95; #100;
A = 8'hE3; B = 8'h96; #100;
A = 8'hE3; B = 8'h97; #100;
A = 8'hE3; B = 8'h98; #100;
A = 8'hE3; B = 8'h99; #100;
A = 8'hE3; B = 8'h9A; #100;
A = 8'hE3; B = 8'h9B; #100;
A = 8'hE3; B = 8'h9C; #100;
A = 8'hE3; B = 8'h9D; #100;
A = 8'hE3; B = 8'h9E; #100;
A = 8'hE3; B = 8'h9F; #100;
A = 8'hE3; B = 8'hA0; #100;
A = 8'hE3; B = 8'hA1; #100;
A = 8'hE3; B = 8'hA2; #100;
A = 8'hE3; B = 8'hA3; #100;
A = 8'hE3; B = 8'hA4; #100;
A = 8'hE3; B = 8'hA5; #100;
A = 8'hE3; B = 8'hA6; #100;
A = 8'hE3; B = 8'hA7; #100;
A = 8'hE3; B = 8'hA8; #100;
A = 8'hE3; B = 8'hA9; #100;
A = 8'hE3; B = 8'hAA; #100;
A = 8'hE3; B = 8'hAB; #100;
A = 8'hE3; B = 8'hAC; #100;
A = 8'hE3; B = 8'hAD; #100;
A = 8'hE3; B = 8'hAE; #100;
A = 8'hE3; B = 8'hAF; #100;
A = 8'hE3; B = 8'hB0; #100;
A = 8'hE3; B = 8'hB1; #100;
A = 8'hE3; B = 8'hB2; #100;
A = 8'hE3; B = 8'hB3; #100;
A = 8'hE3; B = 8'hB4; #100;
A = 8'hE3; B = 8'hB5; #100;
A = 8'hE3; B = 8'hB6; #100;
A = 8'hE3; B = 8'hB7; #100;
A = 8'hE3; B = 8'hB8; #100;
A = 8'hE3; B = 8'hB9; #100;
A = 8'hE3; B = 8'hBA; #100;
A = 8'hE3; B = 8'hBB; #100;
A = 8'hE3; B = 8'hBC; #100;
A = 8'hE3; B = 8'hBD; #100;
A = 8'hE3; B = 8'hBE; #100;
A = 8'hE3; B = 8'hBF; #100;
A = 8'hE3; B = 8'hC0; #100;
A = 8'hE3; B = 8'hC1; #100;
A = 8'hE3; B = 8'hC2; #100;
A = 8'hE3; B = 8'hC3; #100;
A = 8'hE3; B = 8'hC4; #100;
A = 8'hE3; B = 8'hC5; #100;
A = 8'hE3; B = 8'hC6; #100;
A = 8'hE3; B = 8'hC7; #100;
A = 8'hE3; B = 8'hC8; #100;
A = 8'hE3; B = 8'hC9; #100;
A = 8'hE3; B = 8'hCA; #100;
A = 8'hE3; B = 8'hCB; #100;
A = 8'hE3; B = 8'hCC; #100;
A = 8'hE3; B = 8'hCD; #100;
A = 8'hE3; B = 8'hCE; #100;
A = 8'hE3; B = 8'hCF; #100;
A = 8'hE3; B = 8'hD0; #100;
A = 8'hE3; B = 8'hD1; #100;
A = 8'hE3; B = 8'hD2; #100;
A = 8'hE3; B = 8'hD3; #100;
A = 8'hE3; B = 8'hD4; #100;
A = 8'hE3; B = 8'hD5; #100;
A = 8'hE3; B = 8'hD6; #100;
A = 8'hE3; B = 8'hD7; #100;
A = 8'hE3; B = 8'hD8; #100;
A = 8'hE3; B = 8'hD9; #100;
A = 8'hE3; B = 8'hDA; #100;
A = 8'hE3; B = 8'hDB; #100;
A = 8'hE3; B = 8'hDC; #100;
A = 8'hE3; B = 8'hDD; #100;
A = 8'hE3; B = 8'hDE; #100;
A = 8'hE3; B = 8'hDF; #100;
A = 8'hE3; B = 8'hE0; #100;
A = 8'hE3; B = 8'hE1; #100;
A = 8'hE3; B = 8'hE2; #100;
A = 8'hE3; B = 8'hE3; #100;
A = 8'hE3; B = 8'hE4; #100;
A = 8'hE3; B = 8'hE5; #100;
A = 8'hE3; B = 8'hE6; #100;
A = 8'hE3; B = 8'hE7; #100;
A = 8'hE3; B = 8'hE8; #100;
A = 8'hE3; B = 8'hE9; #100;
A = 8'hE3; B = 8'hEA; #100;
A = 8'hE3; B = 8'hEB; #100;
A = 8'hE3; B = 8'hEC; #100;
A = 8'hE3; B = 8'hED; #100;
A = 8'hE3; B = 8'hEE; #100;
A = 8'hE3; B = 8'hEF; #100;
A = 8'hE3; B = 8'hF0; #100;
A = 8'hE3; B = 8'hF1; #100;
A = 8'hE3; B = 8'hF2; #100;
A = 8'hE3; B = 8'hF3; #100;
A = 8'hE3; B = 8'hF4; #100;
A = 8'hE3; B = 8'hF5; #100;
A = 8'hE3; B = 8'hF6; #100;
A = 8'hE3; B = 8'hF7; #100;
A = 8'hE3; B = 8'hF8; #100;
A = 8'hE3; B = 8'hF9; #100;
A = 8'hE3; B = 8'hFA; #100;
A = 8'hE3; B = 8'hFB; #100;
A = 8'hE3; B = 8'hFC; #100;
A = 8'hE3; B = 8'hFD; #100;
A = 8'hE3; B = 8'hFE; #100;
A = 8'hE3; B = 8'hFF; #100;
A = 8'hE4; B = 8'h0; #100;
A = 8'hE4; B = 8'h1; #100;
A = 8'hE4; B = 8'h2; #100;
A = 8'hE4; B = 8'h3; #100;
A = 8'hE4; B = 8'h4; #100;
A = 8'hE4; B = 8'h5; #100;
A = 8'hE4; B = 8'h6; #100;
A = 8'hE4; B = 8'h7; #100;
A = 8'hE4; B = 8'h8; #100;
A = 8'hE4; B = 8'h9; #100;
A = 8'hE4; B = 8'hA; #100;
A = 8'hE4; B = 8'hB; #100;
A = 8'hE4; B = 8'hC; #100;
A = 8'hE4; B = 8'hD; #100;
A = 8'hE4; B = 8'hE; #100;
A = 8'hE4; B = 8'hF; #100;
A = 8'hE4; B = 8'h10; #100;
A = 8'hE4; B = 8'h11; #100;
A = 8'hE4; B = 8'h12; #100;
A = 8'hE4; B = 8'h13; #100;
A = 8'hE4; B = 8'h14; #100;
A = 8'hE4; B = 8'h15; #100;
A = 8'hE4; B = 8'h16; #100;
A = 8'hE4; B = 8'h17; #100;
A = 8'hE4; B = 8'h18; #100;
A = 8'hE4; B = 8'h19; #100;
A = 8'hE4; B = 8'h1A; #100;
A = 8'hE4; B = 8'h1B; #100;
A = 8'hE4; B = 8'h1C; #100;
A = 8'hE4; B = 8'h1D; #100;
A = 8'hE4; B = 8'h1E; #100;
A = 8'hE4; B = 8'h1F; #100;
A = 8'hE4; B = 8'h20; #100;
A = 8'hE4; B = 8'h21; #100;
A = 8'hE4; B = 8'h22; #100;
A = 8'hE4; B = 8'h23; #100;
A = 8'hE4; B = 8'h24; #100;
A = 8'hE4; B = 8'h25; #100;
A = 8'hE4; B = 8'h26; #100;
A = 8'hE4; B = 8'h27; #100;
A = 8'hE4; B = 8'h28; #100;
A = 8'hE4; B = 8'h29; #100;
A = 8'hE4; B = 8'h2A; #100;
A = 8'hE4; B = 8'h2B; #100;
A = 8'hE4; B = 8'h2C; #100;
A = 8'hE4; B = 8'h2D; #100;
A = 8'hE4; B = 8'h2E; #100;
A = 8'hE4; B = 8'h2F; #100;
A = 8'hE4; B = 8'h30; #100;
A = 8'hE4; B = 8'h31; #100;
A = 8'hE4; B = 8'h32; #100;
A = 8'hE4; B = 8'h33; #100;
A = 8'hE4; B = 8'h34; #100;
A = 8'hE4; B = 8'h35; #100;
A = 8'hE4; B = 8'h36; #100;
A = 8'hE4; B = 8'h37; #100;
A = 8'hE4; B = 8'h38; #100;
A = 8'hE4; B = 8'h39; #100;
A = 8'hE4; B = 8'h3A; #100;
A = 8'hE4; B = 8'h3B; #100;
A = 8'hE4; B = 8'h3C; #100;
A = 8'hE4; B = 8'h3D; #100;
A = 8'hE4; B = 8'h3E; #100;
A = 8'hE4; B = 8'h3F; #100;
A = 8'hE4; B = 8'h40; #100;
A = 8'hE4; B = 8'h41; #100;
A = 8'hE4; B = 8'h42; #100;
A = 8'hE4; B = 8'h43; #100;
A = 8'hE4; B = 8'h44; #100;
A = 8'hE4; B = 8'h45; #100;
A = 8'hE4; B = 8'h46; #100;
A = 8'hE4; B = 8'h47; #100;
A = 8'hE4; B = 8'h48; #100;
A = 8'hE4; B = 8'h49; #100;
A = 8'hE4; B = 8'h4A; #100;
A = 8'hE4; B = 8'h4B; #100;
A = 8'hE4; B = 8'h4C; #100;
A = 8'hE4; B = 8'h4D; #100;
A = 8'hE4; B = 8'h4E; #100;
A = 8'hE4; B = 8'h4F; #100;
A = 8'hE4; B = 8'h50; #100;
A = 8'hE4; B = 8'h51; #100;
A = 8'hE4; B = 8'h52; #100;
A = 8'hE4; B = 8'h53; #100;
A = 8'hE4; B = 8'h54; #100;
A = 8'hE4; B = 8'h55; #100;
A = 8'hE4; B = 8'h56; #100;
A = 8'hE4; B = 8'h57; #100;
A = 8'hE4; B = 8'h58; #100;
A = 8'hE4; B = 8'h59; #100;
A = 8'hE4; B = 8'h5A; #100;
A = 8'hE4; B = 8'h5B; #100;
A = 8'hE4; B = 8'h5C; #100;
A = 8'hE4; B = 8'h5D; #100;
A = 8'hE4; B = 8'h5E; #100;
A = 8'hE4; B = 8'h5F; #100;
A = 8'hE4; B = 8'h60; #100;
A = 8'hE4; B = 8'h61; #100;
A = 8'hE4; B = 8'h62; #100;
A = 8'hE4; B = 8'h63; #100;
A = 8'hE4; B = 8'h64; #100;
A = 8'hE4; B = 8'h65; #100;
A = 8'hE4; B = 8'h66; #100;
A = 8'hE4; B = 8'h67; #100;
A = 8'hE4; B = 8'h68; #100;
A = 8'hE4; B = 8'h69; #100;
A = 8'hE4; B = 8'h6A; #100;
A = 8'hE4; B = 8'h6B; #100;
A = 8'hE4; B = 8'h6C; #100;
A = 8'hE4; B = 8'h6D; #100;
A = 8'hE4; B = 8'h6E; #100;
A = 8'hE4; B = 8'h6F; #100;
A = 8'hE4; B = 8'h70; #100;
A = 8'hE4; B = 8'h71; #100;
A = 8'hE4; B = 8'h72; #100;
A = 8'hE4; B = 8'h73; #100;
A = 8'hE4; B = 8'h74; #100;
A = 8'hE4; B = 8'h75; #100;
A = 8'hE4; B = 8'h76; #100;
A = 8'hE4; B = 8'h77; #100;
A = 8'hE4; B = 8'h78; #100;
A = 8'hE4; B = 8'h79; #100;
A = 8'hE4; B = 8'h7A; #100;
A = 8'hE4; B = 8'h7B; #100;
A = 8'hE4; B = 8'h7C; #100;
A = 8'hE4; B = 8'h7D; #100;
A = 8'hE4; B = 8'h7E; #100;
A = 8'hE4; B = 8'h7F; #100;
A = 8'hE4; B = 8'h80; #100;
A = 8'hE4; B = 8'h81; #100;
A = 8'hE4; B = 8'h82; #100;
A = 8'hE4; B = 8'h83; #100;
A = 8'hE4; B = 8'h84; #100;
A = 8'hE4; B = 8'h85; #100;
A = 8'hE4; B = 8'h86; #100;
A = 8'hE4; B = 8'h87; #100;
A = 8'hE4; B = 8'h88; #100;
A = 8'hE4; B = 8'h89; #100;
A = 8'hE4; B = 8'h8A; #100;
A = 8'hE4; B = 8'h8B; #100;
A = 8'hE4; B = 8'h8C; #100;
A = 8'hE4; B = 8'h8D; #100;
A = 8'hE4; B = 8'h8E; #100;
A = 8'hE4; B = 8'h8F; #100;
A = 8'hE4; B = 8'h90; #100;
A = 8'hE4; B = 8'h91; #100;
A = 8'hE4; B = 8'h92; #100;
A = 8'hE4; B = 8'h93; #100;
A = 8'hE4; B = 8'h94; #100;
A = 8'hE4; B = 8'h95; #100;
A = 8'hE4; B = 8'h96; #100;
A = 8'hE4; B = 8'h97; #100;
A = 8'hE4; B = 8'h98; #100;
A = 8'hE4; B = 8'h99; #100;
A = 8'hE4; B = 8'h9A; #100;
A = 8'hE4; B = 8'h9B; #100;
A = 8'hE4; B = 8'h9C; #100;
A = 8'hE4; B = 8'h9D; #100;
A = 8'hE4; B = 8'h9E; #100;
A = 8'hE4; B = 8'h9F; #100;
A = 8'hE4; B = 8'hA0; #100;
A = 8'hE4; B = 8'hA1; #100;
A = 8'hE4; B = 8'hA2; #100;
A = 8'hE4; B = 8'hA3; #100;
A = 8'hE4; B = 8'hA4; #100;
A = 8'hE4; B = 8'hA5; #100;
A = 8'hE4; B = 8'hA6; #100;
A = 8'hE4; B = 8'hA7; #100;
A = 8'hE4; B = 8'hA8; #100;
A = 8'hE4; B = 8'hA9; #100;
A = 8'hE4; B = 8'hAA; #100;
A = 8'hE4; B = 8'hAB; #100;
A = 8'hE4; B = 8'hAC; #100;
A = 8'hE4; B = 8'hAD; #100;
A = 8'hE4; B = 8'hAE; #100;
A = 8'hE4; B = 8'hAF; #100;
A = 8'hE4; B = 8'hB0; #100;
A = 8'hE4; B = 8'hB1; #100;
A = 8'hE4; B = 8'hB2; #100;
A = 8'hE4; B = 8'hB3; #100;
A = 8'hE4; B = 8'hB4; #100;
A = 8'hE4; B = 8'hB5; #100;
A = 8'hE4; B = 8'hB6; #100;
A = 8'hE4; B = 8'hB7; #100;
A = 8'hE4; B = 8'hB8; #100;
A = 8'hE4; B = 8'hB9; #100;
A = 8'hE4; B = 8'hBA; #100;
A = 8'hE4; B = 8'hBB; #100;
A = 8'hE4; B = 8'hBC; #100;
A = 8'hE4; B = 8'hBD; #100;
A = 8'hE4; B = 8'hBE; #100;
A = 8'hE4; B = 8'hBF; #100;
A = 8'hE4; B = 8'hC0; #100;
A = 8'hE4; B = 8'hC1; #100;
A = 8'hE4; B = 8'hC2; #100;
A = 8'hE4; B = 8'hC3; #100;
A = 8'hE4; B = 8'hC4; #100;
A = 8'hE4; B = 8'hC5; #100;
A = 8'hE4; B = 8'hC6; #100;
A = 8'hE4; B = 8'hC7; #100;
A = 8'hE4; B = 8'hC8; #100;
A = 8'hE4; B = 8'hC9; #100;
A = 8'hE4; B = 8'hCA; #100;
A = 8'hE4; B = 8'hCB; #100;
A = 8'hE4; B = 8'hCC; #100;
A = 8'hE4; B = 8'hCD; #100;
A = 8'hE4; B = 8'hCE; #100;
A = 8'hE4; B = 8'hCF; #100;
A = 8'hE4; B = 8'hD0; #100;
A = 8'hE4; B = 8'hD1; #100;
A = 8'hE4; B = 8'hD2; #100;
A = 8'hE4; B = 8'hD3; #100;
A = 8'hE4; B = 8'hD4; #100;
A = 8'hE4; B = 8'hD5; #100;
A = 8'hE4; B = 8'hD6; #100;
A = 8'hE4; B = 8'hD7; #100;
A = 8'hE4; B = 8'hD8; #100;
A = 8'hE4; B = 8'hD9; #100;
A = 8'hE4; B = 8'hDA; #100;
A = 8'hE4; B = 8'hDB; #100;
A = 8'hE4; B = 8'hDC; #100;
A = 8'hE4; B = 8'hDD; #100;
A = 8'hE4; B = 8'hDE; #100;
A = 8'hE4; B = 8'hDF; #100;
A = 8'hE4; B = 8'hE0; #100;
A = 8'hE4; B = 8'hE1; #100;
A = 8'hE4; B = 8'hE2; #100;
A = 8'hE4; B = 8'hE3; #100;
A = 8'hE4; B = 8'hE4; #100;
A = 8'hE4; B = 8'hE5; #100;
A = 8'hE4; B = 8'hE6; #100;
A = 8'hE4; B = 8'hE7; #100;
A = 8'hE4; B = 8'hE8; #100;
A = 8'hE4; B = 8'hE9; #100;
A = 8'hE4; B = 8'hEA; #100;
A = 8'hE4; B = 8'hEB; #100;
A = 8'hE4; B = 8'hEC; #100;
A = 8'hE4; B = 8'hED; #100;
A = 8'hE4; B = 8'hEE; #100;
A = 8'hE4; B = 8'hEF; #100;
A = 8'hE4; B = 8'hF0; #100;
A = 8'hE4; B = 8'hF1; #100;
A = 8'hE4; B = 8'hF2; #100;
A = 8'hE4; B = 8'hF3; #100;
A = 8'hE4; B = 8'hF4; #100;
A = 8'hE4; B = 8'hF5; #100;
A = 8'hE4; B = 8'hF6; #100;
A = 8'hE4; B = 8'hF7; #100;
A = 8'hE4; B = 8'hF8; #100;
A = 8'hE4; B = 8'hF9; #100;
A = 8'hE4; B = 8'hFA; #100;
A = 8'hE4; B = 8'hFB; #100;
A = 8'hE4; B = 8'hFC; #100;
A = 8'hE4; B = 8'hFD; #100;
A = 8'hE4; B = 8'hFE; #100;
A = 8'hE4; B = 8'hFF; #100;
A = 8'hE5; B = 8'h0; #100;
A = 8'hE5; B = 8'h1; #100;
A = 8'hE5; B = 8'h2; #100;
A = 8'hE5; B = 8'h3; #100;
A = 8'hE5; B = 8'h4; #100;
A = 8'hE5; B = 8'h5; #100;
A = 8'hE5; B = 8'h6; #100;
A = 8'hE5; B = 8'h7; #100;
A = 8'hE5; B = 8'h8; #100;
A = 8'hE5; B = 8'h9; #100;
A = 8'hE5; B = 8'hA; #100;
A = 8'hE5; B = 8'hB; #100;
A = 8'hE5; B = 8'hC; #100;
A = 8'hE5; B = 8'hD; #100;
A = 8'hE5; B = 8'hE; #100;
A = 8'hE5; B = 8'hF; #100;
A = 8'hE5; B = 8'h10; #100;
A = 8'hE5; B = 8'h11; #100;
A = 8'hE5; B = 8'h12; #100;
A = 8'hE5; B = 8'h13; #100;
A = 8'hE5; B = 8'h14; #100;
A = 8'hE5; B = 8'h15; #100;
A = 8'hE5; B = 8'h16; #100;
A = 8'hE5; B = 8'h17; #100;
A = 8'hE5; B = 8'h18; #100;
A = 8'hE5; B = 8'h19; #100;
A = 8'hE5; B = 8'h1A; #100;
A = 8'hE5; B = 8'h1B; #100;
A = 8'hE5; B = 8'h1C; #100;
A = 8'hE5; B = 8'h1D; #100;
A = 8'hE5; B = 8'h1E; #100;
A = 8'hE5; B = 8'h1F; #100;
A = 8'hE5; B = 8'h20; #100;
A = 8'hE5; B = 8'h21; #100;
A = 8'hE5; B = 8'h22; #100;
A = 8'hE5; B = 8'h23; #100;
A = 8'hE5; B = 8'h24; #100;
A = 8'hE5; B = 8'h25; #100;
A = 8'hE5; B = 8'h26; #100;
A = 8'hE5; B = 8'h27; #100;
A = 8'hE5; B = 8'h28; #100;
A = 8'hE5; B = 8'h29; #100;
A = 8'hE5; B = 8'h2A; #100;
A = 8'hE5; B = 8'h2B; #100;
A = 8'hE5; B = 8'h2C; #100;
A = 8'hE5; B = 8'h2D; #100;
A = 8'hE5; B = 8'h2E; #100;
A = 8'hE5; B = 8'h2F; #100;
A = 8'hE5; B = 8'h30; #100;
A = 8'hE5; B = 8'h31; #100;
A = 8'hE5; B = 8'h32; #100;
A = 8'hE5; B = 8'h33; #100;
A = 8'hE5; B = 8'h34; #100;
A = 8'hE5; B = 8'h35; #100;
A = 8'hE5; B = 8'h36; #100;
A = 8'hE5; B = 8'h37; #100;
A = 8'hE5; B = 8'h38; #100;
A = 8'hE5; B = 8'h39; #100;
A = 8'hE5; B = 8'h3A; #100;
A = 8'hE5; B = 8'h3B; #100;
A = 8'hE5; B = 8'h3C; #100;
A = 8'hE5; B = 8'h3D; #100;
A = 8'hE5; B = 8'h3E; #100;
A = 8'hE5; B = 8'h3F; #100;
A = 8'hE5; B = 8'h40; #100;
A = 8'hE5; B = 8'h41; #100;
A = 8'hE5; B = 8'h42; #100;
A = 8'hE5; B = 8'h43; #100;
A = 8'hE5; B = 8'h44; #100;
A = 8'hE5; B = 8'h45; #100;
A = 8'hE5; B = 8'h46; #100;
A = 8'hE5; B = 8'h47; #100;
A = 8'hE5; B = 8'h48; #100;
A = 8'hE5; B = 8'h49; #100;
A = 8'hE5; B = 8'h4A; #100;
A = 8'hE5; B = 8'h4B; #100;
A = 8'hE5; B = 8'h4C; #100;
A = 8'hE5; B = 8'h4D; #100;
A = 8'hE5; B = 8'h4E; #100;
A = 8'hE5; B = 8'h4F; #100;
A = 8'hE5; B = 8'h50; #100;
A = 8'hE5; B = 8'h51; #100;
A = 8'hE5; B = 8'h52; #100;
A = 8'hE5; B = 8'h53; #100;
A = 8'hE5; B = 8'h54; #100;
A = 8'hE5; B = 8'h55; #100;
A = 8'hE5; B = 8'h56; #100;
A = 8'hE5; B = 8'h57; #100;
A = 8'hE5; B = 8'h58; #100;
A = 8'hE5; B = 8'h59; #100;
A = 8'hE5; B = 8'h5A; #100;
A = 8'hE5; B = 8'h5B; #100;
A = 8'hE5; B = 8'h5C; #100;
A = 8'hE5; B = 8'h5D; #100;
A = 8'hE5; B = 8'h5E; #100;
A = 8'hE5; B = 8'h5F; #100;
A = 8'hE5; B = 8'h60; #100;
A = 8'hE5; B = 8'h61; #100;
A = 8'hE5; B = 8'h62; #100;
A = 8'hE5; B = 8'h63; #100;
A = 8'hE5; B = 8'h64; #100;
A = 8'hE5; B = 8'h65; #100;
A = 8'hE5; B = 8'h66; #100;
A = 8'hE5; B = 8'h67; #100;
A = 8'hE5; B = 8'h68; #100;
A = 8'hE5; B = 8'h69; #100;
A = 8'hE5; B = 8'h6A; #100;
A = 8'hE5; B = 8'h6B; #100;
A = 8'hE5; B = 8'h6C; #100;
A = 8'hE5; B = 8'h6D; #100;
A = 8'hE5; B = 8'h6E; #100;
A = 8'hE5; B = 8'h6F; #100;
A = 8'hE5; B = 8'h70; #100;
A = 8'hE5; B = 8'h71; #100;
A = 8'hE5; B = 8'h72; #100;
A = 8'hE5; B = 8'h73; #100;
A = 8'hE5; B = 8'h74; #100;
A = 8'hE5; B = 8'h75; #100;
A = 8'hE5; B = 8'h76; #100;
A = 8'hE5; B = 8'h77; #100;
A = 8'hE5; B = 8'h78; #100;
A = 8'hE5; B = 8'h79; #100;
A = 8'hE5; B = 8'h7A; #100;
A = 8'hE5; B = 8'h7B; #100;
A = 8'hE5; B = 8'h7C; #100;
A = 8'hE5; B = 8'h7D; #100;
A = 8'hE5; B = 8'h7E; #100;
A = 8'hE5; B = 8'h7F; #100;
A = 8'hE5; B = 8'h80; #100;
A = 8'hE5; B = 8'h81; #100;
A = 8'hE5; B = 8'h82; #100;
A = 8'hE5; B = 8'h83; #100;
A = 8'hE5; B = 8'h84; #100;
A = 8'hE5; B = 8'h85; #100;
A = 8'hE5; B = 8'h86; #100;
A = 8'hE5; B = 8'h87; #100;
A = 8'hE5; B = 8'h88; #100;
A = 8'hE5; B = 8'h89; #100;
A = 8'hE5; B = 8'h8A; #100;
A = 8'hE5; B = 8'h8B; #100;
A = 8'hE5; B = 8'h8C; #100;
A = 8'hE5; B = 8'h8D; #100;
A = 8'hE5; B = 8'h8E; #100;
A = 8'hE5; B = 8'h8F; #100;
A = 8'hE5; B = 8'h90; #100;
A = 8'hE5; B = 8'h91; #100;
A = 8'hE5; B = 8'h92; #100;
A = 8'hE5; B = 8'h93; #100;
A = 8'hE5; B = 8'h94; #100;
A = 8'hE5; B = 8'h95; #100;
A = 8'hE5; B = 8'h96; #100;
A = 8'hE5; B = 8'h97; #100;
A = 8'hE5; B = 8'h98; #100;
A = 8'hE5; B = 8'h99; #100;
A = 8'hE5; B = 8'h9A; #100;
A = 8'hE5; B = 8'h9B; #100;
A = 8'hE5; B = 8'h9C; #100;
A = 8'hE5; B = 8'h9D; #100;
A = 8'hE5; B = 8'h9E; #100;
A = 8'hE5; B = 8'h9F; #100;
A = 8'hE5; B = 8'hA0; #100;
A = 8'hE5; B = 8'hA1; #100;
A = 8'hE5; B = 8'hA2; #100;
A = 8'hE5; B = 8'hA3; #100;
A = 8'hE5; B = 8'hA4; #100;
A = 8'hE5; B = 8'hA5; #100;
A = 8'hE5; B = 8'hA6; #100;
A = 8'hE5; B = 8'hA7; #100;
A = 8'hE5; B = 8'hA8; #100;
A = 8'hE5; B = 8'hA9; #100;
A = 8'hE5; B = 8'hAA; #100;
A = 8'hE5; B = 8'hAB; #100;
A = 8'hE5; B = 8'hAC; #100;
A = 8'hE5; B = 8'hAD; #100;
A = 8'hE5; B = 8'hAE; #100;
A = 8'hE5; B = 8'hAF; #100;
A = 8'hE5; B = 8'hB0; #100;
A = 8'hE5; B = 8'hB1; #100;
A = 8'hE5; B = 8'hB2; #100;
A = 8'hE5; B = 8'hB3; #100;
A = 8'hE5; B = 8'hB4; #100;
A = 8'hE5; B = 8'hB5; #100;
A = 8'hE5; B = 8'hB6; #100;
A = 8'hE5; B = 8'hB7; #100;
A = 8'hE5; B = 8'hB8; #100;
A = 8'hE5; B = 8'hB9; #100;
A = 8'hE5; B = 8'hBA; #100;
A = 8'hE5; B = 8'hBB; #100;
A = 8'hE5; B = 8'hBC; #100;
A = 8'hE5; B = 8'hBD; #100;
A = 8'hE5; B = 8'hBE; #100;
A = 8'hE5; B = 8'hBF; #100;
A = 8'hE5; B = 8'hC0; #100;
A = 8'hE5; B = 8'hC1; #100;
A = 8'hE5; B = 8'hC2; #100;
A = 8'hE5; B = 8'hC3; #100;
A = 8'hE5; B = 8'hC4; #100;
A = 8'hE5; B = 8'hC5; #100;
A = 8'hE5; B = 8'hC6; #100;
A = 8'hE5; B = 8'hC7; #100;
A = 8'hE5; B = 8'hC8; #100;
A = 8'hE5; B = 8'hC9; #100;
A = 8'hE5; B = 8'hCA; #100;
A = 8'hE5; B = 8'hCB; #100;
A = 8'hE5; B = 8'hCC; #100;
A = 8'hE5; B = 8'hCD; #100;
A = 8'hE5; B = 8'hCE; #100;
A = 8'hE5; B = 8'hCF; #100;
A = 8'hE5; B = 8'hD0; #100;
A = 8'hE5; B = 8'hD1; #100;
A = 8'hE5; B = 8'hD2; #100;
A = 8'hE5; B = 8'hD3; #100;
A = 8'hE5; B = 8'hD4; #100;
A = 8'hE5; B = 8'hD5; #100;
A = 8'hE5; B = 8'hD6; #100;
A = 8'hE5; B = 8'hD7; #100;
A = 8'hE5; B = 8'hD8; #100;
A = 8'hE5; B = 8'hD9; #100;
A = 8'hE5; B = 8'hDA; #100;
A = 8'hE5; B = 8'hDB; #100;
A = 8'hE5; B = 8'hDC; #100;
A = 8'hE5; B = 8'hDD; #100;
A = 8'hE5; B = 8'hDE; #100;
A = 8'hE5; B = 8'hDF; #100;
A = 8'hE5; B = 8'hE0; #100;
A = 8'hE5; B = 8'hE1; #100;
A = 8'hE5; B = 8'hE2; #100;
A = 8'hE5; B = 8'hE3; #100;
A = 8'hE5; B = 8'hE4; #100;
A = 8'hE5; B = 8'hE5; #100;
A = 8'hE5; B = 8'hE6; #100;
A = 8'hE5; B = 8'hE7; #100;
A = 8'hE5; B = 8'hE8; #100;
A = 8'hE5; B = 8'hE9; #100;
A = 8'hE5; B = 8'hEA; #100;
A = 8'hE5; B = 8'hEB; #100;
A = 8'hE5; B = 8'hEC; #100;
A = 8'hE5; B = 8'hED; #100;
A = 8'hE5; B = 8'hEE; #100;
A = 8'hE5; B = 8'hEF; #100;
A = 8'hE5; B = 8'hF0; #100;
A = 8'hE5; B = 8'hF1; #100;
A = 8'hE5; B = 8'hF2; #100;
A = 8'hE5; B = 8'hF3; #100;
A = 8'hE5; B = 8'hF4; #100;
A = 8'hE5; B = 8'hF5; #100;
A = 8'hE5; B = 8'hF6; #100;
A = 8'hE5; B = 8'hF7; #100;
A = 8'hE5; B = 8'hF8; #100;
A = 8'hE5; B = 8'hF9; #100;
A = 8'hE5; B = 8'hFA; #100;
A = 8'hE5; B = 8'hFB; #100;
A = 8'hE5; B = 8'hFC; #100;
A = 8'hE5; B = 8'hFD; #100;
A = 8'hE5; B = 8'hFE; #100;
A = 8'hE5; B = 8'hFF; #100;
A = 8'hE6; B = 8'h0; #100;
A = 8'hE6; B = 8'h1; #100;
A = 8'hE6; B = 8'h2; #100;
A = 8'hE6; B = 8'h3; #100;
A = 8'hE6; B = 8'h4; #100;
A = 8'hE6; B = 8'h5; #100;
A = 8'hE6; B = 8'h6; #100;
A = 8'hE6; B = 8'h7; #100;
A = 8'hE6; B = 8'h8; #100;
A = 8'hE6; B = 8'h9; #100;
A = 8'hE6; B = 8'hA; #100;
A = 8'hE6; B = 8'hB; #100;
A = 8'hE6; B = 8'hC; #100;
A = 8'hE6; B = 8'hD; #100;
A = 8'hE6; B = 8'hE; #100;
A = 8'hE6; B = 8'hF; #100;
A = 8'hE6; B = 8'h10; #100;
A = 8'hE6; B = 8'h11; #100;
A = 8'hE6; B = 8'h12; #100;
A = 8'hE6; B = 8'h13; #100;
A = 8'hE6; B = 8'h14; #100;
A = 8'hE6; B = 8'h15; #100;
A = 8'hE6; B = 8'h16; #100;
A = 8'hE6; B = 8'h17; #100;
A = 8'hE6; B = 8'h18; #100;
A = 8'hE6; B = 8'h19; #100;
A = 8'hE6; B = 8'h1A; #100;
A = 8'hE6; B = 8'h1B; #100;
A = 8'hE6; B = 8'h1C; #100;
A = 8'hE6; B = 8'h1D; #100;
A = 8'hE6; B = 8'h1E; #100;
A = 8'hE6; B = 8'h1F; #100;
A = 8'hE6; B = 8'h20; #100;
A = 8'hE6; B = 8'h21; #100;
A = 8'hE6; B = 8'h22; #100;
A = 8'hE6; B = 8'h23; #100;
A = 8'hE6; B = 8'h24; #100;
A = 8'hE6; B = 8'h25; #100;
A = 8'hE6; B = 8'h26; #100;
A = 8'hE6; B = 8'h27; #100;
A = 8'hE6; B = 8'h28; #100;
A = 8'hE6; B = 8'h29; #100;
A = 8'hE6; B = 8'h2A; #100;
A = 8'hE6; B = 8'h2B; #100;
A = 8'hE6; B = 8'h2C; #100;
A = 8'hE6; B = 8'h2D; #100;
A = 8'hE6; B = 8'h2E; #100;
A = 8'hE6; B = 8'h2F; #100;
A = 8'hE6; B = 8'h30; #100;
A = 8'hE6; B = 8'h31; #100;
A = 8'hE6; B = 8'h32; #100;
A = 8'hE6; B = 8'h33; #100;
A = 8'hE6; B = 8'h34; #100;
A = 8'hE6; B = 8'h35; #100;
A = 8'hE6; B = 8'h36; #100;
A = 8'hE6; B = 8'h37; #100;
A = 8'hE6; B = 8'h38; #100;
A = 8'hE6; B = 8'h39; #100;
A = 8'hE6; B = 8'h3A; #100;
A = 8'hE6; B = 8'h3B; #100;
A = 8'hE6; B = 8'h3C; #100;
A = 8'hE6; B = 8'h3D; #100;
A = 8'hE6; B = 8'h3E; #100;
A = 8'hE6; B = 8'h3F; #100;
A = 8'hE6; B = 8'h40; #100;
A = 8'hE6; B = 8'h41; #100;
A = 8'hE6; B = 8'h42; #100;
A = 8'hE6; B = 8'h43; #100;
A = 8'hE6; B = 8'h44; #100;
A = 8'hE6; B = 8'h45; #100;
A = 8'hE6; B = 8'h46; #100;
A = 8'hE6; B = 8'h47; #100;
A = 8'hE6; B = 8'h48; #100;
A = 8'hE6; B = 8'h49; #100;
A = 8'hE6; B = 8'h4A; #100;
A = 8'hE6; B = 8'h4B; #100;
A = 8'hE6; B = 8'h4C; #100;
A = 8'hE6; B = 8'h4D; #100;
A = 8'hE6; B = 8'h4E; #100;
A = 8'hE6; B = 8'h4F; #100;
A = 8'hE6; B = 8'h50; #100;
A = 8'hE6; B = 8'h51; #100;
A = 8'hE6; B = 8'h52; #100;
A = 8'hE6; B = 8'h53; #100;
A = 8'hE6; B = 8'h54; #100;
A = 8'hE6; B = 8'h55; #100;
A = 8'hE6; B = 8'h56; #100;
A = 8'hE6; B = 8'h57; #100;
A = 8'hE6; B = 8'h58; #100;
A = 8'hE6; B = 8'h59; #100;
A = 8'hE6; B = 8'h5A; #100;
A = 8'hE6; B = 8'h5B; #100;
A = 8'hE6; B = 8'h5C; #100;
A = 8'hE6; B = 8'h5D; #100;
A = 8'hE6; B = 8'h5E; #100;
A = 8'hE6; B = 8'h5F; #100;
A = 8'hE6; B = 8'h60; #100;
A = 8'hE6; B = 8'h61; #100;
A = 8'hE6; B = 8'h62; #100;
A = 8'hE6; B = 8'h63; #100;
A = 8'hE6; B = 8'h64; #100;
A = 8'hE6; B = 8'h65; #100;
A = 8'hE6; B = 8'h66; #100;
A = 8'hE6; B = 8'h67; #100;
A = 8'hE6; B = 8'h68; #100;
A = 8'hE6; B = 8'h69; #100;
A = 8'hE6; B = 8'h6A; #100;
A = 8'hE6; B = 8'h6B; #100;
A = 8'hE6; B = 8'h6C; #100;
A = 8'hE6; B = 8'h6D; #100;
A = 8'hE6; B = 8'h6E; #100;
A = 8'hE6; B = 8'h6F; #100;
A = 8'hE6; B = 8'h70; #100;
A = 8'hE6; B = 8'h71; #100;
A = 8'hE6; B = 8'h72; #100;
A = 8'hE6; B = 8'h73; #100;
A = 8'hE6; B = 8'h74; #100;
A = 8'hE6; B = 8'h75; #100;
A = 8'hE6; B = 8'h76; #100;
A = 8'hE6; B = 8'h77; #100;
A = 8'hE6; B = 8'h78; #100;
A = 8'hE6; B = 8'h79; #100;
A = 8'hE6; B = 8'h7A; #100;
A = 8'hE6; B = 8'h7B; #100;
A = 8'hE6; B = 8'h7C; #100;
A = 8'hE6; B = 8'h7D; #100;
A = 8'hE6; B = 8'h7E; #100;
A = 8'hE6; B = 8'h7F; #100;
A = 8'hE6; B = 8'h80; #100;
A = 8'hE6; B = 8'h81; #100;
A = 8'hE6; B = 8'h82; #100;
A = 8'hE6; B = 8'h83; #100;
A = 8'hE6; B = 8'h84; #100;
A = 8'hE6; B = 8'h85; #100;
A = 8'hE6; B = 8'h86; #100;
A = 8'hE6; B = 8'h87; #100;
A = 8'hE6; B = 8'h88; #100;
A = 8'hE6; B = 8'h89; #100;
A = 8'hE6; B = 8'h8A; #100;
A = 8'hE6; B = 8'h8B; #100;
A = 8'hE6; B = 8'h8C; #100;
A = 8'hE6; B = 8'h8D; #100;
A = 8'hE6; B = 8'h8E; #100;
A = 8'hE6; B = 8'h8F; #100;
A = 8'hE6; B = 8'h90; #100;
A = 8'hE6; B = 8'h91; #100;
A = 8'hE6; B = 8'h92; #100;
A = 8'hE6; B = 8'h93; #100;
A = 8'hE6; B = 8'h94; #100;
A = 8'hE6; B = 8'h95; #100;
A = 8'hE6; B = 8'h96; #100;
A = 8'hE6; B = 8'h97; #100;
A = 8'hE6; B = 8'h98; #100;
A = 8'hE6; B = 8'h99; #100;
A = 8'hE6; B = 8'h9A; #100;
A = 8'hE6; B = 8'h9B; #100;
A = 8'hE6; B = 8'h9C; #100;
A = 8'hE6; B = 8'h9D; #100;
A = 8'hE6; B = 8'h9E; #100;
A = 8'hE6; B = 8'h9F; #100;
A = 8'hE6; B = 8'hA0; #100;
A = 8'hE6; B = 8'hA1; #100;
A = 8'hE6; B = 8'hA2; #100;
A = 8'hE6; B = 8'hA3; #100;
A = 8'hE6; B = 8'hA4; #100;
A = 8'hE6; B = 8'hA5; #100;
A = 8'hE6; B = 8'hA6; #100;
A = 8'hE6; B = 8'hA7; #100;
A = 8'hE6; B = 8'hA8; #100;
A = 8'hE6; B = 8'hA9; #100;
A = 8'hE6; B = 8'hAA; #100;
A = 8'hE6; B = 8'hAB; #100;
A = 8'hE6; B = 8'hAC; #100;
A = 8'hE6; B = 8'hAD; #100;
A = 8'hE6; B = 8'hAE; #100;
A = 8'hE6; B = 8'hAF; #100;
A = 8'hE6; B = 8'hB0; #100;
A = 8'hE6; B = 8'hB1; #100;
A = 8'hE6; B = 8'hB2; #100;
A = 8'hE6; B = 8'hB3; #100;
A = 8'hE6; B = 8'hB4; #100;
A = 8'hE6; B = 8'hB5; #100;
A = 8'hE6; B = 8'hB6; #100;
A = 8'hE6; B = 8'hB7; #100;
A = 8'hE6; B = 8'hB8; #100;
A = 8'hE6; B = 8'hB9; #100;
A = 8'hE6; B = 8'hBA; #100;
A = 8'hE6; B = 8'hBB; #100;
A = 8'hE6; B = 8'hBC; #100;
A = 8'hE6; B = 8'hBD; #100;
A = 8'hE6; B = 8'hBE; #100;
A = 8'hE6; B = 8'hBF; #100;
A = 8'hE6; B = 8'hC0; #100;
A = 8'hE6; B = 8'hC1; #100;
A = 8'hE6; B = 8'hC2; #100;
A = 8'hE6; B = 8'hC3; #100;
A = 8'hE6; B = 8'hC4; #100;
A = 8'hE6; B = 8'hC5; #100;
A = 8'hE6; B = 8'hC6; #100;
A = 8'hE6; B = 8'hC7; #100;
A = 8'hE6; B = 8'hC8; #100;
A = 8'hE6; B = 8'hC9; #100;
A = 8'hE6; B = 8'hCA; #100;
A = 8'hE6; B = 8'hCB; #100;
A = 8'hE6; B = 8'hCC; #100;
A = 8'hE6; B = 8'hCD; #100;
A = 8'hE6; B = 8'hCE; #100;
A = 8'hE6; B = 8'hCF; #100;
A = 8'hE6; B = 8'hD0; #100;
A = 8'hE6; B = 8'hD1; #100;
A = 8'hE6; B = 8'hD2; #100;
A = 8'hE6; B = 8'hD3; #100;
A = 8'hE6; B = 8'hD4; #100;
A = 8'hE6; B = 8'hD5; #100;
A = 8'hE6; B = 8'hD6; #100;
A = 8'hE6; B = 8'hD7; #100;
A = 8'hE6; B = 8'hD8; #100;
A = 8'hE6; B = 8'hD9; #100;
A = 8'hE6; B = 8'hDA; #100;
A = 8'hE6; B = 8'hDB; #100;
A = 8'hE6; B = 8'hDC; #100;
A = 8'hE6; B = 8'hDD; #100;
A = 8'hE6; B = 8'hDE; #100;
A = 8'hE6; B = 8'hDF; #100;
A = 8'hE6; B = 8'hE0; #100;
A = 8'hE6; B = 8'hE1; #100;
A = 8'hE6; B = 8'hE2; #100;
A = 8'hE6; B = 8'hE3; #100;
A = 8'hE6; B = 8'hE4; #100;
A = 8'hE6; B = 8'hE5; #100;
A = 8'hE6; B = 8'hE6; #100;
A = 8'hE6; B = 8'hE7; #100;
A = 8'hE6; B = 8'hE8; #100;
A = 8'hE6; B = 8'hE9; #100;
A = 8'hE6; B = 8'hEA; #100;
A = 8'hE6; B = 8'hEB; #100;
A = 8'hE6; B = 8'hEC; #100;
A = 8'hE6; B = 8'hED; #100;
A = 8'hE6; B = 8'hEE; #100;
A = 8'hE6; B = 8'hEF; #100;
A = 8'hE6; B = 8'hF0; #100;
A = 8'hE6; B = 8'hF1; #100;
A = 8'hE6; B = 8'hF2; #100;
A = 8'hE6; B = 8'hF3; #100;
A = 8'hE6; B = 8'hF4; #100;
A = 8'hE6; B = 8'hF5; #100;
A = 8'hE6; B = 8'hF6; #100;
A = 8'hE6; B = 8'hF7; #100;
A = 8'hE6; B = 8'hF8; #100;
A = 8'hE6; B = 8'hF9; #100;
A = 8'hE6; B = 8'hFA; #100;
A = 8'hE6; B = 8'hFB; #100;
A = 8'hE6; B = 8'hFC; #100;
A = 8'hE6; B = 8'hFD; #100;
A = 8'hE6; B = 8'hFE; #100;
A = 8'hE6; B = 8'hFF; #100;
A = 8'hE7; B = 8'h0; #100;
A = 8'hE7; B = 8'h1; #100;
A = 8'hE7; B = 8'h2; #100;
A = 8'hE7; B = 8'h3; #100;
A = 8'hE7; B = 8'h4; #100;
A = 8'hE7; B = 8'h5; #100;
A = 8'hE7; B = 8'h6; #100;
A = 8'hE7; B = 8'h7; #100;
A = 8'hE7; B = 8'h8; #100;
A = 8'hE7; B = 8'h9; #100;
A = 8'hE7; B = 8'hA; #100;
A = 8'hE7; B = 8'hB; #100;
A = 8'hE7; B = 8'hC; #100;
A = 8'hE7; B = 8'hD; #100;
A = 8'hE7; B = 8'hE; #100;
A = 8'hE7; B = 8'hF; #100;
A = 8'hE7; B = 8'h10; #100;
A = 8'hE7; B = 8'h11; #100;
A = 8'hE7; B = 8'h12; #100;
A = 8'hE7; B = 8'h13; #100;
A = 8'hE7; B = 8'h14; #100;
A = 8'hE7; B = 8'h15; #100;
A = 8'hE7; B = 8'h16; #100;
A = 8'hE7; B = 8'h17; #100;
A = 8'hE7; B = 8'h18; #100;
A = 8'hE7; B = 8'h19; #100;
A = 8'hE7; B = 8'h1A; #100;
A = 8'hE7; B = 8'h1B; #100;
A = 8'hE7; B = 8'h1C; #100;
A = 8'hE7; B = 8'h1D; #100;
A = 8'hE7; B = 8'h1E; #100;
A = 8'hE7; B = 8'h1F; #100;
A = 8'hE7; B = 8'h20; #100;
A = 8'hE7; B = 8'h21; #100;
A = 8'hE7; B = 8'h22; #100;
A = 8'hE7; B = 8'h23; #100;
A = 8'hE7; B = 8'h24; #100;
A = 8'hE7; B = 8'h25; #100;
A = 8'hE7; B = 8'h26; #100;
A = 8'hE7; B = 8'h27; #100;
A = 8'hE7; B = 8'h28; #100;
A = 8'hE7; B = 8'h29; #100;
A = 8'hE7; B = 8'h2A; #100;
A = 8'hE7; B = 8'h2B; #100;
A = 8'hE7; B = 8'h2C; #100;
A = 8'hE7; B = 8'h2D; #100;
A = 8'hE7; B = 8'h2E; #100;
A = 8'hE7; B = 8'h2F; #100;
A = 8'hE7; B = 8'h30; #100;
A = 8'hE7; B = 8'h31; #100;
A = 8'hE7; B = 8'h32; #100;
A = 8'hE7; B = 8'h33; #100;
A = 8'hE7; B = 8'h34; #100;
A = 8'hE7; B = 8'h35; #100;
A = 8'hE7; B = 8'h36; #100;
A = 8'hE7; B = 8'h37; #100;
A = 8'hE7; B = 8'h38; #100;
A = 8'hE7; B = 8'h39; #100;
A = 8'hE7; B = 8'h3A; #100;
A = 8'hE7; B = 8'h3B; #100;
A = 8'hE7; B = 8'h3C; #100;
A = 8'hE7; B = 8'h3D; #100;
A = 8'hE7; B = 8'h3E; #100;
A = 8'hE7; B = 8'h3F; #100;
A = 8'hE7; B = 8'h40; #100;
A = 8'hE7; B = 8'h41; #100;
A = 8'hE7; B = 8'h42; #100;
A = 8'hE7; B = 8'h43; #100;
A = 8'hE7; B = 8'h44; #100;
A = 8'hE7; B = 8'h45; #100;
A = 8'hE7; B = 8'h46; #100;
A = 8'hE7; B = 8'h47; #100;
A = 8'hE7; B = 8'h48; #100;
A = 8'hE7; B = 8'h49; #100;
A = 8'hE7; B = 8'h4A; #100;
A = 8'hE7; B = 8'h4B; #100;
A = 8'hE7; B = 8'h4C; #100;
A = 8'hE7; B = 8'h4D; #100;
A = 8'hE7; B = 8'h4E; #100;
A = 8'hE7; B = 8'h4F; #100;
A = 8'hE7; B = 8'h50; #100;
A = 8'hE7; B = 8'h51; #100;
A = 8'hE7; B = 8'h52; #100;
A = 8'hE7; B = 8'h53; #100;
A = 8'hE7; B = 8'h54; #100;
A = 8'hE7; B = 8'h55; #100;
A = 8'hE7; B = 8'h56; #100;
A = 8'hE7; B = 8'h57; #100;
A = 8'hE7; B = 8'h58; #100;
A = 8'hE7; B = 8'h59; #100;
A = 8'hE7; B = 8'h5A; #100;
A = 8'hE7; B = 8'h5B; #100;
A = 8'hE7; B = 8'h5C; #100;
A = 8'hE7; B = 8'h5D; #100;
A = 8'hE7; B = 8'h5E; #100;
A = 8'hE7; B = 8'h5F; #100;
A = 8'hE7; B = 8'h60; #100;
A = 8'hE7; B = 8'h61; #100;
A = 8'hE7; B = 8'h62; #100;
A = 8'hE7; B = 8'h63; #100;
A = 8'hE7; B = 8'h64; #100;
A = 8'hE7; B = 8'h65; #100;
A = 8'hE7; B = 8'h66; #100;
A = 8'hE7; B = 8'h67; #100;
A = 8'hE7; B = 8'h68; #100;
A = 8'hE7; B = 8'h69; #100;
A = 8'hE7; B = 8'h6A; #100;
A = 8'hE7; B = 8'h6B; #100;
A = 8'hE7; B = 8'h6C; #100;
A = 8'hE7; B = 8'h6D; #100;
A = 8'hE7; B = 8'h6E; #100;
A = 8'hE7; B = 8'h6F; #100;
A = 8'hE7; B = 8'h70; #100;
A = 8'hE7; B = 8'h71; #100;
A = 8'hE7; B = 8'h72; #100;
A = 8'hE7; B = 8'h73; #100;
A = 8'hE7; B = 8'h74; #100;
A = 8'hE7; B = 8'h75; #100;
A = 8'hE7; B = 8'h76; #100;
A = 8'hE7; B = 8'h77; #100;
A = 8'hE7; B = 8'h78; #100;
A = 8'hE7; B = 8'h79; #100;
A = 8'hE7; B = 8'h7A; #100;
A = 8'hE7; B = 8'h7B; #100;
A = 8'hE7; B = 8'h7C; #100;
A = 8'hE7; B = 8'h7D; #100;
A = 8'hE7; B = 8'h7E; #100;
A = 8'hE7; B = 8'h7F; #100;
A = 8'hE7; B = 8'h80; #100;
A = 8'hE7; B = 8'h81; #100;
A = 8'hE7; B = 8'h82; #100;
A = 8'hE7; B = 8'h83; #100;
A = 8'hE7; B = 8'h84; #100;
A = 8'hE7; B = 8'h85; #100;
A = 8'hE7; B = 8'h86; #100;
A = 8'hE7; B = 8'h87; #100;
A = 8'hE7; B = 8'h88; #100;
A = 8'hE7; B = 8'h89; #100;
A = 8'hE7; B = 8'h8A; #100;
A = 8'hE7; B = 8'h8B; #100;
A = 8'hE7; B = 8'h8C; #100;
A = 8'hE7; B = 8'h8D; #100;
A = 8'hE7; B = 8'h8E; #100;
A = 8'hE7; B = 8'h8F; #100;
A = 8'hE7; B = 8'h90; #100;
A = 8'hE7; B = 8'h91; #100;
A = 8'hE7; B = 8'h92; #100;
A = 8'hE7; B = 8'h93; #100;
A = 8'hE7; B = 8'h94; #100;
A = 8'hE7; B = 8'h95; #100;
A = 8'hE7; B = 8'h96; #100;
A = 8'hE7; B = 8'h97; #100;
A = 8'hE7; B = 8'h98; #100;
A = 8'hE7; B = 8'h99; #100;
A = 8'hE7; B = 8'h9A; #100;
A = 8'hE7; B = 8'h9B; #100;
A = 8'hE7; B = 8'h9C; #100;
A = 8'hE7; B = 8'h9D; #100;
A = 8'hE7; B = 8'h9E; #100;
A = 8'hE7; B = 8'h9F; #100;
A = 8'hE7; B = 8'hA0; #100;
A = 8'hE7; B = 8'hA1; #100;
A = 8'hE7; B = 8'hA2; #100;
A = 8'hE7; B = 8'hA3; #100;
A = 8'hE7; B = 8'hA4; #100;
A = 8'hE7; B = 8'hA5; #100;
A = 8'hE7; B = 8'hA6; #100;
A = 8'hE7; B = 8'hA7; #100;
A = 8'hE7; B = 8'hA8; #100;
A = 8'hE7; B = 8'hA9; #100;
A = 8'hE7; B = 8'hAA; #100;
A = 8'hE7; B = 8'hAB; #100;
A = 8'hE7; B = 8'hAC; #100;
A = 8'hE7; B = 8'hAD; #100;
A = 8'hE7; B = 8'hAE; #100;
A = 8'hE7; B = 8'hAF; #100;
A = 8'hE7; B = 8'hB0; #100;
A = 8'hE7; B = 8'hB1; #100;
A = 8'hE7; B = 8'hB2; #100;
A = 8'hE7; B = 8'hB3; #100;
A = 8'hE7; B = 8'hB4; #100;
A = 8'hE7; B = 8'hB5; #100;
A = 8'hE7; B = 8'hB6; #100;
A = 8'hE7; B = 8'hB7; #100;
A = 8'hE7; B = 8'hB8; #100;
A = 8'hE7; B = 8'hB9; #100;
A = 8'hE7; B = 8'hBA; #100;
A = 8'hE7; B = 8'hBB; #100;
A = 8'hE7; B = 8'hBC; #100;
A = 8'hE7; B = 8'hBD; #100;
A = 8'hE7; B = 8'hBE; #100;
A = 8'hE7; B = 8'hBF; #100;
A = 8'hE7; B = 8'hC0; #100;
A = 8'hE7; B = 8'hC1; #100;
A = 8'hE7; B = 8'hC2; #100;
A = 8'hE7; B = 8'hC3; #100;
A = 8'hE7; B = 8'hC4; #100;
A = 8'hE7; B = 8'hC5; #100;
A = 8'hE7; B = 8'hC6; #100;
A = 8'hE7; B = 8'hC7; #100;
A = 8'hE7; B = 8'hC8; #100;
A = 8'hE7; B = 8'hC9; #100;
A = 8'hE7; B = 8'hCA; #100;
A = 8'hE7; B = 8'hCB; #100;
A = 8'hE7; B = 8'hCC; #100;
A = 8'hE7; B = 8'hCD; #100;
A = 8'hE7; B = 8'hCE; #100;
A = 8'hE7; B = 8'hCF; #100;
A = 8'hE7; B = 8'hD0; #100;
A = 8'hE7; B = 8'hD1; #100;
A = 8'hE7; B = 8'hD2; #100;
A = 8'hE7; B = 8'hD3; #100;
A = 8'hE7; B = 8'hD4; #100;
A = 8'hE7; B = 8'hD5; #100;
A = 8'hE7; B = 8'hD6; #100;
A = 8'hE7; B = 8'hD7; #100;
A = 8'hE7; B = 8'hD8; #100;
A = 8'hE7; B = 8'hD9; #100;
A = 8'hE7; B = 8'hDA; #100;
A = 8'hE7; B = 8'hDB; #100;
A = 8'hE7; B = 8'hDC; #100;
A = 8'hE7; B = 8'hDD; #100;
A = 8'hE7; B = 8'hDE; #100;
A = 8'hE7; B = 8'hDF; #100;
A = 8'hE7; B = 8'hE0; #100;
A = 8'hE7; B = 8'hE1; #100;
A = 8'hE7; B = 8'hE2; #100;
A = 8'hE7; B = 8'hE3; #100;
A = 8'hE7; B = 8'hE4; #100;
A = 8'hE7; B = 8'hE5; #100;
A = 8'hE7; B = 8'hE6; #100;
A = 8'hE7; B = 8'hE7; #100;
A = 8'hE7; B = 8'hE8; #100;
A = 8'hE7; B = 8'hE9; #100;
A = 8'hE7; B = 8'hEA; #100;
A = 8'hE7; B = 8'hEB; #100;
A = 8'hE7; B = 8'hEC; #100;
A = 8'hE7; B = 8'hED; #100;
A = 8'hE7; B = 8'hEE; #100;
A = 8'hE7; B = 8'hEF; #100;
A = 8'hE7; B = 8'hF0; #100;
A = 8'hE7; B = 8'hF1; #100;
A = 8'hE7; B = 8'hF2; #100;
A = 8'hE7; B = 8'hF3; #100;
A = 8'hE7; B = 8'hF4; #100;
A = 8'hE7; B = 8'hF5; #100;
A = 8'hE7; B = 8'hF6; #100;
A = 8'hE7; B = 8'hF7; #100;
A = 8'hE7; B = 8'hF8; #100;
A = 8'hE7; B = 8'hF9; #100;
A = 8'hE7; B = 8'hFA; #100;
A = 8'hE7; B = 8'hFB; #100;
A = 8'hE7; B = 8'hFC; #100;
A = 8'hE7; B = 8'hFD; #100;
A = 8'hE7; B = 8'hFE; #100;
A = 8'hE7; B = 8'hFF; #100;
A = 8'hE8; B = 8'h0; #100;
A = 8'hE8; B = 8'h1; #100;
A = 8'hE8; B = 8'h2; #100;
A = 8'hE8; B = 8'h3; #100;
A = 8'hE8; B = 8'h4; #100;
A = 8'hE8; B = 8'h5; #100;
A = 8'hE8; B = 8'h6; #100;
A = 8'hE8; B = 8'h7; #100;
A = 8'hE8; B = 8'h8; #100;
A = 8'hE8; B = 8'h9; #100;
A = 8'hE8; B = 8'hA; #100;
A = 8'hE8; B = 8'hB; #100;
A = 8'hE8; B = 8'hC; #100;
A = 8'hE8; B = 8'hD; #100;
A = 8'hE8; B = 8'hE; #100;
A = 8'hE8; B = 8'hF; #100;
A = 8'hE8; B = 8'h10; #100;
A = 8'hE8; B = 8'h11; #100;
A = 8'hE8; B = 8'h12; #100;
A = 8'hE8; B = 8'h13; #100;
A = 8'hE8; B = 8'h14; #100;
A = 8'hE8; B = 8'h15; #100;
A = 8'hE8; B = 8'h16; #100;
A = 8'hE8; B = 8'h17; #100;
A = 8'hE8; B = 8'h18; #100;
A = 8'hE8; B = 8'h19; #100;
A = 8'hE8; B = 8'h1A; #100;
A = 8'hE8; B = 8'h1B; #100;
A = 8'hE8; B = 8'h1C; #100;
A = 8'hE8; B = 8'h1D; #100;
A = 8'hE8; B = 8'h1E; #100;
A = 8'hE8; B = 8'h1F; #100;
A = 8'hE8; B = 8'h20; #100;
A = 8'hE8; B = 8'h21; #100;
A = 8'hE8; B = 8'h22; #100;
A = 8'hE8; B = 8'h23; #100;
A = 8'hE8; B = 8'h24; #100;
A = 8'hE8; B = 8'h25; #100;
A = 8'hE8; B = 8'h26; #100;
A = 8'hE8; B = 8'h27; #100;
A = 8'hE8; B = 8'h28; #100;
A = 8'hE8; B = 8'h29; #100;
A = 8'hE8; B = 8'h2A; #100;
A = 8'hE8; B = 8'h2B; #100;
A = 8'hE8; B = 8'h2C; #100;
A = 8'hE8; B = 8'h2D; #100;
A = 8'hE8; B = 8'h2E; #100;
A = 8'hE8; B = 8'h2F; #100;
A = 8'hE8; B = 8'h30; #100;
A = 8'hE8; B = 8'h31; #100;
A = 8'hE8; B = 8'h32; #100;
A = 8'hE8; B = 8'h33; #100;
A = 8'hE8; B = 8'h34; #100;
A = 8'hE8; B = 8'h35; #100;
A = 8'hE8; B = 8'h36; #100;
A = 8'hE8; B = 8'h37; #100;
A = 8'hE8; B = 8'h38; #100;
A = 8'hE8; B = 8'h39; #100;
A = 8'hE8; B = 8'h3A; #100;
A = 8'hE8; B = 8'h3B; #100;
A = 8'hE8; B = 8'h3C; #100;
A = 8'hE8; B = 8'h3D; #100;
A = 8'hE8; B = 8'h3E; #100;
A = 8'hE8; B = 8'h3F; #100;
A = 8'hE8; B = 8'h40; #100;
A = 8'hE8; B = 8'h41; #100;
A = 8'hE8; B = 8'h42; #100;
A = 8'hE8; B = 8'h43; #100;
A = 8'hE8; B = 8'h44; #100;
A = 8'hE8; B = 8'h45; #100;
A = 8'hE8; B = 8'h46; #100;
A = 8'hE8; B = 8'h47; #100;
A = 8'hE8; B = 8'h48; #100;
A = 8'hE8; B = 8'h49; #100;
A = 8'hE8; B = 8'h4A; #100;
A = 8'hE8; B = 8'h4B; #100;
A = 8'hE8; B = 8'h4C; #100;
A = 8'hE8; B = 8'h4D; #100;
A = 8'hE8; B = 8'h4E; #100;
A = 8'hE8; B = 8'h4F; #100;
A = 8'hE8; B = 8'h50; #100;
A = 8'hE8; B = 8'h51; #100;
A = 8'hE8; B = 8'h52; #100;
A = 8'hE8; B = 8'h53; #100;
A = 8'hE8; B = 8'h54; #100;
A = 8'hE8; B = 8'h55; #100;
A = 8'hE8; B = 8'h56; #100;
A = 8'hE8; B = 8'h57; #100;
A = 8'hE8; B = 8'h58; #100;
A = 8'hE8; B = 8'h59; #100;
A = 8'hE8; B = 8'h5A; #100;
A = 8'hE8; B = 8'h5B; #100;
A = 8'hE8; B = 8'h5C; #100;
A = 8'hE8; B = 8'h5D; #100;
A = 8'hE8; B = 8'h5E; #100;
A = 8'hE8; B = 8'h5F; #100;
A = 8'hE8; B = 8'h60; #100;
A = 8'hE8; B = 8'h61; #100;
A = 8'hE8; B = 8'h62; #100;
A = 8'hE8; B = 8'h63; #100;
A = 8'hE8; B = 8'h64; #100;
A = 8'hE8; B = 8'h65; #100;
A = 8'hE8; B = 8'h66; #100;
A = 8'hE8; B = 8'h67; #100;
A = 8'hE8; B = 8'h68; #100;
A = 8'hE8; B = 8'h69; #100;
A = 8'hE8; B = 8'h6A; #100;
A = 8'hE8; B = 8'h6B; #100;
A = 8'hE8; B = 8'h6C; #100;
A = 8'hE8; B = 8'h6D; #100;
A = 8'hE8; B = 8'h6E; #100;
A = 8'hE8; B = 8'h6F; #100;
A = 8'hE8; B = 8'h70; #100;
A = 8'hE8; B = 8'h71; #100;
A = 8'hE8; B = 8'h72; #100;
A = 8'hE8; B = 8'h73; #100;
A = 8'hE8; B = 8'h74; #100;
A = 8'hE8; B = 8'h75; #100;
A = 8'hE8; B = 8'h76; #100;
A = 8'hE8; B = 8'h77; #100;
A = 8'hE8; B = 8'h78; #100;
A = 8'hE8; B = 8'h79; #100;
A = 8'hE8; B = 8'h7A; #100;
A = 8'hE8; B = 8'h7B; #100;
A = 8'hE8; B = 8'h7C; #100;
A = 8'hE8; B = 8'h7D; #100;
A = 8'hE8; B = 8'h7E; #100;
A = 8'hE8; B = 8'h7F; #100;
A = 8'hE8; B = 8'h80; #100;
A = 8'hE8; B = 8'h81; #100;
A = 8'hE8; B = 8'h82; #100;
A = 8'hE8; B = 8'h83; #100;
A = 8'hE8; B = 8'h84; #100;
A = 8'hE8; B = 8'h85; #100;
A = 8'hE8; B = 8'h86; #100;
A = 8'hE8; B = 8'h87; #100;
A = 8'hE8; B = 8'h88; #100;
A = 8'hE8; B = 8'h89; #100;
A = 8'hE8; B = 8'h8A; #100;
A = 8'hE8; B = 8'h8B; #100;
A = 8'hE8; B = 8'h8C; #100;
A = 8'hE8; B = 8'h8D; #100;
A = 8'hE8; B = 8'h8E; #100;
A = 8'hE8; B = 8'h8F; #100;
A = 8'hE8; B = 8'h90; #100;
A = 8'hE8; B = 8'h91; #100;
A = 8'hE8; B = 8'h92; #100;
A = 8'hE8; B = 8'h93; #100;
A = 8'hE8; B = 8'h94; #100;
A = 8'hE8; B = 8'h95; #100;
A = 8'hE8; B = 8'h96; #100;
A = 8'hE8; B = 8'h97; #100;
A = 8'hE8; B = 8'h98; #100;
A = 8'hE8; B = 8'h99; #100;
A = 8'hE8; B = 8'h9A; #100;
A = 8'hE8; B = 8'h9B; #100;
A = 8'hE8; B = 8'h9C; #100;
A = 8'hE8; B = 8'h9D; #100;
A = 8'hE8; B = 8'h9E; #100;
A = 8'hE8; B = 8'h9F; #100;
A = 8'hE8; B = 8'hA0; #100;
A = 8'hE8; B = 8'hA1; #100;
A = 8'hE8; B = 8'hA2; #100;
A = 8'hE8; B = 8'hA3; #100;
A = 8'hE8; B = 8'hA4; #100;
A = 8'hE8; B = 8'hA5; #100;
A = 8'hE8; B = 8'hA6; #100;
A = 8'hE8; B = 8'hA7; #100;
A = 8'hE8; B = 8'hA8; #100;
A = 8'hE8; B = 8'hA9; #100;
A = 8'hE8; B = 8'hAA; #100;
A = 8'hE8; B = 8'hAB; #100;
A = 8'hE8; B = 8'hAC; #100;
A = 8'hE8; B = 8'hAD; #100;
A = 8'hE8; B = 8'hAE; #100;
A = 8'hE8; B = 8'hAF; #100;
A = 8'hE8; B = 8'hB0; #100;
A = 8'hE8; B = 8'hB1; #100;
A = 8'hE8; B = 8'hB2; #100;
A = 8'hE8; B = 8'hB3; #100;
A = 8'hE8; B = 8'hB4; #100;
A = 8'hE8; B = 8'hB5; #100;
A = 8'hE8; B = 8'hB6; #100;
A = 8'hE8; B = 8'hB7; #100;
A = 8'hE8; B = 8'hB8; #100;
A = 8'hE8; B = 8'hB9; #100;
A = 8'hE8; B = 8'hBA; #100;
A = 8'hE8; B = 8'hBB; #100;
A = 8'hE8; B = 8'hBC; #100;
A = 8'hE8; B = 8'hBD; #100;
A = 8'hE8; B = 8'hBE; #100;
A = 8'hE8; B = 8'hBF; #100;
A = 8'hE8; B = 8'hC0; #100;
A = 8'hE8; B = 8'hC1; #100;
A = 8'hE8; B = 8'hC2; #100;
A = 8'hE8; B = 8'hC3; #100;
A = 8'hE8; B = 8'hC4; #100;
A = 8'hE8; B = 8'hC5; #100;
A = 8'hE8; B = 8'hC6; #100;
A = 8'hE8; B = 8'hC7; #100;
A = 8'hE8; B = 8'hC8; #100;
A = 8'hE8; B = 8'hC9; #100;
A = 8'hE8; B = 8'hCA; #100;
A = 8'hE8; B = 8'hCB; #100;
A = 8'hE8; B = 8'hCC; #100;
A = 8'hE8; B = 8'hCD; #100;
A = 8'hE8; B = 8'hCE; #100;
A = 8'hE8; B = 8'hCF; #100;
A = 8'hE8; B = 8'hD0; #100;
A = 8'hE8; B = 8'hD1; #100;
A = 8'hE8; B = 8'hD2; #100;
A = 8'hE8; B = 8'hD3; #100;
A = 8'hE8; B = 8'hD4; #100;
A = 8'hE8; B = 8'hD5; #100;
A = 8'hE8; B = 8'hD6; #100;
A = 8'hE8; B = 8'hD7; #100;
A = 8'hE8; B = 8'hD8; #100;
A = 8'hE8; B = 8'hD9; #100;
A = 8'hE8; B = 8'hDA; #100;
A = 8'hE8; B = 8'hDB; #100;
A = 8'hE8; B = 8'hDC; #100;
A = 8'hE8; B = 8'hDD; #100;
A = 8'hE8; B = 8'hDE; #100;
A = 8'hE8; B = 8'hDF; #100;
A = 8'hE8; B = 8'hE0; #100;
A = 8'hE8; B = 8'hE1; #100;
A = 8'hE8; B = 8'hE2; #100;
A = 8'hE8; B = 8'hE3; #100;
A = 8'hE8; B = 8'hE4; #100;
A = 8'hE8; B = 8'hE5; #100;
A = 8'hE8; B = 8'hE6; #100;
A = 8'hE8; B = 8'hE7; #100;
A = 8'hE8; B = 8'hE8; #100;
A = 8'hE8; B = 8'hE9; #100;
A = 8'hE8; B = 8'hEA; #100;
A = 8'hE8; B = 8'hEB; #100;
A = 8'hE8; B = 8'hEC; #100;
A = 8'hE8; B = 8'hED; #100;
A = 8'hE8; B = 8'hEE; #100;
A = 8'hE8; B = 8'hEF; #100;
A = 8'hE8; B = 8'hF0; #100;
A = 8'hE8; B = 8'hF1; #100;
A = 8'hE8; B = 8'hF2; #100;
A = 8'hE8; B = 8'hF3; #100;
A = 8'hE8; B = 8'hF4; #100;
A = 8'hE8; B = 8'hF5; #100;
A = 8'hE8; B = 8'hF6; #100;
A = 8'hE8; B = 8'hF7; #100;
A = 8'hE8; B = 8'hF8; #100;
A = 8'hE8; B = 8'hF9; #100;
A = 8'hE8; B = 8'hFA; #100;
A = 8'hE8; B = 8'hFB; #100;
A = 8'hE8; B = 8'hFC; #100;
A = 8'hE8; B = 8'hFD; #100;
A = 8'hE8; B = 8'hFE; #100;
A = 8'hE8; B = 8'hFF; #100;
A = 8'hE9; B = 8'h0; #100;
A = 8'hE9; B = 8'h1; #100;
A = 8'hE9; B = 8'h2; #100;
A = 8'hE9; B = 8'h3; #100;
A = 8'hE9; B = 8'h4; #100;
A = 8'hE9; B = 8'h5; #100;
A = 8'hE9; B = 8'h6; #100;
A = 8'hE9; B = 8'h7; #100;
A = 8'hE9; B = 8'h8; #100;
A = 8'hE9; B = 8'h9; #100;
A = 8'hE9; B = 8'hA; #100;
A = 8'hE9; B = 8'hB; #100;
A = 8'hE9; B = 8'hC; #100;
A = 8'hE9; B = 8'hD; #100;
A = 8'hE9; B = 8'hE; #100;
A = 8'hE9; B = 8'hF; #100;
A = 8'hE9; B = 8'h10; #100;
A = 8'hE9; B = 8'h11; #100;
A = 8'hE9; B = 8'h12; #100;
A = 8'hE9; B = 8'h13; #100;
A = 8'hE9; B = 8'h14; #100;
A = 8'hE9; B = 8'h15; #100;
A = 8'hE9; B = 8'h16; #100;
A = 8'hE9; B = 8'h17; #100;
A = 8'hE9; B = 8'h18; #100;
A = 8'hE9; B = 8'h19; #100;
A = 8'hE9; B = 8'h1A; #100;
A = 8'hE9; B = 8'h1B; #100;
A = 8'hE9; B = 8'h1C; #100;
A = 8'hE9; B = 8'h1D; #100;
A = 8'hE9; B = 8'h1E; #100;
A = 8'hE9; B = 8'h1F; #100;
A = 8'hE9; B = 8'h20; #100;
A = 8'hE9; B = 8'h21; #100;
A = 8'hE9; B = 8'h22; #100;
A = 8'hE9; B = 8'h23; #100;
A = 8'hE9; B = 8'h24; #100;
A = 8'hE9; B = 8'h25; #100;
A = 8'hE9; B = 8'h26; #100;
A = 8'hE9; B = 8'h27; #100;
A = 8'hE9; B = 8'h28; #100;
A = 8'hE9; B = 8'h29; #100;
A = 8'hE9; B = 8'h2A; #100;
A = 8'hE9; B = 8'h2B; #100;
A = 8'hE9; B = 8'h2C; #100;
A = 8'hE9; B = 8'h2D; #100;
A = 8'hE9; B = 8'h2E; #100;
A = 8'hE9; B = 8'h2F; #100;
A = 8'hE9; B = 8'h30; #100;
A = 8'hE9; B = 8'h31; #100;
A = 8'hE9; B = 8'h32; #100;
A = 8'hE9; B = 8'h33; #100;
A = 8'hE9; B = 8'h34; #100;
A = 8'hE9; B = 8'h35; #100;
A = 8'hE9; B = 8'h36; #100;
A = 8'hE9; B = 8'h37; #100;
A = 8'hE9; B = 8'h38; #100;
A = 8'hE9; B = 8'h39; #100;
A = 8'hE9; B = 8'h3A; #100;
A = 8'hE9; B = 8'h3B; #100;
A = 8'hE9; B = 8'h3C; #100;
A = 8'hE9; B = 8'h3D; #100;
A = 8'hE9; B = 8'h3E; #100;
A = 8'hE9; B = 8'h3F; #100;
A = 8'hE9; B = 8'h40; #100;
A = 8'hE9; B = 8'h41; #100;
A = 8'hE9; B = 8'h42; #100;
A = 8'hE9; B = 8'h43; #100;
A = 8'hE9; B = 8'h44; #100;
A = 8'hE9; B = 8'h45; #100;
A = 8'hE9; B = 8'h46; #100;
A = 8'hE9; B = 8'h47; #100;
A = 8'hE9; B = 8'h48; #100;
A = 8'hE9; B = 8'h49; #100;
A = 8'hE9; B = 8'h4A; #100;
A = 8'hE9; B = 8'h4B; #100;
A = 8'hE9; B = 8'h4C; #100;
A = 8'hE9; B = 8'h4D; #100;
A = 8'hE9; B = 8'h4E; #100;
A = 8'hE9; B = 8'h4F; #100;
A = 8'hE9; B = 8'h50; #100;
A = 8'hE9; B = 8'h51; #100;
A = 8'hE9; B = 8'h52; #100;
A = 8'hE9; B = 8'h53; #100;
A = 8'hE9; B = 8'h54; #100;
A = 8'hE9; B = 8'h55; #100;
A = 8'hE9; B = 8'h56; #100;
A = 8'hE9; B = 8'h57; #100;
A = 8'hE9; B = 8'h58; #100;
A = 8'hE9; B = 8'h59; #100;
A = 8'hE9; B = 8'h5A; #100;
A = 8'hE9; B = 8'h5B; #100;
A = 8'hE9; B = 8'h5C; #100;
A = 8'hE9; B = 8'h5D; #100;
A = 8'hE9; B = 8'h5E; #100;
A = 8'hE9; B = 8'h5F; #100;
A = 8'hE9; B = 8'h60; #100;
A = 8'hE9; B = 8'h61; #100;
A = 8'hE9; B = 8'h62; #100;
A = 8'hE9; B = 8'h63; #100;
A = 8'hE9; B = 8'h64; #100;
A = 8'hE9; B = 8'h65; #100;
A = 8'hE9; B = 8'h66; #100;
A = 8'hE9; B = 8'h67; #100;
A = 8'hE9; B = 8'h68; #100;
A = 8'hE9; B = 8'h69; #100;
A = 8'hE9; B = 8'h6A; #100;
A = 8'hE9; B = 8'h6B; #100;
A = 8'hE9; B = 8'h6C; #100;
A = 8'hE9; B = 8'h6D; #100;
A = 8'hE9; B = 8'h6E; #100;
A = 8'hE9; B = 8'h6F; #100;
A = 8'hE9; B = 8'h70; #100;
A = 8'hE9; B = 8'h71; #100;
A = 8'hE9; B = 8'h72; #100;
A = 8'hE9; B = 8'h73; #100;
A = 8'hE9; B = 8'h74; #100;
A = 8'hE9; B = 8'h75; #100;
A = 8'hE9; B = 8'h76; #100;
A = 8'hE9; B = 8'h77; #100;
A = 8'hE9; B = 8'h78; #100;
A = 8'hE9; B = 8'h79; #100;
A = 8'hE9; B = 8'h7A; #100;
A = 8'hE9; B = 8'h7B; #100;
A = 8'hE9; B = 8'h7C; #100;
A = 8'hE9; B = 8'h7D; #100;
A = 8'hE9; B = 8'h7E; #100;
A = 8'hE9; B = 8'h7F; #100;
A = 8'hE9; B = 8'h80; #100;
A = 8'hE9; B = 8'h81; #100;
A = 8'hE9; B = 8'h82; #100;
A = 8'hE9; B = 8'h83; #100;
A = 8'hE9; B = 8'h84; #100;
A = 8'hE9; B = 8'h85; #100;
A = 8'hE9; B = 8'h86; #100;
A = 8'hE9; B = 8'h87; #100;
A = 8'hE9; B = 8'h88; #100;
A = 8'hE9; B = 8'h89; #100;
A = 8'hE9; B = 8'h8A; #100;
A = 8'hE9; B = 8'h8B; #100;
A = 8'hE9; B = 8'h8C; #100;
A = 8'hE9; B = 8'h8D; #100;
A = 8'hE9; B = 8'h8E; #100;
A = 8'hE9; B = 8'h8F; #100;
A = 8'hE9; B = 8'h90; #100;
A = 8'hE9; B = 8'h91; #100;
A = 8'hE9; B = 8'h92; #100;
A = 8'hE9; B = 8'h93; #100;
A = 8'hE9; B = 8'h94; #100;
A = 8'hE9; B = 8'h95; #100;
A = 8'hE9; B = 8'h96; #100;
A = 8'hE9; B = 8'h97; #100;
A = 8'hE9; B = 8'h98; #100;
A = 8'hE9; B = 8'h99; #100;
A = 8'hE9; B = 8'h9A; #100;
A = 8'hE9; B = 8'h9B; #100;
A = 8'hE9; B = 8'h9C; #100;
A = 8'hE9; B = 8'h9D; #100;
A = 8'hE9; B = 8'h9E; #100;
A = 8'hE9; B = 8'h9F; #100;
A = 8'hE9; B = 8'hA0; #100;
A = 8'hE9; B = 8'hA1; #100;
A = 8'hE9; B = 8'hA2; #100;
A = 8'hE9; B = 8'hA3; #100;
A = 8'hE9; B = 8'hA4; #100;
A = 8'hE9; B = 8'hA5; #100;
A = 8'hE9; B = 8'hA6; #100;
A = 8'hE9; B = 8'hA7; #100;
A = 8'hE9; B = 8'hA8; #100;
A = 8'hE9; B = 8'hA9; #100;
A = 8'hE9; B = 8'hAA; #100;
A = 8'hE9; B = 8'hAB; #100;
A = 8'hE9; B = 8'hAC; #100;
A = 8'hE9; B = 8'hAD; #100;
A = 8'hE9; B = 8'hAE; #100;
A = 8'hE9; B = 8'hAF; #100;
A = 8'hE9; B = 8'hB0; #100;
A = 8'hE9; B = 8'hB1; #100;
A = 8'hE9; B = 8'hB2; #100;
A = 8'hE9; B = 8'hB3; #100;
A = 8'hE9; B = 8'hB4; #100;
A = 8'hE9; B = 8'hB5; #100;
A = 8'hE9; B = 8'hB6; #100;
A = 8'hE9; B = 8'hB7; #100;
A = 8'hE9; B = 8'hB8; #100;
A = 8'hE9; B = 8'hB9; #100;
A = 8'hE9; B = 8'hBA; #100;
A = 8'hE9; B = 8'hBB; #100;
A = 8'hE9; B = 8'hBC; #100;
A = 8'hE9; B = 8'hBD; #100;
A = 8'hE9; B = 8'hBE; #100;
A = 8'hE9; B = 8'hBF; #100;
A = 8'hE9; B = 8'hC0; #100;
A = 8'hE9; B = 8'hC1; #100;
A = 8'hE9; B = 8'hC2; #100;
A = 8'hE9; B = 8'hC3; #100;
A = 8'hE9; B = 8'hC4; #100;
A = 8'hE9; B = 8'hC5; #100;
A = 8'hE9; B = 8'hC6; #100;
A = 8'hE9; B = 8'hC7; #100;
A = 8'hE9; B = 8'hC8; #100;
A = 8'hE9; B = 8'hC9; #100;
A = 8'hE9; B = 8'hCA; #100;
A = 8'hE9; B = 8'hCB; #100;
A = 8'hE9; B = 8'hCC; #100;
A = 8'hE9; B = 8'hCD; #100;
A = 8'hE9; B = 8'hCE; #100;
A = 8'hE9; B = 8'hCF; #100;
A = 8'hE9; B = 8'hD0; #100;
A = 8'hE9; B = 8'hD1; #100;
A = 8'hE9; B = 8'hD2; #100;
A = 8'hE9; B = 8'hD3; #100;
A = 8'hE9; B = 8'hD4; #100;
A = 8'hE9; B = 8'hD5; #100;
A = 8'hE9; B = 8'hD6; #100;
A = 8'hE9; B = 8'hD7; #100;
A = 8'hE9; B = 8'hD8; #100;
A = 8'hE9; B = 8'hD9; #100;
A = 8'hE9; B = 8'hDA; #100;
A = 8'hE9; B = 8'hDB; #100;
A = 8'hE9; B = 8'hDC; #100;
A = 8'hE9; B = 8'hDD; #100;
A = 8'hE9; B = 8'hDE; #100;
A = 8'hE9; B = 8'hDF; #100;
A = 8'hE9; B = 8'hE0; #100;
A = 8'hE9; B = 8'hE1; #100;
A = 8'hE9; B = 8'hE2; #100;
A = 8'hE9; B = 8'hE3; #100;
A = 8'hE9; B = 8'hE4; #100;
A = 8'hE9; B = 8'hE5; #100;
A = 8'hE9; B = 8'hE6; #100;
A = 8'hE9; B = 8'hE7; #100;
A = 8'hE9; B = 8'hE8; #100;
A = 8'hE9; B = 8'hE9; #100;
A = 8'hE9; B = 8'hEA; #100;
A = 8'hE9; B = 8'hEB; #100;
A = 8'hE9; B = 8'hEC; #100;
A = 8'hE9; B = 8'hED; #100;
A = 8'hE9; B = 8'hEE; #100;
A = 8'hE9; B = 8'hEF; #100;
A = 8'hE9; B = 8'hF0; #100;
A = 8'hE9; B = 8'hF1; #100;
A = 8'hE9; B = 8'hF2; #100;
A = 8'hE9; B = 8'hF3; #100;
A = 8'hE9; B = 8'hF4; #100;
A = 8'hE9; B = 8'hF5; #100;
A = 8'hE9; B = 8'hF6; #100;
A = 8'hE9; B = 8'hF7; #100;
A = 8'hE9; B = 8'hF8; #100;
A = 8'hE9; B = 8'hF9; #100;
A = 8'hE9; B = 8'hFA; #100;
A = 8'hE9; B = 8'hFB; #100;
A = 8'hE9; B = 8'hFC; #100;
A = 8'hE9; B = 8'hFD; #100;
A = 8'hE9; B = 8'hFE; #100;
A = 8'hE9; B = 8'hFF; #100;
A = 8'hEA; B = 8'h0; #100;
A = 8'hEA; B = 8'h1; #100;
A = 8'hEA; B = 8'h2; #100;
A = 8'hEA; B = 8'h3; #100;
A = 8'hEA; B = 8'h4; #100;
A = 8'hEA; B = 8'h5; #100;
A = 8'hEA; B = 8'h6; #100;
A = 8'hEA; B = 8'h7; #100;
A = 8'hEA; B = 8'h8; #100;
A = 8'hEA; B = 8'h9; #100;
A = 8'hEA; B = 8'hA; #100;
A = 8'hEA; B = 8'hB; #100;
A = 8'hEA; B = 8'hC; #100;
A = 8'hEA; B = 8'hD; #100;
A = 8'hEA; B = 8'hE; #100;
A = 8'hEA; B = 8'hF; #100;
A = 8'hEA; B = 8'h10; #100;
A = 8'hEA; B = 8'h11; #100;
A = 8'hEA; B = 8'h12; #100;
A = 8'hEA; B = 8'h13; #100;
A = 8'hEA; B = 8'h14; #100;
A = 8'hEA; B = 8'h15; #100;
A = 8'hEA; B = 8'h16; #100;
A = 8'hEA; B = 8'h17; #100;
A = 8'hEA; B = 8'h18; #100;
A = 8'hEA; B = 8'h19; #100;
A = 8'hEA; B = 8'h1A; #100;
A = 8'hEA; B = 8'h1B; #100;
A = 8'hEA; B = 8'h1C; #100;
A = 8'hEA; B = 8'h1D; #100;
A = 8'hEA; B = 8'h1E; #100;
A = 8'hEA; B = 8'h1F; #100;
A = 8'hEA; B = 8'h20; #100;
A = 8'hEA; B = 8'h21; #100;
A = 8'hEA; B = 8'h22; #100;
A = 8'hEA; B = 8'h23; #100;
A = 8'hEA; B = 8'h24; #100;
A = 8'hEA; B = 8'h25; #100;
A = 8'hEA; B = 8'h26; #100;
A = 8'hEA; B = 8'h27; #100;
A = 8'hEA; B = 8'h28; #100;
A = 8'hEA; B = 8'h29; #100;
A = 8'hEA; B = 8'h2A; #100;
A = 8'hEA; B = 8'h2B; #100;
A = 8'hEA; B = 8'h2C; #100;
A = 8'hEA; B = 8'h2D; #100;
A = 8'hEA; B = 8'h2E; #100;
A = 8'hEA; B = 8'h2F; #100;
A = 8'hEA; B = 8'h30; #100;
A = 8'hEA; B = 8'h31; #100;
A = 8'hEA; B = 8'h32; #100;
A = 8'hEA; B = 8'h33; #100;
A = 8'hEA; B = 8'h34; #100;
A = 8'hEA; B = 8'h35; #100;
A = 8'hEA; B = 8'h36; #100;
A = 8'hEA; B = 8'h37; #100;
A = 8'hEA; B = 8'h38; #100;
A = 8'hEA; B = 8'h39; #100;
A = 8'hEA; B = 8'h3A; #100;
A = 8'hEA; B = 8'h3B; #100;
A = 8'hEA; B = 8'h3C; #100;
A = 8'hEA; B = 8'h3D; #100;
A = 8'hEA; B = 8'h3E; #100;
A = 8'hEA; B = 8'h3F; #100;
A = 8'hEA; B = 8'h40; #100;
A = 8'hEA; B = 8'h41; #100;
A = 8'hEA; B = 8'h42; #100;
A = 8'hEA; B = 8'h43; #100;
A = 8'hEA; B = 8'h44; #100;
A = 8'hEA; B = 8'h45; #100;
A = 8'hEA; B = 8'h46; #100;
A = 8'hEA; B = 8'h47; #100;
A = 8'hEA; B = 8'h48; #100;
A = 8'hEA; B = 8'h49; #100;
A = 8'hEA; B = 8'h4A; #100;
A = 8'hEA; B = 8'h4B; #100;
A = 8'hEA; B = 8'h4C; #100;
A = 8'hEA; B = 8'h4D; #100;
A = 8'hEA; B = 8'h4E; #100;
A = 8'hEA; B = 8'h4F; #100;
A = 8'hEA; B = 8'h50; #100;
A = 8'hEA; B = 8'h51; #100;
A = 8'hEA; B = 8'h52; #100;
A = 8'hEA; B = 8'h53; #100;
A = 8'hEA; B = 8'h54; #100;
A = 8'hEA; B = 8'h55; #100;
A = 8'hEA; B = 8'h56; #100;
A = 8'hEA; B = 8'h57; #100;
A = 8'hEA; B = 8'h58; #100;
A = 8'hEA; B = 8'h59; #100;
A = 8'hEA; B = 8'h5A; #100;
A = 8'hEA; B = 8'h5B; #100;
A = 8'hEA; B = 8'h5C; #100;
A = 8'hEA; B = 8'h5D; #100;
A = 8'hEA; B = 8'h5E; #100;
A = 8'hEA; B = 8'h5F; #100;
A = 8'hEA; B = 8'h60; #100;
A = 8'hEA; B = 8'h61; #100;
A = 8'hEA; B = 8'h62; #100;
A = 8'hEA; B = 8'h63; #100;
A = 8'hEA; B = 8'h64; #100;
A = 8'hEA; B = 8'h65; #100;
A = 8'hEA; B = 8'h66; #100;
A = 8'hEA; B = 8'h67; #100;
A = 8'hEA; B = 8'h68; #100;
A = 8'hEA; B = 8'h69; #100;
A = 8'hEA; B = 8'h6A; #100;
A = 8'hEA; B = 8'h6B; #100;
A = 8'hEA; B = 8'h6C; #100;
A = 8'hEA; B = 8'h6D; #100;
A = 8'hEA; B = 8'h6E; #100;
A = 8'hEA; B = 8'h6F; #100;
A = 8'hEA; B = 8'h70; #100;
A = 8'hEA; B = 8'h71; #100;
A = 8'hEA; B = 8'h72; #100;
A = 8'hEA; B = 8'h73; #100;
A = 8'hEA; B = 8'h74; #100;
A = 8'hEA; B = 8'h75; #100;
A = 8'hEA; B = 8'h76; #100;
A = 8'hEA; B = 8'h77; #100;
A = 8'hEA; B = 8'h78; #100;
A = 8'hEA; B = 8'h79; #100;
A = 8'hEA; B = 8'h7A; #100;
A = 8'hEA; B = 8'h7B; #100;
A = 8'hEA; B = 8'h7C; #100;
A = 8'hEA; B = 8'h7D; #100;
A = 8'hEA; B = 8'h7E; #100;
A = 8'hEA; B = 8'h7F; #100;
A = 8'hEA; B = 8'h80; #100;
A = 8'hEA; B = 8'h81; #100;
A = 8'hEA; B = 8'h82; #100;
A = 8'hEA; B = 8'h83; #100;
A = 8'hEA; B = 8'h84; #100;
A = 8'hEA; B = 8'h85; #100;
A = 8'hEA; B = 8'h86; #100;
A = 8'hEA; B = 8'h87; #100;
A = 8'hEA; B = 8'h88; #100;
A = 8'hEA; B = 8'h89; #100;
A = 8'hEA; B = 8'h8A; #100;
A = 8'hEA; B = 8'h8B; #100;
A = 8'hEA; B = 8'h8C; #100;
A = 8'hEA; B = 8'h8D; #100;
A = 8'hEA; B = 8'h8E; #100;
A = 8'hEA; B = 8'h8F; #100;
A = 8'hEA; B = 8'h90; #100;
A = 8'hEA; B = 8'h91; #100;
A = 8'hEA; B = 8'h92; #100;
A = 8'hEA; B = 8'h93; #100;
A = 8'hEA; B = 8'h94; #100;
A = 8'hEA; B = 8'h95; #100;
A = 8'hEA; B = 8'h96; #100;
A = 8'hEA; B = 8'h97; #100;
A = 8'hEA; B = 8'h98; #100;
A = 8'hEA; B = 8'h99; #100;
A = 8'hEA; B = 8'h9A; #100;
A = 8'hEA; B = 8'h9B; #100;
A = 8'hEA; B = 8'h9C; #100;
A = 8'hEA; B = 8'h9D; #100;
A = 8'hEA; B = 8'h9E; #100;
A = 8'hEA; B = 8'h9F; #100;
A = 8'hEA; B = 8'hA0; #100;
A = 8'hEA; B = 8'hA1; #100;
A = 8'hEA; B = 8'hA2; #100;
A = 8'hEA; B = 8'hA3; #100;
A = 8'hEA; B = 8'hA4; #100;
A = 8'hEA; B = 8'hA5; #100;
A = 8'hEA; B = 8'hA6; #100;
A = 8'hEA; B = 8'hA7; #100;
A = 8'hEA; B = 8'hA8; #100;
A = 8'hEA; B = 8'hA9; #100;
A = 8'hEA; B = 8'hAA; #100;
A = 8'hEA; B = 8'hAB; #100;
A = 8'hEA; B = 8'hAC; #100;
A = 8'hEA; B = 8'hAD; #100;
A = 8'hEA; B = 8'hAE; #100;
A = 8'hEA; B = 8'hAF; #100;
A = 8'hEA; B = 8'hB0; #100;
A = 8'hEA; B = 8'hB1; #100;
A = 8'hEA; B = 8'hB2; #100;
A = 8'hEA; B = 8'hB3; #100;
A = 8'hEA; B = 8'hB4; #100;
A = 8'hEA; B = 8'hB5; #100;
A = 8'hEA; B = 8'hB6; #100;
A = 8'hEA; B = 8'hB7; #100;
A = 8'hEA; B = 8'hB8; #100;
A = 8'hEA; B = 8'hB9; #100;
A = 8'hEA; B = 8'hBA; #100;
A = 8'hEA; B = 8'hBB; #100;
A = 8'hEA; B = 8'hBC; #100;
A = 8'hEA; B = 8'hBD; #100;
A = 8'hEA; B = 8'hBE; #100;
A = 8'hEA; B = 8'hBF; #100;
A = 8'hEA; B = 8'hC0; #100;
A = 8'hEA; B = 8'hC1; #100;
A = 8'hEA; B = 8'hC2; #100;
A = 8'hEA; B = 8'hC3; #100;
A = 8'hEA; B = 8'hC4; #100;
A = 8'hEA; B = 8'hC5; #100;
A = 8'hEA; B = 8'hC6; #100;
A = 8'hEA; B = 8'hC7; #100;
A = 8'hEA; B = 8'hC8; #100;
A = 8'hEA; B = 8'hC9; #100;
A = 8'hEA; B = 8'hCA; #100;
A = 8'hEA; B = 8'hCB; #100;
A = 8'hEA; B = 8'hCC; #100;
A = 8'hEA; B = 8'hCD; #100;
A = 8'hEA; B = 8'hCE; #100;
A = 8'hEA; B = 8'hCF; #100;
A = 8'hEA; B = 8'hD0; #100;
A = 8'hEA; B = 8'hD1; #100;
A = 8'hEA; B = 8'hD2; #100;
A = 8'hEA; B = 8'hD3; #100;
A = 8'hEA; B = 8'hD4; #100;
A = 8'hEA; B = 8'hD5; #100;
A = 8'hEA; B = 8'hD6; #100;
A = 8'hEA; B = 8'hD7; #100;
A = 8'hEA; B = 8'hD8; #100;
A = 8'hEA; B = 8'hD9; #100;
A = 8'hEA; B = 8'hDA; #100;
A = 8'hEA; B = 8'hDB; #100;
A = 8'hEA; B = 8'hDC; #100;
A = 8'hEA; B = 8'hDD; #100;
A = 8'hEA; B = 8'hDE; #100;
A = 8'hEA; B = 8'hDF; #100;
A = 8'hEA; B = 8'hE0; #100;
A = 8'hEA; B = 8'hE1; #100;
A = 8'hEA; B = 8'hE2; #100;
A = 8'hEA; B = 8'hE3; #100;
A = 8'hEA; B = 8'hE4; #100;
A = 8'hEA; B = 8'hE5; #100;
A = 8'hEA; B = 8'hE6; #100;
A = 8'hEA; B = 8'hE7; #100;
A = 8'hEA; B = 8'hE8; #100;
A = 8'hEA; B = 8'hE9; #100;
A = 8'hEA; B = 8'hEA; #100;
A = 8'hEA; B = 8'hEB; #100;
A = 8'hEA; B = 8'hEC; #100;
A = 8'hEA; B = 8'hED; #100;
A = 8'hEA; B = 8'hEE; #100;
A = 8'hEA; B = 8'hEF; #100;
A = 8'hEA; B = 8'hF0; #100;
A = 8'hEA; B = 8'hF1; #100;
A = 8'hEA; B = 8'hF2; #100;
A = 8'hEA; B = 8'hF3; #100;
A = 8'hEA; B = 8'hF4; #100;
A = 8'hEA; B = 8'hF5; #100;
A = 8'hEA; B = 8'hF6; #100;
A = 8'hEA; B = 8'hF7; #100;
A = 8'hEA; B = 8'hF8; #100;
A = 8'hEA; B = 8'hF9; #100;
A = 8'hEA; B = 8'hFA; #100;
A = 8'hEA; B = 8'hFB; #100;
A = 8'hEA; B = 8'hFC; #100;
A = 8'hEA; B = 8'hFD; #100;
A = 8'hEA; B = 8'hFE; #100;
A = 8'hEA; B = 8'hFF; #100;
A = 8'hEB; B = 8'h0; #100;
A = 8'hEB; B = 8'h1; #100;
A = 8'hEB; B = 8'h2; #100;
A = 8'hEB; B = 8'h3; #100;
A = 8'hEB; B = 8'h4; #100;
A = 8'hEB; B = 8'h5; #100;
A = 8'hEB; B = 8'h6; #100;
A = 8'hEB; B = 8'h7; #100;
A = 8'hEB; B = 8'h8; #100;
A = 8'hEB; B = 8'h9; #100;
A = 8'hEB; B = 8'hA; #100;
A = 8'hEB; B = 8'hB; #100;
A = 8'hEB; B = 8'hC; #100;
A = 8'hEB; B = 8'hD; #100;
A = 8'hEB; B = 8'hE; #100;
A = 8'hEB; B = 8'hF; #100;
A = 8'hEB; B = 8'h10; #100;
A = 8'hEB; B = 8'h11; #100;
A = 8'hEB; B = 8'h12; #100;
A = 8'hEB; B = 8'h13; #100;
A = 8'hEB; B = 8'h14; #100;
A = 8'hEB; B = 8'h15; #100;
A = 8'hEB; B = 8'h16; #100;
A = 8'hEB; B = 8'h17; #100;
A = 8'hEB; B = 8'h18; #100;
A = 8'hEB; B = 8'h19; #100;
A = 8'hEB; B = 8'h1A; #100;
A = 8'hEB; B = 8'h1B; #100;
A = 8'hEB; B = 8'h1C; #100;
A = 8'hEB; B = 8'h1D; #100;
A = 8'hEB; B = 8'h1E; #100;
A = 8'hEB; B = 8'h1F; #100;
A = 8'hEB; B = 8'h20; #100;
A = 8'hEB; B = 8'h21; #100;
A = 8'hEB; B = 8'h22; #100;
A = 8'hEB; B = 8'h23; #100;
A = 8'hEB; B = 8'h24; #100;
A = 8'hEB; B = 8'h25; #100;
A = 8'hEB; B = 8'h26; #100;
A = 8'hEB; B = 8'h27; #100;
A = 8'hEB; B = 8'h28; #100;
A = 8'hEB; B = 8'h29; #100;
A = 8'hEB; B = 8'h2A; #100;
A = 8'hEB; B = 8'h2B; #100;
A = 8'hEB; B = 8'h2C; #100;
A = 8'hEB; B = 8'h2D; #100;
A = 8'hEB; B = 8'h2E; #100;
A = 8'hEB; B = 8'h2F; #100;
A = 8'hEB; B = 8'h30; #100;
A = 8'hEB; B = 8'h31; #100;
A = 8'hEB; B = 8'h32; #100;
A = 8'hEB; B = 8'h33; #100;
A = 8'hEB; B = 8'h34; #100;
A = 8'hEB; B = 8'h35; #100;
A = 8'hEB; B = 8'h36; #100;
A = 8'hEB; B = 8'h37; #100;
A = 8'hEB; B = 8'h38; #100;
A = 8'hEB; B = 8'h39; #100;
A = 8'hEB; B = 8'h3A; #100;
A = 8'hEB; B = 8'h3B; #100;
A = 8'hEB; B = 8'h3C; #100;
A = 8'hEB; B = 8'h3D; #100;
A = 8'hEB; B = 8'h3E; #100;
A = 8'hEB; B = 8'h3F; #100;
A = 8'hEB; B = 8'h40; #100;
A = 8'hEB; B = 8'h41; #100;
A = 8'hEB; B = 8'h42; #100;
A = 8'hEB; B = 8'h43; #100;
A = 8'hEB; B = 8'h44; #100;
A = 8'hEB; B = 8'h45; #100;
A = 8'hEB; B = 8'h46; #100;
A = 8'hEB; B = 8'h47; #100;
A = 8'hEB; B = 8'h48; #100;
A = 8'hEB; B = 8'h49; #100;
A = 8'hEB; B = 8'h4A; #100;
A = 8'hEB; B = 8'h4B; #100;
A = 8'hEB; B = 8'h4C; #100;
A = 8'hEB; B = 8'h4D; #100;
A = 8'hEB; B = 8'h4E; #100;
A = 8'hEB; B = 8'h4F; #100;
A = 8'hEB; B = 8'h50; #100;
A = 8'hEB; B = 8'h51; #100;
A = 8'hEB; B = 8'h52; #100;
A = 8'hEB; B = 8'h53; #100;
A = 8'hEB; B = 8'h54; #100;
A = 8'hEB; B = 8'h55; #100;
A = 8'hEB; B = 8'h56; #100;
A = 8'hEB; B = 8'h57; #100;
A = 8'hEB; B = 8'h58; #100;
A = 8'hEB; B = 8'h59; #100;
A = 8'hEB; B = 8'h5A; #100;
A = 8'hEB; B = 8'h5B; #100;
A = 8'hEB; B = 8'h5C; #100;
A = 8'hEB; B = 8'h5D; #100;
A = 8'hEB; B = 8'h5E; #100;
A = 8'hEB; B = 8'h5F; #100;
A = 8'hEB; B = 8'h60; #100;
A = 8'hEB; B = 8'h61; #100;
A = 8'hEB; B = 8'h62; #100;
A = 8'hEB; B = 8'h63; #100;
A = 8'hEB; B = 8'h64; #100;
A = 8'hEB; B = 8'h65; #100;
A = 8'hEB; B = 8'h66; #100;
A = 8'hEB; B = 8'h67; #100;
A = 8'hEB; B = 8'h68; #100;
A = 8'hEB; B = 8'h69; #100;
A = 8'hEB; B = 8'h6A; #100;
A = 8'hEB; B = 8'h6B; #100;
A = 8'hEB; B = 8'h6C; #100;
A = 8'hEB; B = 8'h6D; #100;
A = 8'hEB; B = 8'h6E; #100;
A = 8'hEB; B = 8'h6F; #100;
A = 8'hEB; B = 8'h70; #100;
A = 8'hEB; B = 8'h71; #100;
A = 8'hEB; B = 8'h72; #100;
A = 8'hEB; B = 8'h73; #100;
A = 8'hEB; B = 8'h74; #100;
A = 8'hEB; B = 8'h75; #100;
A = 8'hEB; B = 8'h76; #100;
A = 8'hEB; B = 8'h77; #100;
A = 8'hEB; B = 8'h78; #100;
A = 8'hEB; B = 8'h79; #100;
A = 8'hEB; B = 8'h7A; #100;
A = 8'hEB; B = 8'h7B; #100;
A = 8'hEB; B = 8'h7C; #100;
A = 8'hEB; B = 8'h7D; #100;
A = 8'hEB; B = 8'h7E; #100;
A = 8'hEB; B = 8'h7F; #100;
A = 8'hEB; B = 8'h80; #100;
A = 8'hEB; B = 8'h81; #100;
A = 8'hEB; B = 8'h82; #100;
A = 8'hEB; B = 8'h83; #100;
A = 8'hEB; B = 8'h84; #100;
A = 8'hEB; B = 8'h85; #100;
A = 8'hEB; B = 8'h86; #100;
A = 8'hEB; B = 8'h87; #100;
A = 8'hEB; B = 8'h88; #100;
A = 8'hEB; B = 8'h89; #100;
A = 8'hEB; B = 8'h8A; #100;
A = 8'hEB; B = 8'h8B; #100;
A = 8'hEB; B = 8'h8C; #100;
A = 8'hEB; B = 8'h8D; #100;
A = 8'hEB; B = 8'h8E; #100;
A = 8'hEB; B = 8'h8F; #100;
A = 8'hEB; B = 8'h90; #100;
A = 8'hEB; B = 8'h91; #100;
A = 8'hEB; B = 8'h92; #100;
A = 8'hEB; B = 8'h93; #100;
A = 8'hEB; B = 8'h94; #100;
A = 8'hEB; B = 8'h95; #100;
A = 8'hEB; B = 8'h96; #100;
A = 8'hEB; B = 8'h97; #100;
A = 8'hEB; B = 8'h98; #100;
A = 8'hEB; B = 8'h99; #100;
A = 8'hEB; B = 8'h9A; #100;
A = 8'hEB; B = 8'h9B; #100;
A = 8'hEB; B = 8'h9C; #100;
A = 8'hEB; B = 8'h9D; #100;
A = 8'hEB; B = 8'h9E; #100;
A = 8'hEB; B = 8'h9F; #100;
A = 8'hEB; B = 8'hA0; #100;
A = 8'hEB; B = 8'hA1; #100;
A = 8'hEB; B = 8'hA2; #100;
A = 8'hEB; B = 8'hA3; #100;
A = 8'hEB; B = 8'hA4; #100;
A = 8'hEB; B = 8'hA5; #100;
A = 8'hEB; B = 8'hA6; #100;
A = 8'hEB; B = 8'hA7; #100;
A = 8'hEB; B = 8'hA8; #100;
A = 8'hEB; B = 8'hA9; #100;
A = 8'hEB; B = 8'hAA; #100;
A = 8'hEB; B = 8'hAB; #100;
A = 8'hEB; B = 8'hAC; #100;
A = 8'hEB; B = 8'hAD; #100;
A = 8'hEB; B = 8'hAE; #100;
A = 8'hEB; B = 8'hAF; #100;
A = 8'hEB; B = 8'hB0; #100;
A = 8'hEB; B = 8'hB1; #100;
A = 8'hEB; B = 8'hB2; #100;
A = 8'hEB; B = 8'hB3; #100;
A = 8'hEB; B = 8'hB4; #100;
A = 8'hEB; B = 8'hB5; #100;
A = 8'hEB; B = 8'hB6; #100;
A = 8'hEB; B = 8'hB7; #100;
A = 8'hEB; B = 8'hB8; #100;
A = 8'hEB; B = 8'hB9; #100;
A = 8'hEB; B = 8'hBA; #100;
A = 8'hEB; B = 8'hBB; #100;
A = 8'hEB; B = 8'hBC; #100;
A = 8'hEB; B = 8'hBD; #100;
A = 8'hEB; B = 8'hBE; #100;
A = 8'hEB; B = 8'hBF; #100;
A = 8'hEB; B = 8'hC0; #100;
A = 8'hEB; B = 8'hC1; #100;
A = 8'hEB; B = 8'hC2; #100;
A = 8'hEB; B = 8'hC3; #100;
A = 8'hEB; B = 8'hC4; #100;
A = 8'hEB; B = 8'hC5; #100;
A = 8'hEB; B = 8'hC6; #100;
A = 8'hEB; B = 8'hC7; #100;
A = 8'hEB; B = 8'hC8; #100;
A = 8'hEB; B = 8'hC9; #100;
A = 8'hEB; B = 8'hCA; #100;
A = 8'hEB; B = 8'hCB; #100;
A = 8'hEB; B = 8'hCC; #100;
A = 8'hEB; B = 8'hCD; #100;
A = 8'hEB; B = 8'hCE; #100;
A = 8'hEB; B = 8'hCF; #100;
A = 8'hEB; B = 8'hD0; #100;
A = 8'hEB; B = 8'hD1; #100;
A = 8'hEB; B = 8'hD2; #100;
A = 8'hEB; B = 8'hD3; #100;
A = 8'hEB; B = 8'hD4; #100;
A = 8'hEB; B = 8'hD5; #100;
A = 8'hEB; B = 8'hD6; #100;
A = 8'hEB; B = 8'hD7; #100;
A = 8'hEB; B = 8'hD8; #100;
A = 8'hEB; B = 8'hD9; #100;
A = 8'hEB; B = 8'hDA; #100;
A = 8'hEB; B = 8'hDB; #100;
A = 8'hEB; B = 8'hDC; #100;
A = 8'hEB; B = 8'hDD; #100;
A = 8'hEB; B = 8'hDE; #100;
A = 8'hEB; B = 8'hDF; #100;
A = 8'hEB; B = 8'hE0; #100;
A = 8'hEB; B = 8'hE1; #100;
A = 8'hEB; B = 8'hE2; #100;
A = 8'hEB; B = 8'hE3; #100;
A = 8'hEB; B = 8'hE4; #100;
A = 8'hEB; B = 8'hE5; #100;
A = 8'hEB; B = 8'hE6; #100;
A = 8'hEB; B = 8'hE7; #100;
A = 8'hEB; B = 8'hE8; #100;
A = 8'hEB; B = 8'hE9; #100;
A = 8'hEB; B = 8'hEA; #100;
A = 8'hEB; B = 8'hEB; #100;
A = 8'hEB; B = 8'hEC; #100;
A = 8'hEB; B = 8'hED; #100;
A = 8'hEB; B = 8'hEE; #100;
A = 8'hEB; B = 8'hEF; #100;
A = 8'hEB; B = 8'hF0; #100;
A = 8'hEB; B = 8'hF1; #100;
A = 8'hEB; B = 8'hF2; #100;
A = 8'hEB; B = 8'hF3; #100;
A = 8'hEB; B = 8'hF4; #100;
A = 8'hEB; B = 8'hF5; #100;
A = 8'hEB; B = 8'hF6; #100;
A = 8'hEB; B = 8'hF7; #100;
A = 8'hEB; B = 8'hF8; #100;
A = 8'hEB; B = 8'hF9; #100;
A = 8'hEB; B = 8'hFA; #100;
A = 8'hEB; B = 8'hFB; #100;
A = 8'hEB; B = 8'hFC; #100;
A = 8'hEB; B = 8'hFD; #100;
A = 8'hEB; B = 8'hFE; #100;
A = 8'hEB; B = 8'hFF; #100;
A = 8'hEC; B = 8'h0; #100;
A = 8'hEC; B = 8'h1; #100;
A = 8'hEC; B = 8'h2; #100;
A = 8'hEC; B = 8'h3; #100;
A = 8'hEC; B = 8'h4; #100;
A = 8'hEC; B = 8'h5; #100;
A = 8'hEC; B = 8'h6; #100;
A = 8'hEC; B = 8'h7; #100;
A = 8'hEC; B = 8'h8; #100;
A = 8'hEC; B = 8'h9; #100;
A = 8'hEC; B = 8'hA; #100;
A = 8'hEC; B = 8'hB; #100;
A = 8'hEC; B = 8'hC; #100;
A = 8'hEC; B = 8'hD; #100;
A = 8'hEC; B = 8'hE; #100;
A = 8'hEC; B = 8'hF; #100;
A = 8'hEC; B = 8'h10; #100;
A = 8'hEC; B = 8'h11; #100;
A = 8'hEC; B = 8'h12; #100;
A = 8'hEC; B = 8'h13; #100;
A = 8'hEC; B = 8'h14; #100;
A = 8'hEC; B = 8'h15; #100;
A = 8'hEC; B = 8'h16; #100;
A = 8'hEC; B = 8'h17; #100;
A = 8'hEC; B = 8'h18; #100;
A = 8'hEC; B = 8'h19; #100;
A = 8'hEC; B = 8'h1A; #100;
A = 8'hEC; B = 8'h1B; #100;
A = 8'hEC; B = 8'h1C; #100;
A = 8'hEC; B = 8'h1D; #100;
A = 8'hEC; B = 8'h1E; #100;
A = 8'hEC; B = 8'h1F; #100;
A = 8'hEC; B = 8'h20; #100;
A = 8'hEC; B = 8'h21; #100;
A = 8'hEC; B = 8'h22; #100;
A = 8'hEC; B = 8'h23; #100;
A = 8'hEC; B = 8'h24; #100;
A = 8'hEC; B = 8'h25; #100;
A = 8'hEC; B = 8'h26; #100;
A = 8'hEC; B = 8'h27; #100;
A = 8'hEC; B = 8'h28; #100;
A = 8'hEC; B = 8'h29; #100;
A = 8'hEC; B = 8'h2A; #100;
A = 8'hEC; B = 8'h2B; #100;
A = 8'hEC; B = 8'h2C; #100;
A = 8'hEC; B = 8'h2D; #100;
A = 8'hEC; B = 8'h2E; #100;
A = 8'hEC; B = 8'h2F; #100;
A = 8'hEC; B = 8'h30; #100;
A = 8'hEC; B = 8'h31; #100;
A = 8'hEC; B = 8'h32; #100;
A = 8'hEC; B = 8'h33; #100;
A = 8'hEC; B = 8'h34; #100;
A = 8'hEC; B = 8'h35; #100;
A = 8'hEC; B = 8'h36; #100;
A = 8'hEC; B = 8'h37; #100;
A = 8'hEC; B = 8'h38; #100;
A = 8'hEC; B = 8'h39; #100;
A = 8'hEC; B = 8'h3A; #100;
A = 8'hEC; B = 8'h3B; #100;
A = 8'hEC; B = 8'h3C; #100;
A = 8'hEC; B = 8'h3D; #100;
A = 8'hEC; B = 8'h3E; #100;
A = 8'hEC; B = 8'h3F; #100;
A = 8'hEC; B = 8'h40; #100;
A = 8'hEC; B = 8'h41; #100;
A = 8'hEC; B = 8'h42; #100;
A = 8'hEC; B = 8'h43; #100;
A = 8'hEC; B = 8'h44; #100;
A = 8'hEC; B = 8'h45; #100;
A = 8'hEC; B = 8'h46; #100;
A = 8'hEC; B = 8'h47; #100;
A = 8'hEC; B = 8'h48; #100;
A = 8'hEC; B = 8'h49; #100;
A = 8'hEC; B = 8'h4A; #100;
A = 8'hEC; B = 8'h4B; #100;
A = 8'hEC; B = 8'h4C; #100;
A = 8'hEC; B = 8'h4D; #100;
A = 8'hEC; B = 8'h4E; #100;
A = 8'hEC; B = 8'h4F; #100;
A = 8'hEC; B = 8'h50; #100;
A = 8'hEC; B = 8'h51; #100;
A = 8'hEC; B = 8'h52; #100;
A = 8'hEC; B = 8'h53; #100;
A = 8'hEC; B = 8'h54; #100;
A = 8'hEC; B = 8'h55; #100;
A = 8'hEC; B = 8'h56; #100;
A = 8'hEC; B = 8'h57; #100;
A = 8'hEC; B = 8'h58; #100;
A = 8'hEC; B = 8'h59; #100;
A = 8'hEC; B = 8'h5A; #100;
A = 8'hEC; B = 8'h5B; #100;
A = 8'hEC; B = 8'h5C; #100;
A = 8'hEC; B = 8'h5D; #100;
A = 8'hEC; B = 8'h5E; #100;
A = 8'hEC; B = 8'h5F; #100;
A = 8'hEC; B = 8'h60; #100;
A = 8'hEC; B = 8'h61; #100;
A = 8'hEC; B = 8'h62; #100;
A = 8'hEC; B = 8'h63; #100;
A = 8'hEC; B = 8'h64; #100;
A = 8'hEC; B = 8'h65; #100;
A = 8'hEC; B = 8'h66; #100;
A = 8'hEC; B = 8'h67; #100;
A = 8'hEC; B = 8'h68; #100;
A = 8'hEC; B = 8'h69; #100;
A = 8'hEC; B = 8'h6A; #100;
A = 8'hEC; B = 8'h6B; #100;
A = 8'hEC; B = 8'h6C; #100;
A = 8'hEC; B = 8'h6D; #100;
A = 8'hEC; B = 8'h6E; #100;
A = 8'hEC; B = 8'h6F; #100;
A = 8'hEC; B = 8'h70; #100;
A = 8'hEC; B = 8'h71; #100;
A = 8'hEC; B = 8'h72; #100;
A = 8'hEC; B = 8'h73; #100;
A = 8'hEC; B = 8'h74; #100;
A = 8'hEC; B = 8'h75; #100;
A = 8'hEC; B = 8'h76; #100;
A = 8'hEC; B = 8'h77; #100;
A = 8'hEC; B = 8'h78; #100;
A = 8'hEC; B = 8'h79; #100;
A = 8'hEC; B = 8'h7A; #100;
A = 8'hEC; B = 8'h7B; #100;
A = 8'hEC; B = 8'h7C; #100;
A = 8'hEC; B = 8'h7D; #100;
A = 8'hEC; B = 8'h7E; #100;
A = 8'hEC; B = 8'h7F; #100;
A = 8'hEC; B = 8'h80; #100;
A = 8'hEC; B = 8'h81; #100;
A = 8'hEC; B = 8'h82; #100;
A = 8'hEC; B = 8'h83; #100;
A = 8'hEC; B = 8'h84; #100;
A = 8'hEC; B = 8'h85; #100;
A = 8'hEC; B = 8'h86; #100;
A = 8'hEC; B = 8'h87; #100;
A = 8'hEC; B = 8'h88; #100;
A = 8'hEC; B = 8'h89; #100;
A = 8'hEC; B = 8'h8A; #100;
A = 8'hEC; B = 8'h8B; #100;
A = 8'hEC; B = 8'h8C; #100;
A = 8'hEC; B = 8'h8D; #100;
A = 8'hEC; B = 8'h8E; #100;
A = 8'hEC; B = 8'h8F; #100;
A = 8'hEC; B = 8'h90; #100;
A = 8'hEC; B = 8'h91; #100;
A = 8'hEC; B = 8'h92; #100;
A = 8'hEC; B = 8'h93; #100;
A = 8'hEC; B = 8'h94; #100;
A = 8'hEC; B = 8'h95; #100;
A = 8'hEC; B = 8'h96; #100;
A = 8'hEC; B = 8'h97; #100;
A = 8'hEC; B = 8'h98; #100;
A = 8'hEC; B = 8'h99; #100;
A = 8'hEC; B = 8'h9A; #100;
A = 8'hEC; B = 8'h9B; #100;
A = 8'hEC; B = 8'h9C; #100;
A = 8'hEC; B = 8'h9D; #100;
A = 8'hEC; B = 8'h9E; #100;
A = 8'hEC; B = 8'h9F; #100;
A = 8'hEC; B = 8'hA0; #100;
A = 8'hEC; B = 8'hA1; #100;
A = 8'hEC; B = 8'hA2; #100;
A = 8'hEC; B = 8'hA3; #100;
A = 8'hEC; B = 8'hA4; #100;
A = 8'hEC; B = 8'hA5; #100;
A = 8'hEC; B = 8'hA6; #100;
A = 8'hEC; B = 8'hA7; #100;
A = 8'hEC; B = 8'hA8; #100;
A = 8'hEC; B = 8'hA9; #100;
A = 8'hEC; B = 8'hAA; #100;
A = 8'hEC; B = 8'hAB; #100;
A = 8'hEC; B = 8'hAC; #100;
A = 8'hEC; B = 8'hAD; #100;
A = 8'hEC; B = 8'hAE; #100;
A = 8'hEC; B = 8'hAF; #100;
A = 8'hEC; B = 8'hB0; #100;
A = 8'hEC; B = 8'hB1; #100;
A = 8'hEC; B = 8'hB2; #100;
A = 8'hEC; B = 8'hB3; #100;
A = 8'hEC; B = 8'hB4; #100;
A = 8'hEC; B = 8'hB5; #100;
A = 8'hEC; B = 8'hB6; #100;
A = 8'hEC; B = 8'hB7; #100;
A = 8'hEC; B = 8'hB8; #100;
A = 8'hEC; B = 8'hB9; #100;
A = 8'hEC; B = 8'hBA; #100;
A = 8'hEC; B = 8'hBB; #100;
A = 8'hEC; B = 8'hBC; #100;
A = 8'hEC; B = 8'hBD; #100;
A = 8'hEC; B = 8'hBE; #100;
A = 8'hEC; B = 8'hBF; #100;
A = 8'hEC; B = 8'hC0; #100;
A = 8'hEC; B = 8'hC1; #100;
A = 8'hEC; B = 8'hC2; #100;
A = 8'hEC; B = 8'hC3; #100;
A = 8'hEC; B = 8'hC4; #100;
A = 8'hEC; B = 8'hC5; #100;
A = 8'hEC; B = 8'hC6; #100;
A = 8'hEC; B = 8'hC7; #100;
A = 8'hEC; B = 8'hC8; #100;
A = 8'hEC; B = 8'hC9; #100;
A = 8'hEC; B = 8'hCA; #100;
A = 8'hEC; B = 8'hCB; #100;
A = 8'hEC; B = 8'hCC; #100;
A = 8'hEC; B = 8'hCD; #100;
A = 8'hEC; B = 8'hCE; #100;
A = 8'hEC; B = 8'hCF; #100;
A = 8'hEC; B = 8'hD0; #100;
A = 8'hEC; B = 8'hD1; #100;
A = 8'hEC; B = 8'hD2; #100;
A = 8'hEC; B = 8'hD3; #100;
A = 8'hEC; B = 8'hD4; #100;
A = 8'hEC; B = 8'hD5; #100;
A = 8'hEC; B = 8'hD6; #100;
A = 8'hEC; B = 8'hD7; #100;
A = 8'hEC; B = 8'hD8; #100;
A = 8'hEC; B = 8'hD9; #100;
A = 8'hEC; B = 8'hDA; #100;
A = 8'hEC; B = 8'hDB; #100;
A = 8'hEC; B = 8'hDC; #100;
A = 8'hEC; B = 8'hDD; #100;
A = 8'hEC; B = 8'hDE; #100;
A = 8'hEC; B = 8'hDF; #100;
A = 8'hEC; B = 8'hE0; #100;
A = 8'hEC; B = 8'hE1; #100;
A = 8'hEC; B = 8'hE2; #100;
A = 8'hEC; B = 8'hE3; #100;
A = 8'hEC; B = 8'hE4; #100;
A = 8'hEC; B = 8'hE5; #100;
A = 8'hEC; B = 8'hE6; #100;
A = 8'hEC; B = 8'hE7; #100;
A = 8'hEC; B = 8'hE8; #100;
A = 8'hEC; B = 8'hE9; #100;
A = 8'hEC; B = 8'hEA; #100;
A = 8'hEC; B = 8'hEB; #100;
A = 8'hEC; B = 8'hEC; #100;
A = 8'hEC; B = 8'hED; #100;
A = 8'hEC; B = 8'hEE; #100;
A = 8'hEC; B = 8'hEF; #100;
A = 8'hEC; B = 8'hF0; #100;
A = 8'hEC; B = 8'hF1; #100;
A = 8'hEC; B = 8'hF2; #100;
A = 8'hEC; B = 8'hF3; #100;
A = 8'hEC; B = 8'hF4; #100;
A = 8'hEC; B = 8'hF5; #100;
A = 8'hEC; B = 8'hF6; #100;
A = 8'hEC; B = 8'hF7; #100;
A = 8'hEC; B = 8'hF8; #100;
A = 8'hEC; B = 8'hF9; #100;
A = 8'hEC; B = 8'hFA; #100;
A = 8'hEC; B = 8'hFB; #100;
A = 8'hEC; B = 8'hFC; #100;
A = 8'hEC; B = 8'hFD; #100;
A = 8'hEC; B = 8'hFE; #100;
A = 8'hEC; B = 8'hFF; #100;
A = 8'hED; B = 8'h0; #100;
A = 8'hED; B = 8'h1; #100;
A = 8'hED; B = 8'h2; #100;
A = 8'hED; B = 8'h3; #100;
A = 8'hED; B = 8'h4; #100;
A = 8'hED; B = 8'h5; #100;
A = 8'hED; B = 8'h6; #100;
A = 8'hED; B = 8'h7; #100;
A = 8'hED; B = 8'h8; #100;
A = 8'hED; B = 8'h9; #100;
A = 8'hED; B = 8'hA; #100;
A = 8'hED; B = 8'hB; #100;
A = 8'hED; B = 8'hC; #100;
A = 8'hED; B = 8'hD; #100;
A = 8'hED; B = 8'hE; #100;
A = 8'hED; B = 8'hF; #100;
A = 8'hED; B = 8'h10; #100;
A = 8'hED; B = 8'h11; #100;
A = 8'hED; B = 8'h12; #100;
A = 8'hED; B = 8'h13; #100;
A = 8'hED; B = 8'h14; #100;
A = 8'hED; B = 8'h15; #100;
A = 8'hED; B = 8'h16; #100;
A = 8'hED; B = 8'h17; #100;
A = 8'hED; B = 8'h18; #100;
A = 8'hED; B = 8'h19; #100;
A = 8'hED; B = 8'h1A; #100;
A = 8'hED; B = 8'h1B; #100;
A = 8'hED; B = 8'h1C; #100;
A = 8'hED; B = 8'h1D; #100;
A = 8'hED; B = 8'h1E; #100;
A = 8'hED; B = 8'h1F; #100;
A = 8'hED; B = 8'h20; #100;
A = 8'hED; B = 8'h21; #100;
A = 8'hED; B = 8'h22; #100;
A = 8'hED; B = 8'h23; #100;
A = 8'hED; B = 8'h24; #100;
A = 8'hED; B = 8'h25; #100;
A = 8'hED; B = 8'h26; #100;
A = 8'hED; B = 8'h27; #100;
A = 8'hED; B = 8'h28; #100;
A = 8'hED; B = 8'h29; #100;
A = 8'hED; B = 8'h2A; #100;
A = 8'hED; B = 8'h2B; #100;
A = 8'hED; B = 8'h2C; #100;
A = 8'hED; B = 8'h2D; #100;
A = 8'hED; B = 8'h2E; #100;
A = 8'hED; B = 8'h2F; #100;
A = 8'hED; B = 8'h30; #100;
A = 8'hED; B = 8'h31; #100;
A = 8'hED; B = 8'h32; #100;
A = 8'hED; B = 8'h33; #100;
A = 8'hED; B = 8'h34; #100;
A = 8'hED; B = 8'h35; #100;
A = 8'hED; B = 8'h36; #100;
A = 8'hED; B = 8'h37; #100;
A = 8'hED; B = 8'h38; #100;
A = 8'hED; B = 8'h39; #100;
A = 8'hED; B = 8'h3A; #100;
A = 8'hED; B = 8'h3B; #100;
A = 8'hED; B = 8'h3C; #100;
A = 8'hED; B = 8'h3D; #100;
A = 8'hED; B = 8'h3E; #100;
A = 8'hED; B = 8'h3F; #100;
A = 8'hED; B = 8'h40; #100;
A = 8'hED; B = 8'h41; #100;
A = 8'hED; B = 8'h42; #100;
A = 8'hED; B = 8'h43; #100;
A = 8'hED; B = 8'h44; #100;
A = 8'hED; B = 8'h45; #100;
A = 8'hED; B = 8'h46; #100;
A = 8'hED; B = 8'h47; #100;
A = 8'hED; B = 8'h48; #100;
A = 8'hED; B = 8'h49; #100;
A = 8'hED; B = 8'h4A; #100;
A = 8'hED; B = 8'h4B; #100;
A = 8'hED; B = 8'h4C; #100;
A = 8'hED; B = 8'h4D; #100;
A = 8'hED; B = 8'h4E; #100;
A = 8'hED; B = 8'h4F; #100;
A = 8'hED; B = 8'h50; #100;
A = 8'hED; B = 8'h51; #100;
A = 8'hED; B = 8'h52; #100;
A = 8'hED; B = 8'h53; #100;
A = 8'hED; B = 8'h54; #100;
A = 8'hED; B = 8'h55; #100;
A = 8'hED; B = 8'h56; #100;
A = 8'hED; B = 8'h57; #100;
A = 8'hED; B = 8'h58; #100;
A = 8'hED; B = 8'h59; #100;
A = 8'hED; B = 8'h5A; #100;
A = 8'hED; B = 8'h5B; #100;
A = 8'hED; B = 8'h5C; #100;
A = 8'hED; B = 8'h5D; #100;
A = 8'hED; B = 8'h5E; #100;
A = 8'hED; B = 8'h5F; #100;
A = 8'hED; B = 8'h60; #100;
A = 8'hED; B = 8'h61; #100;
A = 8'hED; B = 8'h62; #100;
A = 8'hED; B = 8'h63; #100;
A = 8'hED; B = 8'h64; #100;
A = 8'hED; B = 8'h65; #100;
A = 8'hED; B = 8'h66; #100;
A = 8'hED; B = 8'h67; #100;
A = 8'hED; B = 8'h68; #100;
A = 8'hED; B = 8'h69; #100;
A = 8'hED; B = 8'h6A; #100;
A = 8'hED; B = 8'h6B; #100;
A = 8'hED; B = 8'h6C; #100;
A = 8'hED; B = 8'h6D; #100;
A = 8'hED; B = 8'h6E; #100;
A = 8'hED; B = 8'h6F; #100;
A = 8'hED; B = 8'h70; #100;
A = 8'hED; B = 8'h71; #100;
A = 8'hED; B = 8'h72; #100;
A = 8'hED; B = 8'h73; #100;
A = 8'hED; B = 8'h74; #100;
A = 8'hED; B = 8'h75; #100;
A = 8'hED; B = 8'h76; #100;
A = 8'hED; B = 8'h77; #100;
A = 8'hED; B = 8'h78; #100;
A = 8'hED; B = 8'h79; #100;
A = 8'hED; B = 8'h7A; #100;
A = 8'hED; B = 8'h7B; #100;
A = 8'hED; B = 8'h7C; #100;
A = 8'hED; B = 8'h7D; #100;
A = 8'hED; B = 8'h7E; #100;
A = 8'hED; B = 8'h7F; #100;
A = 8'hED; B = 8'h80; #100;
A = 8'hED; B = 8'h81; #100;
A = 8'hED; B = 8'h82; #100;
A = 8'hED; B = 8'h83; #100;
A = 8'hED; B = 8'h84; #100;
A = 8'hED; B = 8'h85; #100;
A = 8'hED; B = 8'h86; #100;
A = 8'hED; B = 8'h87; #100;
A = 8'hED; B = 8'h88; #100;
A = 8'hED; B = 8'h89; #100;
A = 8'hED; B = 8'h8A; #100;
A = 8'hED; B = 8'h8B; #100;
A = 8'hED; B = 8'h8C; #100;
A = 8'hED; B = 8'h8D; #100;
A = 8'hED; B = 8'h8E; #100;
A = 8'hED; B = 8'h8F; #100;
A = 8'hED; B = 8'h90; #100;
A = 8'hED; B = 8'h91; #100;
A = 8'hED; B = 8'h92; #100;
A = 8'hED; B = 8'h93; #100;
A = 8'hED; B = 8'h94; #100;
A = 8'hED; B = 8'h95; #100;
A = 8'hED; B = 8'h96; #100;
A = 8'hED; B = 8'h97; #100;
A = 8'hED; B = 8'h98; #100;
A = 8'hED; B = 8'h99; #100;
A = 8'hED; B = 8'h9A; #100;
A = 8'hED; B = 8'h9B; #100;
A = 8'hED; B = 8'h9C; #100;
A = 8'hED; B = 8'h9D; #100;
A = 8'hED; B = 8'h9E; #100;
A = 8'hED; B = 8'h9F; #100;
A = 8'hED; B = 8'hA0; #100;
A = 8'hED; B = 8'hA1; #100;
A = 8'hED; B = 8'hA2; #100;
A = 8'hED; B = 8'hA3; #100;
A = 8'hED; B = 8'hA4; #100;
A = 8'hED; B = 8'hA5; #100;
A = 8'hED; B = 8'hA6; #100;
A = 8'hED; B = 8'hA7; #100;
A = 8'hED; B = 8'hA8; #100;
A = 8'hED; B = 8'hA9; #100;
A = 8'hED; B = 8'hAA; #100;
A = 8'hED; B = 8'hAB; #100;
A = 8'hED; B = 8'hAC; #100;
A = 8'hED; B = 8'hAD; #100;
A = 8'hED; B = 8'hAE; #100;
A = 8'hED; B = 8'hAF; #100;
A = 8'hED; B = 8'hB0; #100;
A = 8'hED; B = 8'hB1; #100;
A = 8'hED; B = 8'hB2; #100;
A = 8'hED; B = 8'hB3; #100;
A = 8'hED; B = 8'hB4; #100;
A = 8'hED; B = 8'hB5; #100;
A = 8'hED; B = 8'hB6; #100;
A = 8'hED; B = 8'hB7; #100;
A = 8'hED; B = 8'hB8; #100;
A = 8'hED; B = 8'hB9; #100;
A = 8'hED; B = 8'hBA; #100;
A = 8'hED; B = 8'hBB; #100;
A = 8'hED; B = 8'hBC; #100;
A = 8'hED; B = 8'hBD; #100;
A = 8'hED; B = 8'hBE; #100;
A = 8'hED; B = 8'hBF; #100;
A = 8'hED; B = 8'hC0; #100;
A = 8'hED; B = 8'hC1; #100;
A = 8'hED; B = 8'hC2; #100;
A = 8'hED; B = 8'hC3; #100;
A = 8'hED; B = 8'hC4; #100;
A = 8'hED; B = 8'hC5; #100;
A = 8'hED; B = 8'hC6; #100;
A = 8'hED; B = 8'hC7; #100;
A = 8'hED; B = 8'hC8; #100;
A = 8'hED; B = 8'hC9; #100;
A = 8'hED; B = 8'hCA; #100;
A = 8'hED; B = 8'hCB; #100;
A = 8'hED; B = 8'hCC; #100;
A = 8'hED; B = 8'hCD; #100;
A = 8'hED; B = 8'hCE; #100;
A = 8'hED; B = 8'hCF; #100;
A = 8'hED; B = 8'hD0; #100;
A = 8'hED; B = 8'hD1; #100;
A = 8'hED; B = 8'hD2; #100;
A = 8'hED; B = 8'hD3; #100;
A = 8'hED; B = 8'hD4; #100;
A = 8'hED; B = 8'hD5; #100;
A = 8'hED; B = 8'hD6; #100;
A = 8'hED; B = 8'hD7; #100;
A = 8'hED; B = 8'hD8; #100;
A = 8'hED; B = 8'hD9; #100;
A = 8'hED; B = 8'hDA; #100;
A = 8'hED; B = 8'hDB; #100;
A = 8'hED; B = 8'hDC; #100;
A = 8'hED; B = 8'hDD; #100;
A = 8'hED; B = 8'hDE; #100;
A = 8'hED; B = 8'hDF; #100;
A = 8'hED; B = 8'hE0; #100;
A = 8'hED; B = 8'hE1; #100;
A = 8'hED; B = 8'hE2; #100;
A = 8'hED; B = 8'hE3; #100;
A = 8'hED; B = 8'hE4; #100;
A = 8'hED; B = 8'hE5; #100;
A = 8'hED; B = 8'hE6; #100;
A = 8'hED; B = 8'hE7; #100;
A = 8'hED; B = 8'hE8; #100;
A = 8'hED; B = 8'hE9; #100;
A = 8'hED; B = 8'hEA; #100;
A = 8'hED; B = 8'hEB; #100;
A = 8'hED; B = 8'hEC; #100;
A = 8'hED; B = 8'hED; #100;
A = 8'hED; B = 8'hEE; #100;
A = 8'hED; B = 8'hEF; #100;
A = 8'hED; B = 8'hF0; #100;
A = 8'hED; B = 8'hF1; #100;
A = 8'hED; B = 8'hF2; #100;
A = 8'hED; B = 8'hF3; #100;
A = 8'hED; B = 8'hF4; #100;
A = 8'hED; B = 8'hF5; #100;
A = 8'hED; B = 8'hF6; #100;
A = 8'hED; B = 8'hF7; #100;
A = 8'hED; B = 8'hF8; #100;
A = 8'hED; B = 8'hF9; #100;
A = 8'hED; B = 8'hFA; #100;
A = 8'hED; B = 8'hFB; #100;
A = 8'hED; B = 8'hFC; #100;
A = 8'hED; B = 8'hFD; #100;
A = 8'hED; B = 8'hFE; #100;
A = 8'hED; B = 8'hFF; #100;
A = 8'hEE; B = 8'h0; #100;
A = 8'hEE; B = 8'h1; #100;
A = 8'hEE; B = 8'h2; #100;
A = 8'hEE; B = 8'h3; #100;
A = 8'hEE; B = 8'h4; #100;
A = 8'hEE; B = 8'h5; #100;
A = 8'hEE; B = 8'h6; #100;
A = 8'hEE; B = 8'h7; #100;
A = 8'hEE; B = 8'h8; #100;
A = 8'hEE; B = 8'h9; #100;
A = 8'hEE; B = 8'hA; #100;
A = 8'hEE; B = 8'hB; #100;
A = 8'hEE; B = 8'hC; #100;
A = 8'hEE; B = 8'hD; #100;
A = 8'hEE; B = 8'hE; #100;
A = 8'hEE; B = 8'hF; #100;
A = 8'hEE; B = 8'h10; #100;
A = 8'hEE; B = 8'h11; #100;
A = 8'hEE; B = 8'h12; #100;
A = 8'hEE; B = 8'h13; #100;
A = 8'hEE; B = 8'h14; #100;
A = 8'hEE; B = 8'h15; #100;
A = 8'hEE; B = 8'h16; #100;
A = 8'hEE; B = 8'h17; #100;
A = 8'hEE; B = 8'h18; #100;
A = 8'hEE; B = 8'h19; #100;
A = 8'hEE; B = 8'h1A; #100;
A = 8'hEE; B = 8'h1B; #100;
A = 8'hEE; B = 8'h1C; #100;
A = 8'hEE; B = 8'h1D; #100;
A = 8'hEE; B = 8'h1E; #100;
A = 8'hEE; B = 8'h1F; #100;
A = 8'hEE; B = 8'h20; #100;
A = 8'hEE; B = 8'h21; #100;
A = 8'hEE; B = 8'h22; #100;
A = 8'hEE; B = 8'h23; #100;
A = 8'hEE; B = 8'h24; #100;
A = 8'hEE; B = 8'h25; #100;
A = 8'hEE; B = 8'h26; #100;
A = 8'hEE; B = 8'h27; #100;
A = 8'hEE; B = 8'h28; #100;
A = 8'hEE; B = 8'h29; #100;
A = 8'hEE; B = 8'h2A; #100;
A = 8'hEE; B = 8'h2B; #100;
A = 8'hEE; B = 8'h2C; #100;
A = 8'hEE; B = 8'h2D; #100;
A = 8'hEE; B = 8'h2E; #100;
A = 8'hEE; B = 8'h2F; #100;
A = 8'hEE; B = 8'h30; #100;
A = 8'hEE; B = 8'h31; #100;
A = 8'hEE; B = 8'h32; #100;
A = 8'hEE; B = 8'h33; #100;
A = 8'hEE; B = 8'h34; #100;
A = 8'hEE; B = 8'h35; #100;
A = 8'hEE; B = 8'h36; #100;
A = 8'hEE; B = 8'h37; #100;
A = 8'hEE; B = 8'h38; #100;
A = 8'hEE; B = 8'h39; #100;
A = 8'hEE; B = 8'h3A; #100;
A = 8'hEE; B = 8'h3B; #100;
A = 8'hEE; B = 8'h3C; #100;
A = 8'hEE; B = 8'h3D; #100;
A = 8'hEE; B = 8'h3E; #100;
A = 8'hEE; B = 8'h3F; #100;
A = 8'hEE; B = 8'h40; #100;
A = 8'hEE; B = 8'h41; #100;
A = 8'hEE; B = 8'h42; #100;
A = 8'hEE; B = 8'h43; #100;
A = 8'hEE; B = 8'h44; #100;
A = 8'hEE; B = 8'h45; #100;
A = 8'hEE; B = 8'h46; #100;
A = 8'hEE; B = 8'h47; #100;
A = 8'hEE; B = 8'h48; #100;
A = 8'hEE; B = 8'h49; #100;
A = 8'hEE; B = 8'h4A; #100;
A = 8'hEE; B = 8'h4B; #100;
A = 8'hEE; B = 8'h4C; #100;
A = 8'hEE; B = 8'h4D; #100;
A = 8'hEE; B = 8'h4E; #100;
A = 8'hEE; B = 8'h4F; #100;
A = 8'hEE; B = 8'h50; #100;
A = 8'hEE; B = 8'h51; #100;
A = 8'hEE; B = 8'h52; #100;
A = 8'hEE; B = 8'h53; #100;
A = 8'hEE; B = 8'h54; #100;
A = 8'hEE; B = 8'h55; #100;
A = 8'hEE; B = 8'h56; #100;
A = 8'hEE; B = 8'h57; #100;
A = 8'hEE; B = 8'h58; #100;
A = 8'hEE; B = 8'h59; #100;
A = 8'hEE; B = 8'h5A; #100;
A = 8'hEE; B = 8'h5B; #100;
A = 8'hEE; B = 8'h5C; #100;
A = 8'hEE; B = 8'h5D; #100;
A = 8'hEE; B = 8'h5E; #100;
A = 8'hEE; B = 8'h5F; #100;
A = 8'hEE; B = 8'h60; #100;
A = 8'hEE; B = 8'h61; #100;
A = 8'hEE; B = 8'h62; #100;
A = 8'hEE; B = 8'h63; #100;
A = 8'hEE; B = 8'h64; #100;
A = 8'hEE; B = 8'h65; #100;
A = 8'hEE; B = 8'h66; #100;
A = 8'hEE; B = 8'h67; #100;
A = 8'hEE; B = 8'h68; #100;
A = 8'hEE; B = 8'h69; #100;
A = 8'hEE; B = 8'h6A; #100;
A = 8'hEE; B = 8'h6B; #100;
A = 8'hEE; B = 8'h6C; #100;
A = 8'hEE; B = 8'h6D; #100;
A = 8'hEE; B = 8'h6E; #100;
A = 8'hEE; B = 8'h6F; #100;
A = 8'hEE; B = 8'h70; #100;
A = 8'hEE; B = 8'h71; #100;
A = 8'hEE; B = 8'h72; #100;
A = 8'hEE; B = 8'h73; #100;
A = 8'hEE; B = 8'h74; #100;
A = 8'hEE; B = 8'h75; #100;
A = 8'hEE; B = 8'h76; #100;
A = 8'hEE; B = 8'h77; #100;
A = 8'hEE; B = 8'h78; #100;
A = 8'hEE; B = 8'h79; #100;
A = 8'hEE; B = 8'h7A; #100;
A = 8'hEE; B = 8'h7B; #100;
A = 8'hEE; B = 8'h7C; #100;
A = 8'hEE; B = 8'h7D; #100;
A = 8'hEE; B = 8'h7E; #100;
A = 8'hEE; B = 8'h7F; #100;
A = 8'hEE; B = 8'h80; #100;
A = 8'hEE; B = 8'h81; #100;
A = 8'hEE; B = 8'h82; #100;
A = 8'hEE; B = 8'h83; #100;
A = 8'hEE; B = 8'h84; #100;
A = 8'hEE; B = 8'h85; #100;
A = 8'hEE; B = 8'h86; #100;
A = 8'hEE; B = 8'h87; #100;
A = 8'hEE; B = 8'h88; #100;
A = 8'hEE; B = 8'h89; #100;
A = 8'hEE; B = 8'h8A; #100;
A = 8'hEE; B = 8'h8B; #100;
A = 8'hEE; B = 8'h8C; #100;
A = 8'hEE; B = 8'h8D; #100;
A = 8'hEE; B = 8'h8E; #100;
A = 8'hEE; B = 8'h8F; #100;
A = 8'hEE; B = 8'h90; #100;
A = 8'hEE; B = 8'h91; #100;
A = 8'hEE; B = 8'h92; #100;
A = 8'hEE; B = 8'h93; #100;
A = 8'hEE; B = 8'h94; #100;
A = 8'hEE; B = 8'h95; #100;
A = 8'hEE; B = 8'h96; #100;
A = 8'hEE; B = 8'h97; #100;
A = 8'hEE; B = 8'h98; #100;
A = 8'hEE; B = 8'h99; #100;
A = 8'hEE; B = 8'h9A; #100;
A = 8'hEE; B = 8'h9B; #100;
A = 8'hEE; B = 8'h9C; #100;
A = 8'hEE; B = 8'h9D; #100;
A = 8'hEE; B = 8'h9E; #100;
A = 8'hEE; B = 8'h9F; #100;
A = 8'hEE; B = 8'hA0; #100;
A = 8'hEE; B = 8'hA1; #100;
A = 8'hEE; B = 8'hA2; #100;
A = 8'hEE; B = 8'hA3; #100;
A = 8'hEE; B = 8'hA4; #100;
A = 8'hEE; B = 8'hA5; #100;
A = 8'hEE; B = 8'hA6; #100;
A = 8'hEE; B = 8'hA7; #100;
A = 8'hEE; B = 8'hA8; #100;
A = 8'hEE; B = 8'hA9; #100;
A = 8'hEE; B = 8'hAA; #100;
A = 8'hEE; B = 8'hAB; #100;
A = 8'hEE; B = 8'hAC; #100;
A = 8'hEE; B = 8'hAD; #100;
A = 8'hEE; B = 8'hAE; #100;
A = 8'hEE; B = 8'hAF; #100;
A = 8'hEE; B = 8'hB0; #100;
A = 8'hEE; B = 8'hB1; #100;
A = 8'hEE; B = 8'hB2; #100;
A = 8'hEE; B = 8'hB3; #100;
A = 8'hEE; B = 8'hB4; #100;
A = 8'hEE; B = 8'hB5; #100;
A = 8'hEE; B = 8'hB6; #100;
A = 8'hEE; B = 8'hB7; #100;
A = 8'hEE; B = 8'hB8; #100;
A = 8'hEE; B = 8'hB9; #100;
A = 8'hEE; B = 8'hBA; #100;
A = 8'hEE; B = 8'hBB; #100;
A = 8'hEE; B = 8'hBC; #100;
A = 8'hEE; B = 8'hBD; #100;
A = 8'hEE; B = 8'hBE; #100;
A = 8'hEE; B = 8'hBF; #100;
A = 8'hEE; B = 8'hC0; #100;
A = 8'hEE; B = 8'hC1; #100;
A = 8'hEE; B = 8'hC2; #100;
A = 8'hEE; B = 8'hC3; #100;
A = 8'hEE; B = 8'hC4; #100;
A = 8'hEE; B = 8'hC5; #100;
A = 8'hEE; B = 8'hC6; #100;
A = 8'hEE; B = 8'hC7; #100;
A = 8'hEE; B = 8'hC8; #100;
A = 8'hEE; B = 8'hC9; #100;
A = 8'hEE; B = 8'hCA; #100;
A = 8'hEE; B = 8'hCB; #100;
A = 8'hEE; B = 8'hCC; #100;
A = 8'hEE; B = 8'hCD; #100;
A = 8'hEE; B = 8'hCE; #100;
A = 8'hEE; B = 8'hCF; #100;
A = 8'hEE; B = 8'hD0; #100;
A = 8'hEE; B = 8'hD1; #100;
A = 8'hEE; B = 8'hD2; #100;
A = 8'hEE; B = 8'hD3; #100;
A = 8'hEE; B = 8'hD4; #100;
A = 8'hEE; B = 8'hD5; #100;
A = 8'hEE; B = 8'hD6; #100;
A = 8'hEE; B = 8'hD7; #100;
A = 8'hEE; B = 8'hD8; #100;
A = 8'hEE; B = 8'hD9; #100;
A = 8'hEE; B = 8'hDA; #100;
A = 8'hEE; B = 8'hDB; #100;
A = 8'hEE; B = 8'hDC; #100;
A = 8'hEE; B = 8'hDD; #100;
A = 8'hEE; B = 8'hDE; #100;
A = 8'hEE; B = 8'hDF; #100;
A = 8'hEE; B = 8'hE0; #100;
A = 8'hEE; B = 8'hE1; #100;
A = 8'hEE; B = 8'hE2; #100;
A = 8'hEE; B = 8'hE3; #100;
A = 8'hEE; B = 8'hE4; #100;
A = 8'hEE; B = 8'hE5; #100;
A = 8'hEE; B = 8'hE6; #100;
A = 8'hEE; B = 8'hE7; #100;
A = 8'hEE; B = 8'hE8; #100;
A = 8'hEE; B = 8'hE9; #100;
A = 8'hEE; B = 8'hEA; #100;
A = 8'hEE; B = 8'hEB; #100;
A = 8'hEE; B = 8'hEC; #100;
A = 8'hEE; B = 8'hED; #100;
A = 8'hEE; B = 8'hEE; #100;
A = 8'hEE; B = 8'hEF; #100;
A = 8'hEE; B = 8'hF0; #100;
A = 8'hEE; B = 8'hF1; #100;
A = 8'hEE; B = 8'hF2; #100;
A = 8'hEE; B = 8'hF3; #100;
A = 8'hEE; B = 8'hF4; #100;
A = 8'hEE; B = 8'hF5; #100;
A = 8'hEE; B = 8'hF6; #100;
A = 8'hEE; B = 8'hF7; #100;
A = 8'hEE; B = 8'hF8; #100;
A = 8'hEE; B = 8'hF9; #100;
A = 8'hEE; B = 8'hFA; #100;
A = 8'hEE; B = 8'hFB; #100;
A = 8'hEE; B = 8'hFC; #100;
A = 8'hEE; B = 8'hFD; #100;
A = 8'hEE; B = 8'hFE; #100;
A = 8'hEE; B = 8'hFF; #100;
A = 8'hEF; B = 8'h0; #100;
A = 8'hEF; B = 8'h1; #100;
A = 8'hEF; B = 8'h2; #100;
A = 8'hEF; B = 8'h3; #100;
A = 8'hEF; B = 8'h4; #100;
A = 8'hEF; B = 8'h5; #100;
A = 8'hEF; B = 8'h6; #100;
A = 8'hEF; B = 8'h7; #100;
A = 8'hEF; B = 8'h8; #100;
A = 8'hEF; B = 8'h9; #100;
A = 8'hEF; B = 8'hA; #100;
A = 8'hEF; B = 8'hB; #100;
A = 8'hEF; B = 8'hC; #100;
A = 8'hEF; B = 8'hD; #100;
A = 8'hEF; B = 8'hE; #100;
A = 8'hEF; B = 8'hF; #100;
A = 8'hEF; B = 8'h10; #100;
A = 8'hEF; B = 8'h11; #100;
A = 8'hEF; B = 8'h12; #100;
A = 8'hEF; B = 8'h13; #100;
A = 8'hEF; B = 8'h14; #100;
A = 8'hEF; B = 8'h15; #100;
A = 8'hEF; B = 8'h16; #100;
A = 8'hEF; B = 8'h17; #100;
A = 8'hEF; B = 8'h18; #100;
A = 8'hEF; B = 8'h19; #100;
A = 8'hEF; B = 8'h1A; #100;
A = 8'hEF; B = 8'h1B; #100;
A = 8'hEF; B = 8'h1C; #100;
A = 8'hEF; B = 8'h1D; #100;
A = 8'hEF; B = 8'h1E; #100;
A = 8'hEF; B = 8'h1F; #100;
A = 8'hEF; B = 8'h20; #100;
A = 8'hEF; B = 8'h21; #100;
A = 8'hEF; B = 8'h22; #100;
A = 8'hEF; B = 8'h23; #100;
A = 8'hEF; B = 8'h24; #100;
A = 8'hEF; B = 8'h25; #100;
A = 8'hEF; B = 8'h26; #100;
A = 8'hEF; B = 8'h27; #100;
A = 8'hEF; B = 8'h28; #100;
A = 8'hEF; B = 8'h29; #100;
A = 8'hEF; B = 8'h2A; #100;
A = 8'hEF; B = 8'h2B; #100;
A = 8'hEF; B = 8'h2C; #100;
A = 8'hEF; B = 8'h2D; #100;
A = 8'hEF; B = 8'h2E; #100;
A = 8'hEF; B = 8'h2F; #100;
A = 8'hEF; B = 8'h30; #100;
A = 8'hEF; B = 8'h31; #100;
A = 8'hEF; B = 8'h32; #100;
A = 8'hEF; B = 8'h33; #100;
A = 8'hEF; B = 8'h34; #100;
A = 8'hEF; B = 8'h35; #100;
A = 8'hEF; B = 8'h36; #100;
A = 8'hEF; B = 8'h37; #100;
A = 8'hEF; B = 8'h38; #100;
A = 8'hEF; B = 8'h39; #100;
A = 8'hEF; B = 8'h3A; #100;
A = 8'hEF; B = 8'h3B; #100;
A = 8'hEF; B = 8'h3C; #100;
A = 8'hEF; B = 8'h3D; #100;
A = 8'hEF; B = 8'h3E; #100;
A = 8'hEF; B = 8'h3F; #100;
A = 8'hEF; B = 8'h40; #100;
A = 8'hEF; B = 8'h41; #100;
A = 8'hEF; B = 8'h42; #100;
A = 8'hEF; B = 8'h43; #100;
A = 8'hEF; B = 8'h44; #100;
A = 8'hEF; B = 8'h45; #100;
A = 8'hEF; B = 8'h46; #100;
A = 8'hEF; B = 8'h47; #100;
A = 8'hEF; B = 8'h48; #100;
A = 8'hEF; B = 8'h49; #100;
A = 8'hEF; B = 8'h4A; #100;
A = 8'hEF; B = 8'h4B; #100;
A = 8'hEF; B = 8'h4C; #100;
A = 8'hEF; B = 8'h4D; #100;
A = 8'hEF; B = 8'h4E; #100;
A = 8'hEF; B = 8'h4F; #100;
A = 8'hEF; B = 8'h50; #100;
A = 8'hEF; B = 8'h51; #100;
A = 8'hEF; B = 8'h52; #100;
A = 8'hEF; B = 8'h53; #100;
A = 8'hEF; B = 8'h54; #100;
A = 8'hEF; B = 8'h55; #100;
A = 8'hEF; B = 8'h56; #100;
A = 8'hEF; B = 8'h57; #100;
A = 8'hEF; B = 8'h58; #100;
A = 8'hEF; B = 8'h59; #100;
A = 8'hEF; B = 8'h5A; #100;
A = 8'hEF; B = 8'h5B; #100;
A = 8'hEF; B = 8'h5C; #100;
A = 8'hEF; B = 8'h5D; #100;
A = 8'hEF; B = 8'h5E; #100;
A = 8'hEF; B = 8'h5F; #100;
A = 8'hEF; B = 8'h60; #100;
A = 8'hEF; B = 8'h61; #100;
A = 8'hEF; B = 8'h62; #100;
A = 8'hEF; B = 8'h63; #100;
A = 8'hEF; B = 8'h64; #100;
A = 8'hEF; B = 8'h65; #100;
A = 8'hEF; B = 8'h66; #100;
A = 8'hEF; B = 8'h67; #100;
A = 8'hEF; B = 8'h68; #100;
A = 8'hEF; B = 8'h69; #100;
A = 8'hEF; B = 8'h6A; #100;
A = 8'hEF; B = 8'h6B; #100;
A = 8'hEF; B = 8'h6C; #100;
A = 8'hEF; B = 8'h6D; #100;
A = 8'hEF; B = 8'h6E; #100;
A = 8'hEF; B = 8'h6F; #100;
A = 8'hEF; B = 8'h70; #100;
A = 8'hEF; B = 8'h71; #100;
A = 8'hEF; B = 8'h72; #100;
A = 8'hEF; B = 8'h73; #100;
A = 8'hEF; B = 8'h74; #100;
A = 8'hEF; B = 8'h75; #100;
A = 8'hEF; B = 8'h76; #100;
A = 8'hEF; B = 8'h77; #100;
A = 8'hEF; B = 8'h78; #100;
A = 8'hEF; B = 8'h79; #100;
A = 8'hEF; B = 8'h7A; #100;
A = 8'hEF; B = 8'h7B; #100;
A = 8'hEF; B = 8'h7C; #100;
A = 8'hEF; B = 8'h7D; #100;
A = 8'hEF; B = 8'h7E; #100;
A = 8'hEF; B = 8'h7F; #100;
A = 8'hEF; B = 8'h80; #100;
A = 8'hEF; B = 8'h81; #100;
A = 8'hEF; B = 8'h82; #100;
A = 8'hEF; B = 8'h83; #100;
A = 8'hEF; B = 8'h84; #100;
A = 8'hEF; B = 8'h85; #100;
A = 8'hEF; B = 8'h86; #100;
A = 8'hEF; B = 8'h87; #100;
A = 8'hEF; B = 8'h88; #100;
A = 8'hEF; B = 8'h89; #100;
A = 8'hEF; B = 8'h8A; #100;
A = 8'hEF; B = 8'h8B; #100;
A = 8'hEF; B = 8'h8C; #100;
A = 8'hEF; B = 8'h8D; #100;
A = 8'hEF; B = 8'h8E; #100;
A = 8'hEF; B = 8'h8F; #100;
A = 8'hEF; B = 8'h90; #100;
A = 8'hEF; B = 8'h91; #100;
A = 8'hEF; B = 8'h92; #100;
A = 8'hEF; B = 8'h93; #100;
A = 8'hEF; B = 8'h94; #100;
A = 8'hEF; B = 8'h95; #100;
A = 8'hEF; B = 8'h96; #100;
A = 8'hEF; B = 8'h97; #100;
A = 8'hEF; B = 8'h98; #100;
A = 8'hEF; B = 8'h99; #100;
A = 8'hEF; B = 8'h9A; #100;
A = 8'hEF; B = 8'h9B; #100;
A = 8'hEF; B = 8'h9C; #100;
A = 8'hEF; B = 8'h9D; #100;
A = 8'hEF; B = 8'h9E; #100;
A = 8'hEF; B = 8'h9F; #100;
A = 8'hEF; B = 8'hA0; #100;
A = 8'hEF; B = 8'hA1; #100;
A = 8'hEF; B = 8'hA2; #100;
A = 8'hEF; B = 8'hA3; #100;
A = 8'hEF; B = 8'hA4; #100;
A = 8'hEF; B = 8'hA5; #100;
A = 8'hEF; B = 8'hA6; #100;
A = 8'hEF; B = 8'hA7; #100;
A = 8'hEF; B = 8'hA8; #100;
A = 8'hEF; B = 8'hA9; #100;
A = 8'hEF; B = 8'hAA; #100;
A = 8'hEF; B = 8'hAB; #100;
A = 8'hEF; B = 8'hAC; #100;
A = 8'hEF; B = 8'hAD; #100;
A = 8'hEF; B = 8'hAE; #100;
A = 8'hEF; B = 8'hAF; #100;
A = 8'hEF; B = 8'hB0; #100;
A = 8'hEF; B = 8'hB1; #100;
A = 8'hEF; B = 8'hB2; #100;
A = 8'hEF; B = 8'hB3; #100;
A = 8'hEF; B = 8'hB4; #100;
A = 8'hEF; B = 8'hB5; #100;
A = 8'hEF; B = 8'hB6; #100;
A = 8'hEF; B = 8'hB7; #100;
A = 8'hEF; B = 8'hB8; #100;
A = 8'hEF; B = 8'hB9; #100;
A = 8'hEF; B = 8'hBA; #100;
A = 8'hEF; B = 8'hBB; #100;
A = 8'hEF; B = 8'hBC; #100;
A = 8'hEF; B = 8'hBD; #100;
A = 8'hEF; B = 8'hBE; #100;
A = 8'hEF; B = 8'hBF; #100;
A = 8'hEF; B = 8'hC0; #100;
A = 8'hEF; B = 8'hC1; #100;
A = 8'hEF; B = 8'hC2; #100;
A = 8'hEF; B = 8'hC3; #100;
A = 8'hEF; B = 8'hC4; #100;
A = 8'hEF; B = 8'hC5; #100;
A = 8'hEF; B = 8'hC6; #100;
A = 8'hEF; B = 8'hC7; #100;
A = 8'hEF; B = 8'hC8; #100;
A = 8'hEF; B = 8'hC9; #100;
A = 8'hEF; B = 8'hCA; #100;
A = 8'hEF; B = 8'hCB; #100;
A = 8'hEF; B = 8'hCC; #100;
A = 8'hEF; B = 8'hCD; #100;
A = 8'hEF; B = 8'hCE; #100;
A = 8'hEF; B = 8'hCF; #100;
A = 8'hEF; B = 8'hD0; #100;
A = 8'hEF; B = 8'hD1; #100;
A = 8'hEF; B = 8'hD2; #100;
A = 8'hEF; B = 8'hD3; #100;
A = 8'hEF; B = 8'hD4; #100;
A = 8'hEF; B = 8'hD5; #100;
A = 8'hEF; B = 8'hD6; #100;
A = 8'hEF; B = 8'hD7; #100;
A = 8'hEF; B = 8'hD8; #100;
A = 8'hEF; B = 8'hD9; #100;
A = 8'hEF; B = 8'hDA; #100;
A = 8'hEF; B = 8'hDB; #100;
A = 8'hEF; B = 8'hDC; #100;
A = 8'hEF; B = 8'hDD; #100;
A = 8'hEF; B = 8'hDE; #100;
A = 8'hEF; B = 8'hDF; #100;
A = 8'hEF; B = 8'hE0; #100;
A = 8'hEF; B = 8'hE1; #100;
A = 8'hEF; B = 8'hE2; #100;
A = 8'hEF; B = 8'hE3; #100;
A = 8'hEF; B = 8'hE4; #100;
A = 8'hEF; B = 8'hE5; #100;
A = 8'hEF; B = 8'hE6; #100;
A = 8'hEF; B = 8'hE7; #100;
A = 8'hEF; B = 8'hE8; #100;
A = 8'hEF; B = 8'hE9; #100;
A = 8'hEF; B = 8'hEA; #100;
A = 8'hEF; B = 8'hEB; #100;
A = 8'hEF; B = 8'hEC; #100;
A = 8'hEF; B = 8'hED; #100;
A = 8'hEF; B = 8'hEE; #100;
A = 8'hEF; B = 8'hEF; #100;
A = 8'hEF; B = 8'hF0; #100;
A = 8'hEF; B = 8'hF1; #100;
A = 8'hEF; B = 8'hF2; #100;
A = 8'hEF; B = 8'hF3; #100;
A = 8'hEF; B = 8'hF4; #100;
A = 8'hEF; B = 8'hF5; #100;
A = 8'hEF; B = 8'hF6; #100;
A = 8'hEF; B = 8'hF7; #100;
A = 8'hEF; B = 8'hF8; #100;
A = 8'hEF; B = 8'hF9; #100;
A = 8'hEF; B = 8'hFA; #100;
A = 8'hEF; B = 8'hFB; #100;
A = 8'hEF; B = 8'hFC; #100;
A = 8'hEF; B = 8'hFD; #100;
A = 8'hEF; B = 8'hFE; #100;
A = 8'hEF; B = 8'hFF; #100;
A = 8'hF0; B = 8'h0; #100;
A = 8'hF0; B = 8'h1; #100;
A = 8'hF0; B = 8'h2; #100;
A = 8'hF0; B = 8'h3; #100;
A = 8'hF0; B = 8'h4; #100;
A = 8'hF0; B = 8'h5; #100;
A = 8'hF0; B = 8'h6; #100;
A = 8'hF0; B = 8'h7; #100;
A = 8'hF0; B = 8'h8; #100;
A = 8'hF0; B = 8'h9; #100;
A = 8'hF0; B = 8'hA; #100;
A = 8'hF0; B = 8'hB; #100;
A = 8'hF0; B = 8'hC; #100;
A = 8'hF0; B = 8'hD; #100;
A = 8'hF0; B = 8'hE; #100;
A = 8'hF0; B = 8'hF; #100;
A = 8'hF0; B = 8'h10; #100;
A = 8'hF0; B = 8'h11; #100;
A = 8'hF0; B = 8'h12; #100;
A = 8'hF0; B = 8'h13; #100;
A = 8'hF0; B = 8'h14; #100;
A = 8'hF0; B = 8'h15; #100;
A = 8'hF0; B = 8'h16; #100;
A = 8'hF0; B = 8'h17; #100;
A = 8'hF0; B = 8'h18; #100;
A = 8'hF0; B = 8'h19; #100;
A = 8'hF0; B = 8'h1A; #100;
A = 8'hF0; B = 8'h1B; #100;
A = 8'hF0; B = 8'h1C; #100;
A = 8'hF0; B = 8'h1D; #100;
A = 8'hF0; B = 8'h1E; #100;
A = 8'hF0; B = 8'h1F; #100;
A = 8'hF0; B = 8'h20; #100;
A = 8'hF0; B = 8'h21; #100;
A = 8'hF0; B = 8'h22; #100;
A = 8'hF0; B = 8'h23; #100;
A = 8'hF0; B = 8'h24; #100;
A = 8'hF0; B = 8'h25; #100;
A = 8'hF0; B = 8'h26; #100;
A = 8'hF0; B = 8'h27; #100;
A = 8'hF0; B = 8'h28; #100;
A = 8'hF0; B = 8'h29; #100;
A = 8'hF0; B = 8'h2A; #100;
A = 8'hF0; B = 8'h2B; #100;
A = 8'hF0; B = 8'h2C; #100;
A = 8'hF0; B = 8'h2D; #100;
A = 8'hF0; B = 8'h2E; #100;
A = 8'hF0; B = 8'h2F; #100;
A = 8'hF0; B = 8'h30; #100;
A = 8'hF0; B = 8'h31; #100;
A = 8'hF0; B = 8'h32; #100;
A = 8'hF0; B = 8'h33; #100;
A = 8'hF0; B = 8'h34; #100;
A = 8'hF0; B = 8'h35; #100;
A = 8'hF0; B = 8'h36; #100;
A = 8'hF0; B = 8'h37; #100;
A = 8'hF0; B = 8'h38; #100;
A = 8'hF0; B = 8'h39; #100;
A = 8'hF0; B = 8'h3A; #100;
A = 8'hF0; B = 8'h3B; #100;
A = 8'hF0; B = 8'h3C; #100;
A = 8'hF0; B = 8'h3D; #100;
A = 8'hF0; B = 8'h3E; #100;
A = 8'hF0; B = 8'h3F; #100;
A = 8'hF0; B = 8'h40; #100;
A = 8'hF0; B = 8'h41; #100;
A = 8'hF0; B = 8'h42; #100;
A = 8'hF0; B = 8'h43; #100;
A = 8'hF0; B = 8'h44; #100;
A = 8'hF0; B = 8'h45; #100;
A = 8'hF0; B = 8'h46; #100;
A = 8'hF0; B = 8'h47; #100;
A = 8'hF0; B = 8'h48; #100;
A = 8'hF0; B = 8'h49; #100;
A = 8'hF0; B = 8'h4A; #100;
A = 8'hF0; B = 8'h4B; #100;
A = 8'hF0; B = 8'h4C; #100;
A = 8'hF0; B = 8'h4D; #100;
A = 8'hF0; B = 8'h4E; #100;
A = 8'hF0; B = 8'h4F; #100;
A = 8'hF0; B = 8'h50; #100;
A = 8'hF0; B = 8'h51; #100;
A = 8'hF0; B = 8'h52; #100;
A = 8'hF0; B = 8'h53; #100;
A = 8'hF0; B = 8'h54; #100;
A = 8'hF0; B = 8'h55; #100;
A = 8'hF0; B = 8'h56; #100;
A = 8'hF0; B = 8'h57; #100;
A = 8'hF0; B = 8'h58; #100;
A = 8'hF0; B = 8'h59; #100;
A = 8'hF0; B = 8'h5A; #100;
A = 8'hF0; B = 8'h5B; #100;
A = 8'hF0; B = 8'h5C; #100;
A = 8'hF0; B = 8'h5D; #100;
A = 8'hF0; B = 8'h5E; #100;
A = 8'hF0; B = 8'h5F; #100;
A = 8'hF0; B = 8'h60; #100;
A = 8'hF0; B = 8'h61; #100;
A = 8'hF0; B = 8'h62; #100;
A = 8'hF0; B = 8'h63; #100;
A = 8'hF0; B = 8'h64; #100;
A = 8'hF0; B = 8'h65; #100;
A = 8'hF0; B = 8'h66; #100;
A = 8'hF0; B = 8'h67; #100;
A = 8'hF0; B = 8'h68; #100;
A = 8'hF0; B = 8'h69; #100;
A = 8'hF0; B = 8'h6A; #100;
A = 8'hF0; B = 8'h6B; #100;
A = 8'hF0; B = 8'h6C; #100;
A = 8'hF0; B = 8'h6D; #100;
A = 8'hF0; B = 8'h6E; #100;
A = 8'hF0; B = 8'h6F; #100;
A = 8'hF0; B = 8'h70; #100;
A = 8'hF0; B = 8'h71; #100;
A = 8'hF0; B = 8'h72; #100;
A = 8'hF0; B = 8'h73; #100;
A = 8'hF0; B = 8'h74; #100;
A = 8'hF0; B = 8'h75; #100;
A = 8'hF0; B = 8'h76; #100;
A = 8'hF0; B = 8'h77; #100;
A = 8'hF0; B = 8'h78; #100;
A = 8'hF0; B = 8'h79; #100;
A = 8'hF0; B = 8'h7A; #100;
A = 8'hF0; B = 8'h7B; #100;
A = 8'hF0; B = 8'h7C; #100;
A = 8'hF0; B = 8'h7D; #100;
A = 8'hF0; B = 8'h7E; #100;
A = 8'hF0; B = 8'h7F; #100;
A = 8'hF0; B = 8'h80; #100;
A = 8'hF0; B = 8'h81; #100;
A = 8'hF0; B = 8'h82; #100;
A = 8'hF0; B = 8'h83; #100;
A = 8'hF0; B = 8'h84; #100;
A = 8'hF0; B = 8'h85; #100;
A = 8'hF0; B = 8'h86; #100;
A = 8'hF0; B = 8'h87; #100;
A = 8'hF0; B = 8'h88; #100;
A = 8'hF0; B = 8'h89; #100;
A = 8'hF0; B = 8'h8A; #100;
A = 8'hF0; B = 8'h8B; #100;
A = 8'hF0; B = 8'h8C; #100;
A = 8'hF0; B = 8'h8D; #100;
A = 8'hF0; B = 8'h8E; #100;
A = 8'hF0; B = 8'h8F; #100;
A = 8'hF0; B = 8'h90; #100;
A = 8'hF0; B = 8'h91; #100;
A = 8'hF0; B = 8'h92; #100;
A = 8'hF0; B = 8'h93; #100;
A = 8'hF0; B = 8'h94; #100;
A = 8'hF0; B = 8'h95; #100;
A = 8'hF0; B = 8'h96; #100;
A = 8'hF0; B = 8'h97; #100;
A = 8'hF0; B = 8'h98; #100;
A = 8'hF0; B = 8'h99; #100;
A = 8'hF0; B = 8'h9A; #100;
A = 8'hF0; B = 8'h9B; #100;
A = 8'hF0; B = 8'h9C; #100;
A = 8'hF0; B = 8'h9D; #100;
A = 8'hF0; B = 8'h9E; #100;
A = 8'hF0; B = 8'h9F; #100;
A = 8'hF0; B = 8'hA0; #100;
A = 8'hF0; B = 8'hA1; #100;
A = 8'hF0; B = 8'hA2; #100;
A = 8'hF0; B = 8'hA3; #100;
A = 8'hF0; B = 8'hA4; #100;
A = 8'hF0; B = 8'hA5; #100;
A = 8'hF0; B = 8'hA6; #100;
A = 8'hF0; B = 8'hA7; #100;
A = 8'hF0; B = 8'hA8; #100;
A = 8'hF0; B = 8'hA9; #100;
A = 8'hF0; B = 8'hAA; #100;
A = 8'hF0; B = 8'hAB; #100;
A = 8'hF0; B = 8'hAC; #100;
A = 8'hF0; B = 8'hAD; #100;
A = 8'hF0; B = 8'hAE; #100;
A = 8'hF0; B = 8'hAF; #100;
A = 8'hF0; B = 8'hB0; #100;
A = 8'hF0; B = 8'hB1; #100;
A = 8'hF0; B = 8'hB2; #100;
A = 8'hF0; B = 8'hB3; #100;
A = 8'hF0; B = 8'hB4; #100;
A = 8'hF0; B = 8'hB5; #100;
A = 8'hF0; B = 8'hB6; #100;
A = 8'hF0; B = 8'hB7; #100;
A = 8'hF0; B = 8'hB8; #100;
A = 8'hF0; B = 8'hB9; #100;
A = 8'hF0; B = 8'hBA; #100;
A = 8'hF0; B = 8'hBB; #100;
A = 8'hF0; B = 8'hBC; #100;
A = 8'hF0; B = 8'hBD; #100;
A = 8'hF0; B = 8'hBE; #100;
A = 8'hF0; B = 8'hBF; #100;
A = 8'hF0; B = 8'hC0; #100;
A = 8'hF0; B = 8'hC1; #100;
A = 8'hF0; B = 8'hC2; #100;
A = 8'hF0; B = 8'hC3; #100;
A = 8'hF0; B = 8'hC4; #100;
A = 8'hF0; B = 8'hC5; #100;
A = 8'hF0; B = 8'hC6; #100;
A = 8'hF0; B = 8'hC7; #100;
A = 8'hF0; B = 8'hC8; #100;
A = 8'hF0; B = 8'hC9; #100;
A = 8'hF0; B = 8'hCA; #100;
A = 8'hF0; B = 8'hCB; #100;
A = 8'hF0; B = 8'hCC; #100;
A = 8'hF0; B = 8'hCD; #100;
A = 8'hF0; B = 8'hCE; #100;
A = 8'hF0; B = 8'hCF; #100;
A = 8'hF0; B = 8'hD0; #100;
A = 8'hF0; B = 8'hD1; #100;
A = 8'hF0; B = 8'hD2; #100;
A = 8'hF0; B = 8'hD3; #100;
A = 8'hF0; B = 8'hD4; #100;
A = 8'hF0; B = 8'hD5; #100;
A = 8'hF0; B = 8'hD6; #100;
A = 8'hF0; B = 8'hD7; #100;
A = 8'hF0; B = 8'hD8; #100;
A = 8'hF0; B = 8'hD9; #100;
A = 8'hF0; B = 8'hDA; #100;
A = 8'hF0; B = 8'hDB; #100;
A = 8'hF0; B = 8'hDC; #100;
A = 8'hF0; B = 8'hDD; #100;
A = 8'hF0; B = 8'hDE; #100;
A = 8'hF0; B = 8'hDF; #100;
A = 8'hF0; B = 8'hE0; #100;
A = 8'hF0; B = 8'hE1; #100;
A = 8'hF0; B = 8'hE2; #100;
A = 8'hF0; B = 8'hE3; #100;
A = 8'hF0; B = 8'hE4; #100;
A = 8'hF0; B = 8'hE5; #100;
A = 8'hF0; B = 8'hE6; #100;
A = 8'hF0; B = 8'hE7; #100;
A = 8'hF0; B = 8'hE8; #100;
A = 8'hF0; B = 8'hE9; #100;
A = 8'hF0; B = 8'hEA; #100;
A = 8'hF0; B = 8'hEB; #100;
A = 8'hF0; B = 8'hEC; #100;
A = 8'hF0; B = 8'hED; #100;
A = 8'hF0; B = 8'hEE; #100;
A = 8'hF0; B = 8'hEF; #100;
A = 8'hF0; B = 8'hF0; #100;
A = 8'hF0; B = 8'hF1; #100;
A = 8'hF0; B = 8'hF2; #100;
A = 8'hF0; B = 8'hF3; #100;
A = 8'hF0; B = 8'hF4; #100;
A = 8'hF0; B = 8'hF5; #100;
A = 8'hF0; B = 8'hF6; #100;
A = 8'hF0; B = 8'hF7; #100;
A = 8'hF0; B = 8'hF8; #100;
A = 8'hF0; B = 8'hF9; #100;
A = 8'hF0; B = 8'hFA; #100;
A = 8'hF0; B = 8'hFB; #100;
A = 8'hF0; B = 8'hFC; #100;
A = 8'hF0; B = 8'hFD; #100;
A = 8'hF0; B = 8'hFE; #100;
A = 8'hF0; B = 8'hFF; #100;
A = 8'hF1; B = 8'h0; #100;
A = 8'hF1; B = 8'h1; #100;
A = 8'hF1; B = 8'h2; #100;
A = 8'hF1; B = 8'h3; #100;
A = 8'hF1; B = 8'h4; #100;
A = 8'hF1; B = 8'h5; #100;
A = 8'hF1; B = 8'h6; #100;
A = 8'hF1; B = 8'h7; #100;
A = 8'hF1; B = 8'h8; #100;
A = 8'hF1; B = 8'h9; #100;
A = 8'hF1; B = 8'hA; #100;
A = 8'hF1; B = 8'hB; #100;
A = 8'hF1; B = 8'hC; #100;
A = 8'hF1; B = 8'hD; #100;
A = 8'hF1; B = 8'hE; #100;
A = 8'hF1; B = 8'hF; #100;
A = 8'hF1; B = 8'h10; #100;
A = 8'hF1; B = 8'h11; #100;
A = 8'hF1; B = 8'h12; #100;
A = 8'hF1; B = 8'h13; #100;
A = 8'hF1; B = 8'h14; #100;
A = 8'hF1; B = 8'h15; #100;
A = 8'hF1; B = 8'h16; #100;
A = 8'hF1; B = 8'h17; #100;
A = 8'hF1; B = 8'h18; #100;
A = 8'hF1; B = 8'h19; #100;
A = 8'hF1; B = 8'h1A; #100;
A = 8'hF1; B = 8'h1B; #100;
A = 8'hF1; B = 8'h1C; #100;
A = 8'hF1; B = 8'h1D; #100;
A = 8'hF1; B = 8'h1E; #100;
A = 8'hF1; B = 8'h1F; #100;
A = 8'hF1; B = 8'h20; #100;
A = 8'hF1; B = 8'h21; #100;
A = 8'hF1; B = 8'h22; #100;
A = 8'hF1; B = 8'h23; #100;
A = 8'hF1; B = 8'h24; #100;
A = 8'hF1; B = 8'h25; #100;
A = 8'hF1; B = 8'h26; #100;
A = 8'hF1; B = 8'h27; #100;
A = 8'hF1; B = 8'h28; #100;
A = 8'hF1; B = 8'h29; #100;
A = 8'hF1; B = 8'h2A; #100;
A = 8'hF1; B = 8'h2B; #100;
A = 8'hF1; B = 8'h2C; #100;
A = 8'hF1; B = 8'h2D; #100;
A = 8'hF1; B = 8'h2E; #100;
A = 8'hF1; B = 8'h2F; #100;
A = 8'hF1; B = 8'h30; #100;
A = 8'hF1; B = 8'h31; #100;
A = 8'hF1; B = 8'h32; #100;
A = 8'hF1; B = 8'h33; #100;
A = 8'hF1; B = 8'h34; #100;
A = 8'hF1; B = 8'h35; #100;
A = 8'hF1; B = 8'h36; #100;
A = 8'hF1; B = 8'h37; #100;
A = 8'hF1; B = 8'h38; #100;
A = 8'hF1; B = 8'h39; #100;
A = 8'hF1; B = 8'h3A; #100;
A = 8'hF1; B = 8'h3B; #100;
A = 8'hF1; B = 8'h3C; #100;
A = 8'hF1; B = 8'h3D; #100;
A = 8'hF1; B = 8'h3E; #100;
A = 8'hF1; B = 8'h3F; #100;
A = 8'hF1; B = 8'h40; #100;
A = 8'hF1; B = 8'h41; #100;
A = 8'hF1; B = 8'h42; #100;
A = 8'hF1; B = 8'h43; #100;
A = 8'hF1; B = 8'h44; #100;
A = 8'hF1; B = 8'h45; #100;
A = 8'hF1; B = 8'h46; #100;
A = 8'hF1; B = 8'h47; #100;
A = 8'hF1; B = 8'h48; #100;
A = 8'hF1; B = 8'h49; #100;
A = 8'hF1; B = 8'h4A; #100;
A = 8'hF1; B = 8'h4B; #100;
A = 8'hF1; B = 8'h4C; #100;
A = 8'hF1; B = 8'h4D; #100;
A = 8'hF1; B = 8'h4E; #100;
A = 8'hF1; B = 8'h4F; #100;
A = 8'hF1; B = 8'h50; #100;
A = 8'hF1; B = 8'h51; #100;
A = 8'hF1; B = 8'h52; #100;
A = 8'hF1; B = 8'h53; #100;
A = 8'hF1; B = 8'h54; #100;
A = 8'hF1; B = 8'h55; #100;
A = 8'hF1; B = 8'h56; #100;
A = 8'hF1; B = 8'h57; #100;
A = 8'hF1; B = 8'h58; #100;
A = 8'hF1; B = 8'h59; #100;
A = 8'hF1; B = 8'h5A; #100;
A = 8'hF1; B = 8'h5B; #100;
A = 8'hF1; B = 8'h5C; #100;
A = 8'hF1; B = 8'h5D; #100;
A = 8'hF1; B = 8'h5E; #100;
A = 8'hF1; B = 8'h5F; #100;
A = 8'hF1; B = 8'h60; #100;
A = 8'hF1; B = 8'h61; #100;
A = 8'hF1; B = 8'h62; #100;
A = 8'hF1; B = 8'h63; #100;
A = 8'hF1; B = 8'h64; #100;
A = 8'hF1; B = 8'h65; #100;
A = 8'hF1; B = 8'h66; #100;
A = 8'hF1; B = 8'h67; #100;
A = 8'hF1; B = 8'h68; #100;
A = 8'hF1; B = 8'h69; #100;
A = 8'hF1; B = 8'h6A; #100;
A = 8'hF1; B = 8'h6B; #100;
A = 8'hF1; B = 8'h6C; #100;
A = 8'hF1; B = 8'h6D; #100;
A = 8'hF1; B = 8'h6E; #100;
A = 8'hF1; B = 8'h6F; #100;
A = 8'hF1; B = 8'h70; #100;
A = 8'hF1; B = 8'h71; #100;
A = 8'hF1; B = 8'h72; #100;
A = 8'hF1; B = 8'h73; #100;
A = 8'hF1; B = 8'h74; #100;
A = 8'hF1; B = 8'h75; #100;
A = 8'hF1; B = 8'h76; #100;
A = 8'hF1; B = 8'h77; #100;
A = 8'hF1; B = 8'h78; #100;
A = 8'hF1; B = 8'h79; #100;
A = 8'hF1; B = 8'h7A; #100;
A = 8'hF1; B = 8'h7B; #100;
A = 8'hF1; B = 8'h7C; #100;
A = 8'hF1; B = 8'h7D; #100;
A = 8'hF1; B = 8'h7E; #100;
A = 8'hF1; B = 8'h7F; #100;
A = 8'hF1; B = 8'h80; #100;
A = 8'hF1; B = 8'h81; #100;
A = 8'hF1; B = 8'h82; #100;
A = 8'hF1; B = 8'h83; #100;
A = 8'hF1; B = 8'h84; #100;
A = 8'hF1; B = 8'h85; #100;
A = 8'hF1; B = 8'h86; #100;
A = 8'hF1; B = 8'h87; #100;
A = 8'hF1; B = 8'h88; #100;
A = 8'hF1; B = 8'h89; #100;
A = 8'hF1; B = 8'h8A; #100;
A = 8'hF1; B = 8'h8B; #100;
A = 8'hF1; B = 8'h8C; #100;
A = 8'hF1; B = 8'h8D; #100;
A = 8'hF1; B = 8'h8E; #100;
A = 8'hF1; B = 8'h8F; #100;
A = 8'hF1; B = 8'h90; #100;
A = 8'hF1; B = 8'h91; #100;
A = 8'hF1; B = 8'h92; #100;
A = 8'hF1; B = 8'h93; #100;
A = 8'hF1; B = 8'h94; #100;
A = 8'hF1; B = 8'h95; #100;
A = 8'hF1; B = 8'h96; #100;
A = 8'hF1; B = 8'h97; #100;
A = 8'hF1; B = 8'h98; #100;
A = 8'hF1; B = 8'h99; #100;
A = 8'hF1; B = 8'h9A; #100;
A = 8'hF1; B = 8'h9B; #100;
A = 8'hF1; B = 8'h9C; #100;
A = 8'hF1; B = 8'h9D; #100;
A = 8'hF1; B = 8'h9E; #100;
A = 8'hF1; B = 8'h9F; #100;
A = 8'hF1; B = 8'hA0; #100;
A = 8'hF1; B = 8'hA1; #100;
A = 8'hF1; B = 8'hA2; #100;
A = 8'hF1; B = 8'hA3; #100;
A = 8'hF1; B = 8'hA4; #100;
A = 8'hF1; B = 8'hA5; #100;
A = 8'hF1; B = 8'hA6; #100;
A = 8'hF1; B = 8'hA7; #100;
A = 8'hF1; B = 8'hA8; #100;
A = 8'hF1; B = 8'hA9; #100;
A = 8'hF1; B = 8'hAA; #100;
A = 8'hF1; B = 8'hAB; #100;
A = 8'hF1; B = 8'hAC; #100;
A = 8'hF1; B = 8'hAD; #100;
A = 8'hF1; B = 8'hAE; #100;
A = 8'hF1; B = 8'hAF; #100;
A = 8'hF1; B = 8'hB0; #100;
A = 8'hF1; B = 8'hB1; #100;
A = 8'hF1; B = 8'hB2; #100;
A = 8'hF1; B = 8'hB3; #100;
A = 8'hF1; B = 8'hB4; #100;
A = 8'hF1; B = 8'hB5; #100;
A = 8'hF1; B = 8'hB6; #100;
A = 8'hF1; B = 8'hB7; #100;
A = 8'hF1; B = 8'hB8; #100;
A = 8'hF1; B = 8'hB9; #100;
A = 8'hF1; B = 8'hBA; #100;
A = 8'hF1; B = 8'hBB; #100;
A = 8'hF1; B = 8'hBC; #100;
A = 8'hF1; B = 8'hBD; #100;
A = 8'hF1; B = 8'hBE; #100;
A = 8'hF1; B = 8'hBF; #100;
A = 8'hF1; B = 8'hC0; #100;
A = 8'hF1; B = 8'hC1; #100;
A = 8'hF1; B = 8'hC2; #100;
A = 8'hF1; B = 8'hC3; #100;
A = 8'hF1; B = 8'hC4; #100;
A = 8'hF1; B = 8'hC5; #100;
A = 8'hF1; B = 8'hC6; #100;
A = 8'hF1; B = 8'hC7; #100;
A = 8'hF1; B = 8'hC8; #100;
A = 8'hF1; B = 8'hC9; #100;
A = 8'hF1; B = 8'hCA; #100;
A = 8'hF1; B = 8'hCB; #100;
A = 8'hF1; B = 8'hCC; #100;
A = 8'hF1; B = 8'hCD; #100;
A = 8'hF1; B = 8'hCE; #100;
A = 8'hF1; B = 8'hCF; #100;
A = 8'hF1; B = 8'hD0; #100;
A = 8'hF1; B = 8'hD1; #100;
A = 8'hF1; B = 8'hD2; #100;
A = 8'hF1; B = 8'hD3; #100;
A = 8'hF1; B = 8'hD4; #100;
A = 8'hF1; B = 8'hD5; #100;
A = 8'hF1; B = 8'hD6; #100;
A = 8'hF1; B = 8'hD7; #100;
A = 8'hF1; B = 8'hD8; #100;
A = 8'hF1; B = 8'hD9; #100;
A = 8'hF1; B = 8'hDA; #100;
A = 8'hF1; B = 8'hDB; #100;
A = 8'hF1; B = 8'hDC; #100;
A = 8'hF1; B = 8'hDD; #100;
A = 8'hF1; B = 8'hDE; #100;
A = 8'hF1; B = 8'hDF; #100;
A = 8'hF1; B = 8'hE0; #100;
A = 8'hF1; B = 8'hE1; #100;
A = 8'hF1; B = 8'hE2; #100;
A = 8'hF1; B = 8'hE3; #100;
A = 8'hF1; B = 8'hE4; #100;
A = 8'hF1; B = 8'hE5; #100;
A = 8'hF1; B = 8'hE6; #100;
A = 8'hF1; B = 8'hE7; #100;
A = 8'hF1; B = 8'hE8; #100;
A = 8'hF1; B = 8'hE9; #100;
A = 8'hF1; B = 8'hEA; #100;
A = 8'hF1; B = 8'hEB; #100;
A = 8'hF1; B = 8'hEC; #100;
A = 8'hF1; B = 8'hED; #100;
A = 8'hF1; B = 8'hEE; #100;
A = 8'hF1; B = 8'hEF; #100;
A = 8'hF1; B = 8'hF0; #100;
A = 8'hF1; B = 8'hF1; #100;
A = 8'hF1; B = 8'hF2; #100;
A = 8'hF1; B = 8'hF3; #100;
A = 8'hF1; B = 8'hF4; #100;
A = 8'hF1; B = 8'hF5; #100;
A = 8'hF1; B = 8'hF6; #100;
A = 8'hF1; B = 8'hF7; #100;
A = 8'hF1; B = 8'hF8; #100;
A = 8'hF1; B = 8'hF9; #100;
A = 8'hF1; B = 8'hFA; #100;
A = 8'hF1; B = 8'hFB; #100;
A = 8'hF1; B = 8'hFC; #100;
A = 8'hF1; B = 8'hFD; #100;
A = 8'hF1; B = 8'hFE; #100;
A = 8'hF1; B = 8'hFF; #100;
A = 8'hF2; B = 8'h0; #100;
A = 8'hF2; B = 8'h1; #100;
A = 8'hF2; B = 8'h2; #100;
A = 8'hF2; B = 8'h3; #100;
A = 8'hF2; B = 8'h4; #100;
A = 8'hF2; B = 8'h5; #100;
A = 8'hF2; B = 8'h6; #100;
A = 8'hF2; B = 8'h7; #100;
A = 8'hF2; B = 8'h8; #100;
A = 8'hF2; B = 8'h9; #100;
A = 8'hF2; B = 8'hA; #100;
A = 8'hF2; B = 8'hB; #100;
A = 8'hF2; B = 8'hC; #100;
A = 8'hF2; B = 8'hD; #100;
A = 8'hF2; B = 8'hE; #100;
A = 8'hF2; B = 8'hF; #100;
A = 8'hF2; B = 8'h10; #100;
A = 8'hF2; B = 8'h11; #100;
A = 8'hF2; B = 8'h12; #100;
A = 8'hF2; B = 8'h13; #100;
A = 8'hF2; B = 8'h14; #100;
A = 8'hF2; B = 8'h15; #100;
A = 8'hF2; B = 8'h16; #100;
A = 8'hF2; B = 8'h17; #100;
A = 8'hF2; B = 8'h18; #100;
A = 8'hF2; B = 8'h19; #100;
A = 8'hF2; B = 8'h1A; #100;
A = 8'hF2; B = 8'h1B; #100;
A = 8'hF2; B = 8'h1C; #100;
A = 8'hF2; B = 8'h1D; #100;
A = 8'hF2; B = 8'h1E; #100;
A = 8'hF2; B = 8'h1F; #100;
A = 8'hF2; B = 8'h20; #100;
A = 8'hF2; B = 8'h21; #100;
A = 8'hF2; B = 8'h22; #100;
A = 8'hF2; B = 8'h23; #100;
A = 8'hF2; B = 8'h24; #100;
A = 8'hF2; B = 8'h25; #100;
A = 8'hF2; B = 8'h26; #100;
A = 8'hF2; B = 8'h27; #100;
A = 8'hF2; B = 8'h28; #100;
A = 8'hF2; B = 8'h29; #100;
A = 8'hF2; B = 8'h2A; #100;
A = 8'hF2; B = 8'h2B; #100;
A = 8'hF2; B = 8'h2C; #100;
A = 8'hF2; B = 8'h2D; #100;
A = 8'hF2; B = 8'h2E; #100;
A = 8'hF2; B = 8'h2F; #100;
A = 8'hF2; B = 8'h30; #100;
A = 8'hF2; B = 8'h31; #100;
A = 8'hF2; B = 8'h32; #100;
A = 8'hF2; B = 8'h33; #100;
A = 8'hF2; B = 8'h34; #100;
A = 8'hF2; B = 8'h35; #100;
A = 8'hF2; B = 8'h36; #100;
A = 8'hF2; B = 8'h37; #100;
A = 8'hF2; B = 8'h38; #100;
A = 8'hF2; B = 8'h39; #100;
A = 8'hF2; B = 8'h3A; #100;
A = 8'hF2; B = 8'h3B; #100;
A = 8'hF2; B = 8'h3C; #100;
A = 8'hF2; B = 8'h3D; #100;
A = 8'hF2; B = 8'h3E; #100;
A = 8'hF2; B = 8'h3F; #100;
A = 8'hF2; B = 8'h40; #100;
A = 8'hF2; B = 8'h41; #100;
A = 8'hF2; B = 8'h42; #100;
A = 8'hF2; B = 8'h43; #100;
A = 8'hF2; B = 8'h44; #100;
A = 8'hF2; B = 8'h45; #100;
A = 8'hF2; B = 8'h46; #100;
A = 8'hF2; B = 8'h47; #100;
A = 8'hF2; B = 8'h48; #100;
A = 8'hF2; B = 8'h49; #100;
A = 8'hF2; B = 8'h4A; #100;
A = 8'hF2; B = 8'h4B; #100;
A = 8'hF2; B = 8'h4C; #100;
A = 8'hF2; B = 8'h4D; #100;
A = 8'hF2; B = 8'h4E; #100;
A = 8'hF2; B = 8'h4F; #100;
A = 8'hF2; B = 8'h50; #100;
A = 8'hF2; B = 8'h51; #100;
A = 8'hF2; B = 8'h52; #100;
A = 8'hF2; B = 8'h53; #100;
A = 8'hF2; B = 8'h54; #100;
A = 8'hF2; B = 8'h55; #100;
A = 8'hF2; B = 8'h56; #100;
A = 8'hF2; B = 8'h57; #100;
A = 8'hF2; B = 8'h58; #100;
A = 8'hF2; B = 8'h59; #100;
A = 8'hF2; B = 8'h5A; #100;
A = 8'hF2; B = 8'h5B; #100;
A = 8'hF2; B = 8'h5C; #100;
A = 8'hF2; B = 8'h5D; #100;
A = 8'hF2; B = 8'h5E; #100;
A = 8'hF2; B = 8'h5F; #100;
A = 8'hF2; B = 8'h60; #100;
A = 8'hF2; B = 8'h61; #100;
A = 8'hF2; B = 8'h62; #100;
A = 8'hF2; B = 8'h63; #100;
A = 8'hF2; B = 8'h64; #100;
A = 8'hF2; B = 8'h65; #100;
A = 8'hF2; B = 8'h66; #100;
A = 8'hF2; B = 8'h67; #100;
A = 8'hF2; B = 8'h68; #100;
A = 8'hF2; B = 8'h69; #100;
A = 8'hF2; B = 8'h6A; #100;
A = 8'hF2; B = 8'h6B; #100;
A = 8'hF2; B = 8'h6C; #100;
A = 8'hF2; B = 8'h6D; #100;
A = 8'hF2; B = 8'h6E; #100;
A = 8'hF2; B = 8'h6F; #100;
A = 8'hF2; B = 8'h70; #100;
A = 8'hF2; B = 8'h71; #100;
A = 8'hF2; B = 8'h72; #100;
A = 8'hF2; B = 8'h73; #100;
A = 8'hF2; B = 8'h74; #100;
A = 8'hF2; B = 8'h75; #100;
A = 8'hF2; B = 8'h76; #100;
A = 8'hF2; B = 8'h77; #100;
A = 8'hF2; B = 8'h78; #100;
A = 8'hF2; B = 8'h79; #100;
A = 8'hF2; B = 8'h7A; #100;
A = 8'hF2; B = 8'h7B; #100;
A = 8'hF2; B = 8'h7C; #100;
A = 8'hF2; B = 8'h7D; #100;
A = 8'hF2; B = 8'h7E; #100;
A = 8'hF2; B = 8'h7F; #100;
A = 8'hF2; B = 8'h80; #100;
A = 8'hF2; B = 8'h81; #100;
A = 8'hF2; B = 8'h82; #100;
A = 8'hF2; B = 8'h83; #100;
A = 8'hF2; B = 8'h84; #100;
A = 8'hF2; B = 8'h85; #100;
A = 8'hF2; B = 8'h86; #100;
A = 8'hF2; B = 8'h87; #100;
A = 8'hF2; B = 8'h88; #100;
A = 8'hF2; B = 8'h89; #100;
A = 8'hF2; B = 8'h8A; #100;
A = 8'hF2; B = 8'h8B; #100;
A = 8'hF2; B = 8'h8C; #100;
A = 8'hF2; B = 8'h8D; #100;
A = 8'hF2; B = 8'h8E; #100;
A = 8'hF2; B = 8'h8F; #100;
A = 8'hF2; B = 8'h90; #100;
A = 8'hF2; B = 8'h91; #100;
A = 8'hF2; B = 8'h92; #100;
A = 8'hF2; B = 8'h93; #100;
A = 8'hF2; B = 8'h94; #100;
A = 8'hF2; B = 8'h95; #100;
A = 8'hF2; B = 8'h96; #100;
A = 8'hF2; B = 8'h97; #100;
A = 8'hF2; B = 8'h98; #100;
A = 8'hF2; B = 8'h99; #100;
A = 8'hF2; B = 8'h9A; #100;
A = 8'hF2; B = 8'h9B; #100;
A = 8'hF2; B = 8'h9C; #100;
A = 8'hF2; B = 8'h9D; #100;
A = 8'hF2; B = 8'h9E; #100;
A = 8'hF2; B = 8'h9F; #100;
A = 8'hF2; B = 8'hA0; #100;
A = 8'hF2; B = 8'hA1; #100;
A = 8'hF2; B = 8'hA2; #100;
A = 8'hF2; B = 8'hA3; #100;
A = 8'hF2; B = 8'hA4; #100;
A = 8'hF2; B = 8'hA5; #100;
A = 8'hF2; B = 8'hA6; #100;
A = 8'hF2; B = 8'hA7; #100;
A = 8'hF2; B = 8'hA8; #100;
A = 8'hF2; B = 8'hA9; #100;
A = 8'hF2; B = 8'hAA; #100;
A = 8'hF2; B = 8'hAB; #100;
A = 8'hF2; B = 8'hAC; #100;
A = 8'hF2; B = 8'hAD; #100;
A = 8'hF2; B = 8'hAE; #100;
A = 8'hF2; B = 8'hAF; #100;
A = 8'hF2; B = 8'hB0; #100;
A = 8'hF2; B = 8'hB1; #100;
A = 8'hF2; B = 8'hB2; #100;
A = 8'hF2; B = 8'hB3; #100;
A = 8'hF2; B = 8'hB4; #100;
A = 8'hF2; B = 8'hB5; #100;
A = 8'hF2; B = 8'hB6; #100;
A = 8'hF2; B = 8'hB7; #100;
A = 8'hF2; B = 8'hB8; #100;
A = 8'hF2; B = 8'hB9; #100;
A = 8'hF2; B = 8'hBA; #100;
A = 8'hF2; B = 8'hBB; #100;
A = 8'hF2; B = 8'hBC; #100;
A = 8'hF2; B = 8'hBD; #100;
A = 8'hF2; B = 8'hBE; #100;
A = 8'hF2; B = 8'hBF; #100;
A = 8'hF2; B = 8'hC0; #100;
A = 8'hF2; B = 8'hC1; #100;
A = 8'hF2; B = 8'hC2; #100;
A = 8'hF2; B = 8'hC3; #100;
A = 8'hF2; B = 8'hC4; #100;
A = 8'hF2; B = 8'hC5; #100;
A = 8'hF2; B = 8'hC6; #100;
A = 8'hF2; B = 8'hC7; #100;
A = 8'hF2; B = 8'hC8; #100;
A = 8'hF2; B = 8'hC9; #100;
A = 8'hF2; B = 8'hCA; #100;
A = 8'hF2; B = 8'hCB; #100;
A = 8'hF2; B = 8'hCC; #100;
A = 8'hF2; B = 8'hCD; #100;
A = 8'hF2; B = 8'hCE; #100;
A = 8'hF2; B = 8'hCF; #100;
A = 8'hF2; B = 8'hD0; #100;
A = 8'hF2; B = 8'hD1; #100;
A = 8'hF2; B = 8'hD2; #100;
A = 8'hF2; B = 8'hD3; #100;
A = 8'hF2; B = 8'hD4; #100;
A = 8'hF2; B = 8'hD5; #100;
A = 8'hF2; B = 8'hD6; #100;
A = 8'hF2; B = 8'hD7; #100;
A = 8'hF2; B = 8'hD8; #100;
A = 8'hF2; B = 8'hD9; #100;
A = 8'hF2; B = 8'hDA; #100;
A = 8'hF2; B = 8'hDB; #100;
A = 8'hF2; B = 8'hDC; #100;
A = 8'hF2; B = 8'hDD; #100;
A = 8'hF2; B = 8'hDE; #100;
A = 8'hF2; B = 8'hDF; #100;
A = 8'hF2; B = 8'hE0; #100;
A = 8'hF2; B = 8'hE1; #100;
A = 8'hF2; B = 8'hE2; #100;
A = 8'hF2; B = 8'hE3; #100;
A = 8'hF2; B = 8'hE4; #100;
A = 8'hF2; B = 8'hE5; #100;
A = 8'hF2; B = 8'hE6; #100;
A = 8'hF2; B = 8'hE7; #100;
A = 8'hF2; B = 8'hE8; #100;
A = 8'hF2; B = 8'hE9; #100;
A = 8'hF2; B = 8'hEA; #100;
A = 8'hF2; B = 8'hEB; #100;
A = 8'hF2; B = 8'hEC; #100;
A = 8'hF2; B = 8'hED; #100;
A = 8'hF2; B = 8'hEE; #100;
A = 8'hF2; B = 8'hEF; #100;
A = 8'hF2; B = 8'hF0; #100;
A = 8'hF2; B = 8'hF1; #100;
A = 8'hF2; B = 8'hF2; #100;
A = 8'hF2; B = 8'hF3; #100;
A = 8'hF2; B = 8'hF4; #100;
A = 8'hF2; B = 8'hF5; #100;
A = 8'hF2; B = 8'hF6; #100;
A = 8'hF2; B = 8'hF7; #100;
A = 8'hF2; B = 8'hF8; #100;
A = 8'hF2; B = 8'hF9; #100;
A = 8'hF2; B = 8'hFA; #100;
A = 8'hF2; B = 8'hFB; #100;
A = 8'hF2; B = 8'hFC; #100;
A = 8'hF2; B = 8'hFD; #100;
A = 8'hF2; B = 8'hFE; #100;
A = 8'hF2; B = 8'hFF; #100;
A = 8'hF3; B = 8'h0; #100;
A = 8'hF3; B = 8'h1; #100;
A = 8'hF3; B = 8'h2; #100;
A = 8'hF3; B = 8'h3; #100;
A = 8'hF3; B = 8'h4; #100;
A = 8'hF3; B = 8'h5; #100;
A = 8'hF3; B = 8'h6; #100;
A = 8'hF3; B = 8'h7; #100;
A = 8'hF3; B = 8'h8; #100;
A = 8'hF3; B = 8'h9; #100;
A = 8'hF3; B = 8'hA; #100;
A = 8'hF3; B = 8'hB; #100;
A = 8'hF3; B = 8'hC; #100;
A = 8'hF3; B = 8'hD; #100;
A = 8'hF3; B = 8'hE; #100;
A = 8'hF3; B = 8'hF; #100;
A = 8'hF3; B = 8'h10; #100;
A = 8'hF3; B = 8'h11; #100;
A = 8'hF3; B = 8'h12; #100;
A = 8'hF3; B = 8'h13; #100;
A = 8'hF3; B = 8'h14; #100;
A = 8'hF3; B = 8'h15; #100;
A = 8'hF3; B = 8'h16; #100;
A = 8'hF3; B = 8'h17; #100;
A = 8'hF3; B = 8'h18; #100;
A = 8'hF3; B = 8'h19; #100;
A = 8'hF3; B = 8'h1A; #100;
A = 8'hF3; B = 8'h1B; #100;
A = 8'hF3; B = 8'h1C; #100;
A = 8'hF3; B = 8'h1D; #100;
A = 8'hF3; B = 8'h1E; #100;
A = 8'hF3; B = 8'h1F; #100;
A = 8'hF3; B = 8'h20; #100;
A = 8'hF3; B = 8'h21; #100;
A = 8'hF3; B = 8'h22; #100;
A = 8'hF3; B = 8'h23; #100;
A = 8'hF3; B = 8'h24; #100;
A = 8'hF3; B = 8'h25; #100;
A = 8'hF3; B = 8'h26; #100;
A = 8'hF3; B = 8'h27; #100;
A = 8'hF3; B = 8'h28; #100;
A = 8'hF3; B = 8'h29; #100;
A = 8'hF3; B = 8'h2A; #100;
A = 8'hF3; B = 8'h2B; #100;
A = 8'hF3; B = 8'h2C; #100;
A = 8'hF3; B = 8'h2D; #100;
A = 8'hF3; B = 8'h2E; #100;
A = 8'hF3; B = 8'h2F; #100;
A = 8'hF3; B = 8'h30; #100;
A = 8'hF3; B = 8'h31; #100;
A = 8'hF3; B = 8'h32; #100;
A = 8'hF3; B = 8'h33; #100;
A = 8'hF3; B = 8'h34; #100;
A = 8'hF3; B = 8'h35; #100;
A = 8'hF3; B = 8'h36; #100;
A = 8'hF3; B = 8'h37; #100;
A = 8'hF3; B = 8'h38; #100;
A = 8'hF3; B = 8'h39; #100;
A = 8'hF3; B = 8'h3A; #100;
A = 8'hF3; B = 8'h3B; #100;
A = 8'hF3; B = 8'h3C; #100;
A = 8'hF3; B = 8'h3D; #100;
A = 8'hF3; B = 8'h3E; #100;
A = 8'hF3; B = 8'h3F; #100;
A = 8'hF3; B = 8'h40; #100;
A = 8'hF3; B = 8'h41; #100;
A = 8'hF3; B = 8'h42; #100;
A = 8'hF3; B = 8'h43; #100;
A = 8'hF3; B = 8'h44; #100;
A = 8'hF3; B = 8'h45; #100;
A = 8'hF3; B = 8'h46; #100;
A = 8'hF3; B = 8'h47; #100;
A = 8'hF3; B = 8'h48; #100;
A = 8'hF3; B = 8'h49; #100;
A = 8'hF3; B = 8'h4A; #100;
A = 8'hF3; B = 8'h4B; #100;
A = 8'hF3; B = 8'h4C; #100;
A = 8'hF3; B = 8'h4D; #100;
A = 8'hF3; B = 8'h4E; #100;
A = 8'hF3; B = 8'h4F; #100;
A = 8'hF3; B = 8'h50; #100;
A = 8'hF3; B = 8'h51; #100;
A = 8'hF3; B = 8'h52; #100;
A = 8'hF3; B = 8'h53; #100;
A = 8'hF3; B = 8'h54; #100;
A = 8'hF3; B = 8'h55; #100;
A = 8'hF3; B = 8'h56; #100;
A = 8'hF3; B = 8'h57; #100;
A = 8'hF3; B = 8'h58; #100;
A = 8'hF3; B = 8'h59; #100;
A = 8'hF3; B = 8'h5A; #100;
A = 8'hF3; B = 8'h5B; #100;
A = 8'hF3; B = 8'h5C; #100;
A = 8'hF3; B = 8'h5D; #100;
A = 8'hF3; B = 8'h5E; #100;
A = 8'hF3; B = 8'h5F; #100;
A = 8'hF3; B = 8'h60; #100;
A = 8'hF3; B = 8'h61; #100;
A = 8'hF3; B = 8'h62; #100;
A = 8'hF3; B = 8'h63; #100;
A = 8'hF3; B = 8'h64; #100;
A = 8'hF3; B = 8'h65; #100;
A = 8'hF3; B = 8'h66; #100;
A = 8'hF3; B = 8'h67; #100;
A = 8'hF3; B = 8'h68; #100;
A = 8'hF3; B = 8'h69; #100;
A = 8'hF3; B = 8'h6A; #100;
A = 8'hF3; B = 8'h6B; #100;
A = 8'hF3; B = 8'h6C; #100;
A = 8'hF3; B = 8'h6D; #100;
A = 8'hF3; B = 8'h6E; #100;
A = 8'hF3; B = 8'h6F; #100;
A = 8'hF3; B = 8'h70; #100;
A = 8'hF3; B = 8'h71; #100;
A = 8'hF3; B = 8'h72; #100;
A = 8'hF3; B = 8'h73; #100;
A = 8'hF3; B = 8'h74; #100;
A = 8'hF3; B = 8'h75; #100;
A = 8'hF3; B = 8'h76; #100;
A = 8'hF3; B = 8'h77; #100;
A = 8'hF3; B = 8'h78; #100;
A = 8'hF3; B = 8'h79; #100;
A = 8'hF3; B = 8'h7A; #100;
A = 8'hF3; B = 8'h7B; #100;
A = 8'hF3; B = 8'h7C; #100;
A = 8'hF3; B = 8'h7D; #100;
A = 8'hF3; B = 8'h7E; #100;
A = 8'hF3; B = 8'h7F; #100;
A = 8'hF3; B = 8'h80; #100;
A = 8'hF3; B = 8'h81; #100;
A = 8'hF3; B = 8'h82; #100;
A = 8'hF3; B = 8'h83; #100;
A = 8'hF3; B = 8'h84; #100;
A = 8'hF3; B = 8'h85; #100;
A = 8'hF3; B = 8'h86; #100;
A = 8'hF3; B = 8'h87; #100;
A = 8'hF3; B = 8'h88; #100;
A = 8'hF3; B = 8'h89; #100;
A = 8'hF3; B = 8'h8A; #100;
A = 8'hF3; B = 8'h8B; #100;
A = 8'hF3; B = 8'h8C; #100;
A = 8'hF3; B = 8'h8D; #100;
A = 8'hF3; B = 8'h8E; #100;
A = 8'hF3; B = 8'h8F; #100;
A = 8'hF3; B = 8'h90; #100;
A = 8'hF3; B = 8'h91; #100;
A = 8'hF3; B = 8'h92; #100;
A = 8'hF3; B = 8'h93; #100;
A = 8'hF3; B = 8'h94; #100;
A = 8'hF3; B = 8'h95; #100;
A = 8'hF3; B = 8'h96; #100;
A = 8'hF3; B = 8'h97; #100;
A = 8'hF3; B = 8'h98; #100;
A = 8'hF3; B = 8'h99; #100;
A = 8'hF3; B = 8'h9A; #100;
A = 8'hF3; B = 8'h9B; #100;
A = 8'hF3; B = 8'h9C; #100;
A = 8'hF3; B = 8'h9D; #100;
A = 8'hF3; B = 8'h9E; #100;
A = 8'hF3; B = 8'h9F; #100;
A = 8'hF3; B = 8'hA0; #100;
A = 8'hF3; B = 8'hA1; #100;
A = 8'hF3; B = 8'hA2; #100;
A = 8'hF3; B = 8'hA3; #100;
A = 8'hF3; B = 8'hA4; #100;
A = 8'hF3; B = 8'hA5; #100;
A = 8'hF3; B = 8'hA6; #100;
A = 8'hF3; B = 8'hA7; #100;
A = 8'hF3; B = 8'hA8; #100;
A = 8'hF3; B = 8'hA9; #100;
A = 8'hF3; B = 8'hAA; #100;
A = 8'hF3; B = 8'hAB; #100;
A = 8'hF3; B = 8'hAC; #100;
A = 8'hF3; B = 8'hAD; #100;
A = 8'hF3; B = 8'hAE; #100;
A = 8'hF3; B = 8'hAF; #100;
A = 8'hF3; B = 8'hB0; #100;
A = 8'hF3; B = 8'hB1; #100;
A = 8'hF3; B = 8'hB2; #100;
A = 8'hF3; B = 8'hB3; #100;
A = 8'hF3; B = 8'hB4; #100;
A = 8'hF3; B = 8'hB5; #100;
A = 8'hF3; B = 8'hB6; #100;
A = 8'hF3; B = 8'hB7; #100;
A = 8'hF3; B = 8'hB8; #100;
A = 8'hF3; B = 8'hB9; #100;
A = 8'hF3; B = 8'hBA; #100;
A = 8'hF3; B = 8'hBB; #100;
A = 8'hF3; B = 8'hBC; #100;
A = 8'hF3; B = 8'hBD; #100;
A = 8'hF3; B = 8'hBE; #100;
A = 8'hF3; B = 8'hBF; #100;
A = 8'hF3; B = 8'hC0; #100;
A = 8'hF3; B = 8'hC1; #100;
A = 8'hF3; B = 8'hC2; #100;
A = 8'hF3; B = 8'hC3; #100;
A = 8'hF3; B = 8'hC4; #100;
A = 8'hF3; B = 8'hC5; #100;
A = 8'hF3; B = 8'hC6; #100;
A = 8'hF3; B = 8'hC7; #100;
A = 8'hF3; B = 8'hC8; #100;
A = 8'hF3; B = 8'hC9; #100;
A = 8'hF3; B = 8'hCA; #100;
A = 8'hF3; B = 8'hCB; #100;
A = 8'hF3; B = 8'hCC; #100;
A = 8'hF3; B = 8'hCD; #100;
A = 8'hF3; B = 8'hCE; #100;
A = 8'hF3; B = 8'hCF; #100;
A = 8'hF3; B = 8'hD0; #100;
A = 8'hF3; B = 8'hD1; #100;
A = 8'hF3; B = 8'hD2; #100;
A = 8'hF3; B = 8'hD3; #100;
A = 8'hF3; B = 8'hD4; #100;
A = 8'hF3; B = 8'hD5; #100;
A = 8'hF3; B = 8'hD6; #100;
A = 8'hF3; B = 8'hD7; #100;
A = 8'hF3; B = 8'hD8; #100;
A = 8'hF3; B = 8'hD9; #100;
A = 8'hF3; B = 8'hDA; #100;
A = 8'hF3; B = 8'hDB; #100;
A = 8'hF3; B = 8'hDC; #100;
A = 8'hF3; B = 8'hDD; #100;
A = 8'hF3; B = 8'hDE; #100;
A = 8'hF3; B = 8'hDF; #100;
A = 8'hF3; B = 8'hE0; #100;
A = 8'hF3; B = 8'hE1; #100;
A = 8'hF3; B = 8'hE2; #100;
A = 8'hF3; B = 8'hE3; #100;
A = 8'hF3; B = 8'hE4; #100;
A = 8'hF3; B = 8'hE5; #100;
A = 8'hF3; B = 8'hE6; #100;
A = 8'hF3; B = 8'hE7; #100;
A = 8'hF3; B = 8'hE8; #100;
A = 8'hF3; B = 8'hE9; #100;
A = 8'hF3; B = 8'hEA; #100;
A = 8'hF3; B = 8'hEB; #100;
A = 8'hF3; B = 8'hEC; #100;
A = 8'hF3; B = 8'hED; #100;
A = 8'hF3; B = 8'hEE; #100;
A = 8'hF3; B = 8'hEF; #100;
A = 8'hF3; B = 8'hF0; #100;
A = 8'hF3; B = 8'hF1; #100;
A = 8'hF3; B = 8'hF2; #100;
A = 8'hF3; B = 8'hF3; #100;
A = 8'hF3; B = 8'hF4; #100;
A = 8'hF3; B = 8'hF5; #100;
A = 8'hF3; B = 8'hF6; #100;
A = 8'hF3; B = 8'hF7; #100;
A = 8'hF3; B = 8'hF8; #100;
A = 8'hF3; B = 8'hF9; #100;
A = 8'hF3; B = 8'hFA; #100;
A = 8'hF3; B = 8'hFB; #100;
A = 8'hF3; B = 8'hFC; #100;
A = 8'hF3; B = 8'hFD; #100;
A = 8'hF3; B = 8'hFE; #100;
A = 8'hF3; B = 8'hFF; #100;
A = 8'hF4; B = 8'h0; #100;
A = 8'hF4; B = 8'h1; #100;
A = 8'hF4; B = 8'h2; #100;
A = 8'hF4; B = 8'h3; #100;
A = 8'hF4; B = 8'h4; #100;
A = 8'hF4; B = 8'h5; #100;
A = 8'hF4; B = 8'h6; #100;
A = 8'hF4; B = 8'h7; #100;
A = 8'hF4; B = 8'h8; #100;
A = 8'hF4; B = 8'h9; #100;
A = 8'hF4; B = 8'hA; #100;
A = 8'hF4; B = 8'hB; #100;
A = 8'hF4; B = 8'hC; #100;
A = 8'hF4; B = 8'hD; #100;
A = 8'hF4; B = 8'hE; #100;
A = 8'hF4; B = 8'hF; #100;
A = 8'hF4; B = 8'h10; #100;
A = 8'hF4; B = 8'h11; #100;
A = 8'hF4; B = 8'h12; #100;
A = 8'hF4; B = 8'h13; #100;
A = 8'hF4; B = 8'h14; #100;
A = 8'hF4; B = 8'h15; #100;
A = 8'hF4; B = 8'h16; #100;
A = 8'hF4; B = 8'h17; #100;
A = 8'hF4; B = 8'h18; #100;
A = 8'hF4; B = 8'h19; #100;
A = 8'hF4; B = 8'h1A; #100;
A = 8'hF4; B = 8'h1B; #100;
A = 8'hF4; B = 8'h1C; #100;
A = 8'hF4; B = 8'h1D; #100;
A = 8'hF4; B = 8'h1E; #100;
A = 8'hF4; B = 8'h1F; #100;
A = 8'hF4; B = 8'h20; #100;
A = 8'hF4; B = 8'h21; #100;
A = 8'hF4; B = 8'h22; #100;
A = 8'hF4; B = 8'h23; #100;
A = 8'hF4; B = 8'h24; #100;
A = 8'hF4; B = 8'h25; #100;
A = 8'hF4; B = 8'h26; #100;
A = 8'hF4; B = 8'h27; #100;
A = 8'hF4; B = 8'h28; #100;
A = 8'hF4; B = 8'h29; #100;
A = 8'hF4; B = 8'h2A; #100;
A = 8'hF4; B = 8'h2B; #100;
A = 8'hF4; B = 8'h2C; #100;
A = 8'hF4; B = 8'h2D; #100;
A = 8'hF4; B = 8'h2E; #100;
A = 8'hF4; B = 8'h2F; #100;
A = 8'hF4; B = 8'h30; #100;
A = 8'hF4; B = 8'h31; #100;
A = 8'hF4; B = 8'h32; #100;
A = 8'hF4; B = 8'h33; #100;
A = 8'hF4; B = 8'h34; #100;
A = 8'hF4; B = 8'h35; #100;
A = 8'hF4; B = 8'h36; #100;
A = 8'hF4; B = 8'h37; #100;
A = 8'hF4; B = 8'h38; #100;
A = 8'hF4; B = 8'h39; #100;
A = 8'hF4; B = 8'h3A; #100;
A = 8'hF4; B = 8'h3B; #100;
A = 8'hF4; B = 8'h3C; #100;
A = 8'hF4; B = 8'h3D; #100;
A = 8'hF4; B = 8'h3E; #100;
A = 8'hF4; B = 8'h3F; #100;
A = 8'hF4; B = 8'h40; #100;
A = 8'hF4; B = 8'h41; #100;
A = 8'hF4; B = 8'h42; #100;
A = 8'hF4; B = 8'h43; #100;
A = 8'hF4; B = 8'h44; #100;
A = 8'hF4; B = 8'h45; #100;
A = 8'hF4; B = 8'h46; #100;
A = 8'hF4; B = 8'h47; #100;
A = 8'hF4; B = 8'h48; #100;
A = 8'hF4; B = 8'h49; #100;
A = 8'hF4; B = 8'h4A; #100;
A = 8'hF4; B = 8'h4B; #100;
A = 8'hF4; B = 8'h4C; #100;
A = 8'hF4; B = 8'h4D; #100;
A = 8'hF4; B = 8'h4E; #100;
A = 8'hF4; B = 8'h4F; #100;
A = 8'hF4; B = 8'h50; #100;
A = 8'hF4; B = 8'h51; #100;
A = 8'hF4; B = 8'h52; #100;
A = 8'hF4; B = 8'h53; #100;
A = 8'hF4; B = 8'h54; #100;
A = 8'hF4; B = 8'h55; #100;
A = 8'hF4; B = 8'h56; #100;
A = 8'hF4; B = 8'h57; #100;
A = 8'hF4; B = 8'h58; #100;
A = 8'hF4; B = 8'h59; #100;
A = 8'hF4; B = 8'h5A; #100;
A = 8'hF4; B = 8'h5B; #100;
A = 8'hF4; B = 8'h5C; #100;
A = 8'hF4; B = 8'h5D; #100;
A = 8'hF4; B = 8'h5E; #100;
A = 8'hF4; B = 8'h5F; #100;
A = 8'hF4; B = 8'h60; #100;
A = 8'hF4; B = 8'h61; #100;
A = 8'hF4; B = 8'h62; #100;
A = 8'hF4; B = 8'h63; #100;
A = 8'hF4; B = 8'h64; #100;
A = 8'hF4; B = 8'h65; #100;
A = 8'hF4; B = 8'h66; #100;
A = 8'hF4; B = 8'h67; #100;
A = 8'hF4; B = 8'h68; #100;
A = 8'hF4; B = 8'h69; #100;
A = 8'hF4; B = 8'h6A; #100;
A = 8'hF4; B = 8'h6B; #100;
A = 8'hF4; B = 8'h6C; #100;
A = 8'hF4; B = 8'h6D; #100;
A = 8'hF4; B = 8'h6E; #100;
A = 8'hF4; B = 8'h6F; #100;
A = 8'hF4; B = 8'h70; #100;
A = 8'hF4; B = 8'h71; #100;
A = 8'hF4; B = 8'h72; #100;
A = 8'hF4; B = 8'h73; #100;
A = 8'hF4; B = 8'h74; #100;
A = 8'hF4; B = 8'h75; #100;
A = 8'hF4; B = 8'h76; #100;
A = 8'hF4; B = 8'h77; #100;
A = 8'hF4; B = 8'h78; #100;
A = 8'hF4; B = 8'h79; #100;
A = 8'hF4; B = 8'h7A; #100;
A = 8'hF4; B = 8'h7B; #100;
A = 8'hF4; B = 8'h7C; #100;
A = 8'hF4; B = 8'h7D; #100;
A = 8'hF4; B = 8'h7E; #100;
A = 8'hF4; B = 8'h7F; #100;
A = 8'hF4; B = 8'h80; #100;
A = 8'hF4; B = 8'h81; #100;
A = 8'hF4; B = 8'h82; #100;
A = 8'hF4; B = 8'h83; #100;
A = 8'hF4; B = 8'h84; #100;
A = 8'hF4; B = 8'h85; #100;
A = 8'hF4; B = 8'h86; #100;
A = 8'hF4; B = 8'h87; #100;
A = 8'hF4; B = 8'h88; #100;
A = 8'hF4; B = 8'h89; #100;
A = 8'hF4; B = 8'h8A; #100;
A = 8'hF4; B = 8'h8B; #100;
A = 8'hF4; B = 8'h8C; #100;
A = 8'hF4; B = 8'h8D; #100;
A = 8'hF4; B = 8'h8E; #100;
A = 8'hF4; B = 8'h8F; #100;
A = 8'hF4; B = 8'h90; #100;
A = 8'hF4; B = 8'h91; #100;
A = 8'hF4; B = 8'h92; #100;
A = 8'hF4; B = 8'h93; #100;
A = 8'hF4; B = 8'h94; #100;
A = 8'hF4; B = 8'h95; #100;
A = 8'hF4; B = 8'h96; #100;
A = 8'hF4; B = 8'h97; #100;
A = 8'hF4; B = 8'h98; #100;
A = 8'hF4; B = 8'h99; #100;
A = 8'hF4; B = 8'h9A; #100;
A = 8'hF4; B = 8'h9B; #100;
A = 8'hF4; B = 8'h9C; #100;
A = 8'hF4; B = 8'h9D; #100;
A = 8'hF4; B = 8'h9E; #100;
A = 8'hF4; B = 8'h9F; #100;
A = 8'hF4; B = 8'hA0; #100;
A = 8'hF4; B = 8'hA1; #100;
A = 8'hF4; B = 8'hA2; #100;
A = 8'hF4; B = 8'hA3; #100;
A = 8'hF4; B = 8'hA4; #100;
A = 8'hF4; B = 8'hA5; #100;
A = 8'hF4; B = 8'hA6; #100;
A = 8'hF4; B = 8'hA7; #100;
A = 8'hF4; B = 8'hA8; #100;
A = 8'hF4; B = 8'hA9; #100;
A = 8'hF4; B = 8'hAA; #100;
A = 8'hF4; B = 8'hAB; #100;
A = 8'hF4; B = 8'hAC; #100;
A = 8'hF4; B = 8'hAD; #100;
A = 8'hF4; B = 8'hAE; #100;
A = 8'hF4; B = 8'hAF; #100;
A = 8'hF4; B = 8'hB0; #100;
A = 8'hF4; B = 8'hB1; #100;
A = 8'hF4; B = 8'hB2; #100;
A = 8'hF4; B = 8'hB3; #100;
A = 8'hF4; B = 8'hB4; #100;
A = 8'hF4; B = 8'hB5; #100;
A = 8'hF4; B = 8'hB6; #100;
A = 8'hF4; B = 8'hB7; #100;
A = 8'hF4; B = 8'hB8; #100;
A = 8'hF4; B = 8'hB9; #100;
A = 8'hF4; B = 8'hBA; #100;
A = 8'hF4; B = 8'hBB; #100;
A = 8'hF4; B = 8'hBC; #100;
A = 8'hF4; B = 8'hBD; #100;
A = 8'hF4; B = 8'hBE; #100;
A = 8'hF4; B = 8'hBF; #100;
A = 8'hF4; B = 8'hC0; #100;
A = 8'hF4; B = 8'hC1; #100;
A = 8'hF4; B = 8'hC2; #100;
A = 8'hF4; B = 8'hC3; #100;
A = 8'hF4; B = 8'hC4; #100;
A = 8'hF4; B = 8'hC5; #100;
A = 8'hF4; B = 8'hC6; #100;
A = 8'hF4; B = 8'hC7; #100;
A = 8'hF4; B = 8'hC8; #100;
A = 8'hF4; B = 8'hC9; #100;
A = 8'hF4; B = 8'hCA; #100;
A = 8'hF4; B = 8'hCB; #100;
A = 8'hF4; B = 8'hCC; #100;
A = 8'hF4; B = 8'hCD; #100;
A = 8'hF4; B = 8'hCE; #100;
A = 8'hF4; B = 8'hCF; #100;
A = 8'hF4; B = 8'hD0; #100;
A = 8'hF4; B = 8'hD1; #100;
A = 8'hF4; B = 8'hD2; #100;
A = 8'hF4; B = 8'hD3; #100;
A = 8'hF4; B = 8'hD4; #100;
A = 8'hF4; B = 8'hD5; #100;
A = 8'hF4; B = 8'hD6; #100;
A = 8'hF4; B = 8'hD7; #100;
A = 8'hF4; B = 8'hD8; #100;
A = 8'hF4; B = 8'hD9; #100;
A = 8'hF4; B = 8'hDA; #100;
A = 8'hF4; B = 8'hDB; #100;
A = 8'hF4; B = 8'hDC; #100;
A = 8'hF4; B = 8'hDD; #100;
A = 8'hF4; B = 8'hDE; #100;
A = 8'hF4; B = 8'hDF; #100;
A = 8'hF4; B = 8'hE0; #100;
A = 8'hF4; B = 8'hE1; #100;
A = 8'hF4; B = 8'hE2; #100;
A = 8'hF4; B = 8'hE3; #100;
A = 8'hF4; B = 8'hE4; #100;
A = 8'hF4; B = 8'hE5; #100;
A = 8'hF4; B = 8'hE6; #100;
A = 8'hF4; B = 8'hE7; #100;
A = 8'hF4; B = 8'hE8; #100;
A = 8'hF4; B = 8'hE9; #100;
A = 8'hF4; B = 8'hEA; #100;
A = 8'hF4; B = 8'hEB; #100;
A = 8'hF4; B = 8'hEC; #100;
A = 8'hF4; B = 8'hED; #100;
A = 8'hF4; B = 8'hEE; #100;
A = 8'hF4; B = 8'hEF; #100;
A = 8'hF4; B = 8'hF0; #100;
A = 8'hF4; B = 8'hF1; #100;
A = 8'hF4; B = 8'hF2; #100;
A = 8'hF4; B = 8'hF3; #100;
A = 8'hF4; B = 8'hF4; #100;
A = 8'hF4; B = 8'hF5; #100;
A = 8'hF4; B = 8'hF6; #100;
A = 8'hF4; B = 8'hF7; #100;
A = 8'hF4; B = 8'hF8; #100;
A = 8'hF4; B = 8'hF9; #100;
A = 8'hF4; B = 8'hFA; #100;
A = 8'hF4; B = 8'hFB; #100;
A = 8'hF4; B = 8'hFC; #100;
A = 8'hF4; B = 8'hFD; #100;
A = 8'hF4; B = 8'hFE; #100;
A = 8'hF4; B = 8'hFF; #100;
A = 8'hF5; B = 8'h0; #100;
A = 8'hF5; B = 8'h1; #100;
A = 8'hF5; B = 8'h2; #100;
A = 8'hF5; B = 8'h3; #100;
A = 8'hF5; B = 8'h4; #100;
A = 8'hF5; B = 8'h5; #100;
A = 8'hF5; B = 8'h6; #100;
A = 8'hF5; B = 8'h7; #100;
A = 8'hF5; B = 8'h8; #100;
A = 8'hF5; B = 8'h9; #100;
A = 8'hF5; B = 8'hA; #100;
A = 8'hF5; B = 8'hB; #100;
A = 8'hF5; B = 8'hC; #100;
A = 8'hF5; B = 8'hD; #100;
A = 8'hF5; B = 8'hE; #100;
A = 8'hF5; B = 8'hF; #100;
A = 8'hF5; B = 8'h10; #100;
A = 8'hF5; B = 8'h11; #100;
A = 8'hF5; B = 8'h12; #100;
A = 8'hF5; B = 8'h13; #100;
A = 8'hF5; B = 8'h14; #100;
A = 8'hF5; B = 8'h15; #100;
A = 8'hF5; B = 8'h16; #100;
A = 8'hF5; B = 8'h17; #100;
A = 8'hF5; B = 8'h18; #100;
A = 8'hF5; B = 8'h19; #100;
A = 8'hF5; B = 8'h1A; #100;
A = 8'hF5; B = 8'h1B; #100;
A = 8'hF5; B = 8'h1C; #100;
A = 8'hF5; B = 8'h1D; #100;
A = 8'hF5; B = 8'h1E; #100;
A = 8'hF5; B = 8'h1F; #100;
A = 8'hF5; B = 8'h20; #100;
A = 8'hF5; B = 8'h21; #100;
A = 8'hF5; B = 8'h22; #100;
A = 8'hF5; B = 8'h23; #100;
A = 8'hF5; B = 8'h24; #100;
A = 8'hF5; B = 8'h25; #100;
A = 8'hF5; B = 8'h26; #100;
A = 8'hF5; B = 8'h27; #100;
A = 8'hF5; B = 8'h28; #100;
A = 8'hF5; B = 8'h29; #100;
A = 8'hF5; B = 8'h2A; #100;
A = 8'hF5; B = 8'h2B; #100;
A = 8'hF5; B = 8'h2C; #100;
A = 8'hF5; B = 8'h2D; #100;
A = 8'hF5; B = 8'h2E; #100;
A = 8'hF5; B = 8'h2F; #100;
A = 8'hF5; B = 8'h30; #100;
A = 8'hF5; B = 8'h31; #100;
A = 8'hF5; B = 8'h32; #100;
A = 8'hF5; B = 8'h33; #100;
A = 8'hF5; B = 8'h34; #100;
A = 8'hF5; B = 8'h35; #100;
A = 8'hF5; B = 8'h36; #100;
A = 8'hF5; B = 8'h37; #100;
A = 8'hF5; B = 8'h38; #100;
A = 8'hF5; B = 8'h39; #100;
A = 8'hF5; B = 8'h3A; #100;
A = 8'hF5; B = 8'h3B; #100;
A = 8'hF5; B = 8'h3C; #100;
A = 8'hF5; B = 8'h3D; #100;
A = 8'hF5; B = 8'h3E; #100;
A = 8'hF5; B = 8'h3F; #100;
A = 8'hF5; B = 8'h40; #100;
A = 8'hF5; B = 8'h41; #100;
A = 8'hF5; B = 8'h42; #100;
A = 8'hF5; B = 8'h43; #100;
A = 8'hF5; B = 8'h44; #100;
A = 8'hF5; B = 8'h45; #100;
A = 8'hF5; B = 8'h46; #100;
A = 8'hF5; B = 8'h47; #100;
A = 8'hF5; B = 8'h48; #100;
A = 8'hF5; B = 8'h49; #100;
A = 8'hF5; B = 8'h4A; #100;
A = 8'hF5; B = 8'h4B; #100;
A = 8'hF5; B = 8'h4C; #100;
A = 8'hF5; B = 8'h4D; #100;
A = 8'hF5; B = 8'h4E; #100;
A = 8'hF5; B = 8'h4F; #100;
A = 8'hF5; B = 8'h50; #100;
A = 8'hF5; B = 8'h51; #100;
A = 8'hF5; B = 8'h52; #100;
A = 8'hF5; B = 8'h53; #100;
A = 8'hF5; B = 8'h54; #100;
A = 8'hF5; B = 8'h55; #100;
A = 8'hF5; B = 8'h56; #100;
A = 8'hF5; B = 8'h57; #100;
A = 8'hF5; B = 8'h58; #100;
A = 8'hF5; B = 8'h59; #100;
A = 8'hF5; B = 8'h5A; #100;
A = 8'hF5; B = 8'h5B; #100;
A = 8'hF5; B = 8'h5C; #100;
A = 8'hF5; B = 8'h5D; #100;
A = 8'hF5; B = 8'h5E; #100;
A = 8'hF5; B = 8'h5F; #100;
A = 8'hF5; B = 8'h60; #100;
A = 8'hF5; B = 8'h61; #100;
A = 8'hF5; B = 8'h62; #100;
A = 8'hF5; B = 8'h63; #100;
A = 8'hF5; B = 8'h64; #100;
A = 8'hF5; B = 8'h65; #100;
A = 8'hF5; B = 8'h66; #100;
A = 8'hF5; B = 8'h67; #100;
A = 8'hF5; B = 8'h68; #100;
A = 8'hF5; B = 8'h69; #100;
A = 8'hF5; B = 8'h6A; #100;
A = 8'hF5; B = 8'h6B; #100;
A = 8'hF5; B = 8'h6C; #100;
A = 8'hF5; B = 8'h6D; #100;
A = 8'hF5; B = 8'h6E; #100;
A = 8'hF5; B = 8'h6F; #100;
A = 8'hF5; B = 8'h70; #100;
A = 8'hF5; B = 8'h71; #100;
A = 8'hF5; B = 8'h72; #100;
A = 8'hF5; B = 8'h73; #100;
A = 8'hF5; B = 8'h74; #100;
A = 8'hF5; B = 8'h75; #100;
A = 8'hF5; B = 8'h76; #100;
A = 8'hF5; B = 8'h77; #100;
A = 8'hF5; B = 8'h78; #100;
A = 8'hF5; B = 8'h79; #100;
A = 8'hF5; B = 8'h7A; #100;
A = 8'hF5; B = 8'h7B; #100;
A = 8'hF5; B = 8'h7C; #100;
A = 8'hF5; B = 8'h7D; #100;
A = 8'hF5; B = 8'h7E; #100;
A = 8'hF5; B = 8'h7F; #100;
A = 8'hF5; B = 8'h80; #100;
A = 8'hF5; B = 8'h81; #100;
A = 8'hF5; B = 8'h82; #100;
A = 8'hF5; B = 8'h83; #100;
A = 8'hF5; B = 8'h84; #100;
A = 8'hF5; B = 8'h85; #100;
A = 8'hF5; B = 8'h86; #100;
A = 8'hF5; B = 8'h87; #100;
A = 8'hF5; B = 8'h88; #100;
A = 8'hF5; B = 8'h89; #100;
A = 8'hF5; B = 8'h8A; #100;
A = 8'hF5; B = 8'h8B; #100;
A = 8'hF5; B = 8'h8C; #100;
A = 8'hF5; B = 8'h8D; #100;
A = 8'hF5; B = 8'h8E; #100;
A = 8'hF5; B = 8'h8F; #100;
A = 8'hF5; B = 8'h90; #100;
A = 8'hF5; B = 8'h91; #100;
A = 8'hF5; B = 8'h92; #100;
A = 8'hF5; B = 8'h93; #100;
A = 8'hF5; B = 8'h94; #100;
A = 8'hF5; B = 8'h95; #100;
A = 8'hF5; B = 8'h96; #100;
A = 8'hF5; B = 8'h97; #100;
A = 8'hF5; B = 8'h98; #100;
A = 8'hF5; B = 8'h99; #100;
A = 8'hF5; B = 8'h9A; #100;
A = 8'hF5; B = 8'h9B; #100;
A = 8'hF5; B = 8'h9C; #100;
A = 8'hF5; B = 8'h9D; #100;
A = 8'hF5; B = 8'h9E; #100;
A = 8'hF5; B = 8'h9F; #100;
A = 8'hF5; B = 8'hA0; #100;
A = 8'hF5; B = 8'hA1; #100;
A = 8'hF5; B = 8'hA2; #100;
A = 8'hF5; B = 8'hA3; #100;
A = 8'hF5; B = 8'hA4; #100;
A = 8'hF5; B = 8'hA5; #100;
A = 8'hF5; B = 8'hA6; #100;
A = 8'hF5; B = 8'hA7; #100;
A = 8'hF5; B = 8'hA8; #100;
A = 8'hF5; B = 8'hA9; #100;
A = 8'hF5; B = 8'hAA; #100;
A = 8'hF5; B = 8'hAB; #100;
A = 8'hF5; B = 8'hAC; #100;
A = 8'hF5; B = 8'hAD; #100;
A = 8'hF5; B = 8'hAE; #100;
A = 8'hF5; B = 8'hAF; #100;
A = 8'hF5; B = 8'hB0; #100;
A = 8'hF5; B = 8'hB1; #100;
A = 8'hF5; B = 8'hB2; #100;
A = 8'hF5; B = 8'hB3; #100;
A = 8'hF5; B = 8'hB4; #100;
A = 8'hF5; B = 8'hB5; #100;
A = 8'hF5; B = 8'hB6; #100;
A = 8'hF5; B = 8'hB7; #100;
A = 8'hF5; B = 8'hB8; #100;
A = 8'hF5; B = 8'hB9; #100;
A = 8'hF5; B = 8'hBA; #100;
A = 8'hF5; B = 8'hBB; #100;
A = 8'hF5; B = 8'hBC; #100;
A = 8'hF5; B = 8'hBD; #100;
A = 8'hF5; B = 8'hBE; #100;
A = 8'hF5; B = 8'hBF; #100;
A = 8'hF5; B = 8'hC0; #100;
A = 8'hF5; B = 8'hC1; #100;
A = 8'hF5; B = 8'hC2; #100;
A = 8'hF5; B = 8'hC3; #100;
A = 8'hF5; B = 8'hC4; #100;
A = 8'hF5; B = 8'hC5; #100;
A = 8'hF5; B = 8'hC6; #100;
A = 8'hF5; B = 8'hC7; #100;
A = 8'hF5; B = 8'hC8; #100;
A = 8'hF5; B = 8'hC9; #100;
A = 8'hF5; B = 8'hCA; #100;
A = 8'hF5; B = 8'hCB; #100;
A = 8'hF5; B = 8'hCC; #100;
A = 8'hF5; B = 8'hCD; #100;
A = 8'hF5; B = 8'hCE; #100;
A = 8'hF5; B = 8'hCF; #100;
A = 8'hF5; B = 8'hD0; #100;
A = 8'hF5; B = 8'hD1; #100;
A = 8'hF5; B = 8'hD2; #100;
A = 8'hF5; B = 8'hD3; #100;
A = 8'hF5; B = 8'hD4; #100;
A = 8'hF5; B = 8'hD5; #100;
A = 8'hF5; B = 8'hD6; #100;
A = 8'hF5; B = 8'hD7; #100;
A = 8'hF5; B = 8'hD8; #100;
A = 8'hF5; B = 8'hD9; #100;
A = 8'hF5; B = 8'hDA; #100;
A = 8'hF5; B = 8'hDB; #100;
A = 8'hF5; B = 8'hDC; #100;
A = 8'hF5; B = 8'hDD; #100;
A = 8'hF5; B = 8'hDE; #100;
A = 8'hF5; B = 8'hDF; #100;
A = 8'hF5; B = 8'hE0; #100;
A = 8'hF5; B = 8'hE1; #100;
A = 8'hF5; B = 8'hE2; #100;
A = 8'hF5; B = 8'hE3; #100;
A = 8'hF5; B = 8'hE4; #100;
A = 8'hF5; B = 8'hE5; #100;
A = 8'hF5; B = 8'hE6; #100;
A = 8'hF5; B = 8'hE7; #100;
A = 8'hF5; B = 8'hE8; #100;
A = 8'hF5; B = 8'hE9; #100;
A = 8'hF5; B = 8'hEA; #100;
A = 8'hF5; B = 8'hEB; #100;
A = 8'hF5; B = 8'hEC; #100;
A = 8'hF5; B = 8'hED; #100;
A = 8'hF5; B = 8'hEE; #100;
A = 8'hF5; B = 8'hEF; #100;
A = 8'hF5; B = 8'hF0; #100;
A = 8'hF5; B = 8'hF1; #100;
A = 8'hF5; B = 8'hF2; #100;
A = 8'hF5; B = 8'hF3; #100;
A = 8'hF5; B = 8'hF4; #100;
A = 8'hF5; B = 8'hF5; #100;
A = 8'hF5; B = 8'hF6; #100;
A = 8'hF5; B = 8'hF7; #100;
A = 8'hF5; B = 8'hF8; #100;
A = 8'hF5; B = 8'hF9; #100;
A = 8'hF5; B = 8'hFA; #100;
A = 8'hF5; B = 8'hFB; #100;
A = 8'hF5; B = 8'hFC; #100;
A = 8'hF5; B = 8'hFD; #100;
A = 8'hF5; B = 8'hFE; #100;
A = 8'hF5; B = 8'hFF; #100;
A = 8'hF6; B = 8'h0; #100;
A = 8'hF6; B = 8'h1; #100;
A = 8'hF6; B = 8'h2; #100;
A = 8'hF6; B = 8'h3; #100;
A = 8'hF6; B = 8'h4; #100;
A = 8'hF6; B = 8'h5; #100;
A = 8'hF6; B = 8'h6; #100;
A = 8'hF6; B = 8'h7; #100;
A = 8'hF6; B = 8'h8; #100;
A = 8'hF6; B = 8'h9; #100;
A = 8'hF6; B = 8'hA; #100;
A = 8'hF6; B = 8'hB; #100;
A = 8'hF6; B = 8'hC; #100;
A = 8'hF6; B = 8'hD; #100;
A = 8'hF6; B = 8'hE; #100;
A = 8'hF6; B = 8'hF; #100;
A = 8'hF6; B = 8'h10; #100;
A = 8'hF6; B = 8'h11; #100;
A = 8'hF6; B = 8'h12; #100;
A = 8'hF6; B = 8'h13; #100;
A = 8'hF6; B = 8'h14; #100;
A = 8'hF6; B = 8'h15; #100;
A = 8'hF6; B = 8'h16; #100;
A = 8'hF6; B = 8'h17; #100;
A = 8'hF6; B = 8'h18; #100;
A = 8'hF6; B = 8'h19; #100;
A = 8'hF6; B = 8'h1A; #100;
A = 8'hF6; B = 8'h1B; #100;
A = 8'hF6; B = 8'h1C; #100;
A = 8'hF6; B = 8'h1D; #100;
A = 8'hF6; B = 8'h1E; #100;
A = 8'hF6; B = 8'h1F; #100;
A = 8'hF6; B = 8'h20; #100;
A = 8'hF6; B = 8'h21; #100;
A = 8'hF6; B = 8'h22; #100;
A = 8'hF6; B = 8'h23; #100;
A = 8'hF6; B = 8'h24; #100;
A = 8'hF6; B = 8'h25; #100;
A = 8'hF6; B = 8'h26; #100;
A = 8'hF6; B = 8'h27; #100;
A = 8'hF6; B = 8'h28; #100;
A = 8'hF6; B = 8'h29; #100;
A = 8'hF6; B = 8'h2A; #100;
A = 8'hF6; B = 8'h2B; #100;
A = 8'hF6; B = 8'h2C; #100;
A = 8'hF6; B = 8'h2D; #100;
A = 8'hF6; B = 8'h2E; #100;
A = 8'hF6; B = 8'h2F; #100;
A = 8'hF6; B = 8'h30; #100;
A = 8'hF6; B = 8'h31; #100;
A = 8'hF6; B = 8'h32; #100;
A = 8'hF6; B = 8'h33; #100;
A = 8'hF6; B = 8'h34; #100;
A = 8'hF6; B = 8'h35; #100;
A = 8'hF6; B = 8'h36; #100;
A = 8'hF6; B = 8'h37; #100;
A = 8'hF6; B = 8'h38; #100;
A = 8'hF6; B = 8'h39; #100;
A = 8'hF6; B = 8'h3A; #100;
A = 8'hF6; B = 8'h3B; #100;
A = 8'hF6; B = 8'h3C; #100;
A = 8'hF6; B = 8'h3D; #100;
A = 8'hF6; B = 8'h3E; #100;
A = 8'hF6; B = 8'h3F; #100;
A = 8'hF6; B = 8'h40; #100;
A = 8'hF6; B = 8'h41; #100;
A = 8'hF6; B = 8'h42; #100;
A = 8'hF6; B = 8'h43; #100;
A = 8'hF6; B = 8'h44; #100;
A = 8'hF6; B = 8'h45; #100;
A = 8'hF6; B = 8'h46; #100;
A = 8'hF6; B = 8'h47; #100;
A = 8'hF6; B = 8'h48; #100;
A = 8'hF6; B = 8'h49; #100;
A = 8'hF6; B = 8'h4A; #100;
A = 8'hF6; B = 8'h4B; #100;
A = 8'hF6; B = 8'h4C; #100;
A = 8'hF6; B = 8'h4D; #100;
A = 8'hF6; B = 8'h4E; #100;
A = 8'hF6; B = 8'h4F; #100;
A = 8'hF6; B = 8'h50; #100;
A = 8'hF6; B = 8'h51; #100;
A = 8'hF6; B = 8'h52; #100;
A = 8'hF6; B = 8'h53; #100;
A = 8'hF6; B = 8'h54; #100;
A = 8'hF6; B = 8'h55; #100;
A = 8'hF6; B = 8'h56; #100;
A = 8'hF6; B = 8'h57; #100;
A = 8'hF6; B = 8'h58; #100;
A = 8'hF6; B = 8'h59; #100;
A = 8'hF6; B = 8'h5A; #100;
A = 8'hF6; B = 8'h5B; #100;
A = 8'hF6; B = 8'h5C; #100;
A = 8'hF6; B = 8'h5D; #100;
A = 8'hF6; B = 8'h5E; #100;
A = 8'hF6; B = 8'h5F; #100;
A = 8'hF6; B = 8'h60; #100;
A = 8'hF6; B = 8'h61; #100;
A = 8'hF6; B = 8'h62; #100;
A = 8'hF6; B = 8'h63; #100;
A = 8'hF6; B = 8'h64; #100;
A = 8'hF6; B = 8'h65; #100;
A = 8'hF6; B = 8'h66; #100;
A = 8'hF6; B = 8'h67; #100;
A = 8'hF6; B = 8'h68; #100;
A = 8'hF6; B = 8'h69; #100;
A = 8'hF6; B = 8'h6A; #100;
A = 8'hF6; B = 8'h6B; #100;
A = 8'hF6; B = 8'h6C; #100;
A = 8'hF6; B = 8'h6D; #100;
A = 8'hF6; B = 8'h6E; #100;
A = 8'hF6; B = 8'h6F; #100;
A = 8'hF6; B = 8'h70; #100;
A = 8'hF6; B = 8'h71; #100;
A = 8'hF6; B = 8'h72; #100;
A = 8'hF6; B = 8'h73; #100;
A = 8'hF6; B = 8'h74; #100;
A = 8'hF6; B = 8'h75; #100;
A = 8'hF6; B = 8'h76; #100;
A = 8'hF6; B = 8'h77; #100;
A = 8'hF6; B = 8'h78; #100;
A = 8'hF6; B = 8'h79; #100;
A = 8'hF6; B = 8'h7A; #100;
A = 8'hF6; B = 8'h7B; #100;
A = 8'hF6; B = 8'h7C; #100;
A = 8'hF6; B = 8'h7D; #100;
A = 8'hF6; B = 8'h7E; #100;
A = 8'hF6; B = 8'h7F; #100;
A = 8'hF6; B = 8'h80; #100;
A = 8'hF6; B = 8'h81; #100;
A = 8'hF6; B = 8'h82; #100;
A = 8'hF6; B = 8'h83; #100;
A = 8'hF6; B = 8'h84; #100;
A = 8'hF6; B = 8'h85; #100;
A = 8'hF6; B = 8'h86; #100;
A = 8'hF6; B = 8'h87; #100;
A = 8'hF6; B = 8'h88; #100;
A = 8'hF6; B = 8'h89; #100;
A = 8'hF6; B = 8'h8A; #100;
A = 8'hF6; B = 8'h8B; #100;
A = 8'hF6; B = 8'h8C; #100;
A = 8'hF6; B = 8'h8D; #100;
A = 8'hF6; B = 8'h8E; #100;
A = 8'hF6; B = 8'h8F; #100;
A = 8'hF6; B = 8'h90; #100;
A = 8'hF6; B = 8'h91; #100;
A = 8'hF6; B = 8'h92; #100;
A = 8'hF6; B = 8'h93; #100;
A = 8'hF6; B = 8'h94; #100;
A = 8'hF6; B = 8'h95; #100;
A = 8'hF6; B = 8'h96; #100;
A = 8'hF6; B = 8'h97; #100;
A = 8'hF6; B = 8'h98; #100;
A = 8'hF6; B = 8'h99; #100;
A = 8'hF6; B = 8'h9A; #100;
A = 8'hF6; B = 8'h9B; #100;
A = 8'hF6; B = 8'h9C; #100;
A = 8'hF6; B = 8'h9D; #100;
A = 8'hF6; B = 8'h9E; #100;
A = 8'hF6; B = 8'h9F; #100;
A = 8'hF6; B = 8'hA0; #100;
A = 8'hF6; B = 8'hA1; #100;
A = 8'hF6; B = 8'hA2; #100;
A = 8'hF6; B = 8'hA3; #100;
A = 8'hF6; B = 8'hA4; #100;
A = 8'hF6; B = 8'hA5; #100;
A = 8'hF6; B = 8'hA6; #100;
A = 8'hF6; B = 8'hA7; #100;
A = 8'hF6; B = 8'hA8; #100;
A = 8'hF6; B = 8'hA9; #100;
A = 8'hF6; B = 8'hAA; #100;
A = 8'hF6; B = 8'hAB; #100;
A = 8'hF6; B = 8'hAC; #100;
A = 8'hF6; B = 8'hAD; #100;
A = 8'hF6; B = 8'hAE; #100;
A = 8'hF6; B = 8'hAF; #100;
A = 8'hF6; B = 8'hB0; #100;
A = 8'hF6; B = 8'hB1; #100;
A = 8'hF6; B = 8'hB2; #100;
A = 8'hF6; B = 8'hB3; #100;
A = 8'hF6; B = 8'hB4; #100;
A = 8'hF6; B = 8'hB5; #100;
A = 8'hF6; B = 8'hB6; #100;
A = 8'hF6; B = 8'hB7; #100;
A = 8'hF6; B = 8'hB8; #100;
A = 8'hF6; B = 8'hB9; #100;
A = 8'hF6; B = 8'hBA; #100;
A = 8'hF6; B = 8'hBB; #100;
A = 8'hF6; B = 8'hBC; #100;
A = 8'hF6; B = 8'hBD; #100;
A = 8'hF6; B = 8'hBE; #100;
A = 8'hF6; B = 8'hBF; #100;
A = 8'hF6; B = 8'hC0; #100;
A = 8'hF6; B = 8'hC1; #100;
A = 8'hF6; B = 8'hC2; #100;
A = 8'hF6; B = 8'hC3; #100;
A = 8'hF6; B = 8'hC4; #100;
A = 8'hF6; B = 8'hC5; #100;
A = 8'hF6; B = 8'hC6; #100;
A = 8'hF6; B = 8'hC7; #100;
A = 8'hF6; B = 8'hC8; #100;
A = 8'hF6; B = 8'hC9; #100;
A = 8'hF6; B = 8'hCA; #100;
A = 8'hF6; B = 8'hCB; #100;
A = 8'hF6; B = 8'hCC; #100;
A = 8'hF6; B = 8'hCD; #100;
A = 8'hF6; B = 8'hCE; #100;
A = 8'hF6; B = 8'hCF; #100;
A = 8'hF6; B = 8'hD0; #100;
A = 8'hF6; B = 8'hD1; #100;
A = 8'hF6; B = 8'hD2; #100;
A = 8'hF6; B = 8'hD3; #100;
A = 8'hF6; B = 8'hD4; #100;
A = 8'hF6; B = 8'hD5; #100;
A = 8'hF6; B = 8'hD6; #100;
A = 8'hF6; B = 8'hD7; #100;
A = 8'hF6; B = 8'hD8; #100;
A = 8'hF6; B = 8'hD9; #100;
A = 8'hF6; B = 8'hDA; #100;
A = 8'hF6; B = 8'hDB; #100;
A = 8'hF6; B = 8'hDC; #100;
A = 8'hF6; B = 8'hDD; #100;
A = 8'hF6; B = 8'hDE; #100;
A = 8'hF6; B = 8'hDF; #100;
A = 8'hF6; B = 8'hE0; #100;
A = 8'hF6; B = 8'hE1; #100;
A = 8'hF6; B = 8'hE2; #100;
A = 8'hF6; B = 8'hE3; #100;
A = 8'hF6; B = 8'hE4; #100;
A = 8'hF6; B = 8'hE5; #100;
A = 8'hF6; B = 8'hE6; #100;
A = 8'hF6; B = 8'hE7; #100;
A = 8'hF6; B = 8'hE8; #100;
A = 8'hF6; B = 8'hE9; #100;
A = 8'hF6; B = 8'hEA; #100;
A = 8'hF6; B = 8'hEB; #100;
A = 8'hF6; B = 8'hEC; #100;
A = 8'hF6; B = 8'hED; #100;
A = 8'hF6; B = 8'hEE; #100;
A = 8'hF6; B = 8'hEF; #100;
A = 8'hF6; B = 8'hF0; #100;
A = 8'hF6; B = 8'hF1; #100;
A = 8'hF6; B = 8'hF2; #100;
A = 8'hF6; B = 8'hF3; #100;
A = 8'hF6; B = 8'hF4; #100;
A = 8'hF6; B = 8'hF5; #100;
A = 8'hF6; B = 8'hF6; #100;
A = 8'hF6; B = 8'hF7; #100;
A = 8'hF6; B = 8'hF8; #100;
A = 8'hF6; B = 8'hF9; #100;
A = 8'hF6; B = 8'hFA; #100;
A = 8'hF6; B = 8'hFB; #100;
A = 8'hF6; B = 8'hFC; #100;
A = 8'hF6; B = 8'hFD; #100;
A = 8'hF6; B = 8'hFE; #100;
A = 8'hF6; B = 8'hFF; #100;
A = 8'hF7; B = 8'h0; #100;
A = 8'hF7; B = 8'h1; #100;
A = 8'hF7; B = 8'h2; #100;
A = 8'hF7; B = 8'h3; #100;
A = 8'hF7; B = 8'h4; #100;
A = 8'hF7; B = 8'h5; #100;
A = 8'hF7; B = 8'h6; #100;
A = 8'hF7; B = 8'h7; #100;
A = 8'hF7; B = 8'h8; #100;
A = 8'hF7; B = 8'h9; #100;
A = 8'hF7; B = 8'hA; #100;
A = 8'hF7; B = 8'hB; #100;
A = 8'hF7; B = 8'hC; #100;
A = 8'hF7; B = 8'hD; #100;
A = 8'hF7; B = 8'hE; #100;
A = 8'hF7; B = 8'hF; #100;
A = 8'hF7; B = 8'h10; #100;
A = 8'hF7; B = 8'h11; #100;
A = 8'hF7; B = 8'h12; #100;
A = 8'hF7; B = 8'h13; #100;
A = 8'hF7; B = 8'h14; #100;
A = 8'hF7; B = 8'h15; #100;
A = 8'hF7; B = 8'h16; #100;
A = 8'hF7; B = 8'h17; #100;
A = 8'hF7; B = 8'h18; #100;
A = 8'hF7; B = 8'h19; #100;
A = 8'hF7; B = 8'h1A; #100;
A = 8'hF7; B = 8'h1B; #100;
A = 8'hF7; B = 8'h1C; #100;
A = 8'hF7; B = 8'h1D; #100;
A = 8'hF7; B = 8'h1E; #100;
A = 8'hF7; B = 8'h1F; #100;
A = 8'hF7; B = 8'h20; #100;
A = 8'hF7; B = 8'h21; #100;
A = 8'hF7; B = 8'h22; #100;
A = 8'hF7; B = 8'h23; #100;
A = 8'hF7; B = 8'h24; #100;
A = 8'hF7; B = 8'h25; #100;
A = 8'hF7; B = 8'h26; #100;
A = 8'hF7; B = 8'h27; #100;
A = 8'hF7; B = 8'h28; #100;
A = 8'hF7; B = 8'h29; #100;
A = 8'hF7; B = 8'h2A; #100;
A = 8'hF7; B = 8'h2B; #100;
A = 8'hF7; B = 8'h2C; #100;
A = 8'hF7; B = 8'h2D; #100;
A = 8'hF7; B = 8'h2E; #100;
A = 8'hF7; B = 8'h2F; #100;
A = 8'hF7; B = 8'h30; #100;
A = 8'hF7; B = 8'h31; #100;
A = 8'hF7; B = 8'h32; #100;
A = 8'hF7; B = 8'h33; #100;
A = 8'hF7; B = 8'h34; #100;
A = 8'hF7; B = 8'h35; #100;
A = 8'hF7; B = 8'h36; #100;
A = 8'hF7; B = 8'h37; #100;
A = 8'hF7; B = 8'h38; #100;
A = 8'hF7; B = 8'h39; #100;
A = 8'hF7; B = 8'h3A; #100;
A = 8'hF7; B = 8'h3B; #100;
A = 8'hF7; B = 8'h3C; #100;
A = 8'hF7; B = 8'h3D; #100;
A = 8'hF7; B = 8'h3E; #100;
A = 8'hF7; B = 8'h3F; #100;
A = 8'hF7; B = 8'h40; #100;
A = 8'hF7; B = 8'h41; #100;
A = 8'hF7; B = 8'h42; #100;
A = 8'hF7; B = 8'h43; #100;
A = 8'hF7; B = 8'h44; #100;
A = 8'hF7; B = 8'h45; #100;
A = 8'hF7; B = 8'h46; #100;
A = 8'hF7; B = 8'h47; #100;
A = 8'hF7; B = 8'h48; #100;
A = 8'hF7; B = 8'h49; #100;
A = 8'hF7; B = 8'h4A; #100;
A = 8'hF7; B = 8'h4B; #100;
A = 8'hF7; B = 8'h4C; #100;
A = 8'hF7; B = 8'h4D; #100;
A = 8'hF7; B = 8'h4E; #100;
A = 8'hF7; B = 8'h4F; #100;
A = 8'hF7; B = 8'h50; #100;
A = 8'hF7; B = 8'h51; #100;
A = 8'hF7; B = 8'h52; #100;
A = 8'hF7; B = 8'h53; #100;
A = 8'hF7; B = 8'h54; #100;
A = 8'hF7; B = 8'h55; #100;
A = 8'hF7; B = 8'h56; #100;
A = 8'hF7; B = 8'h57; #100;
A = 8'hF7; B = 8'h58; #100;
A = 8'hF7; B = 8'h59; #100;
A = 8'hF7; B = 8'h5A; #100;
A = 8'hF7; B = 8'h5B; #100;
A = 8'hF7; B = 8'h5C; #100;
A = 8'hF7; B = 8'h5D; #100;
A = 8'hF7; B = 8'h5E; #100;
A = 8'hF7; B = 8'h5F; #100;
A = 8'hF7; B = 8'h60; #100;
A = 8'hF7; B = 8'h61; #100;
A = 8'hF7; B = 8'h62; #100;
A = 8'hF7; B = 8'h63; #100;
A = 8'hF7; B = 8'h64; #100;
A = 8'hF7; B = 8'h65; #100;
A = 8'hF7; B = 8'h66; #100;
A = 8'hF7; B = 8'h67; #100;
A = 8'hF7; B = 8'h68; #100;
A = 8'hF7; B = 8'h69; #100;
A = 8'hF7; B = 8'h6A; #100;
A = 8'hF7; B = 8'h6B; #100;
A = 8'hF7; B = 8'h6C; #100;
A = 8'hF7; B = 8'h6D; #100;
A = 8'hF7; B = 8'h6E; #100;
A = 8'hF7; B = 8'h6F; #100;
A = 8'hF7; B = 8'h70; #100;
A = 8'hF7; B = 8'h71; #100;
A = 8'hF7; B = 8'h72; #100;
A = 8'hF7; B = 8'h73; #100;
A = 8'hF7; B = 8'h74; #100;
A = 8'hF7; B = 8'h75; #100;
A = 8'hF7; B = 8'h76; #100;
A = 8'hF7; B = 8'h77; #100;
A = 8'hF7; B = 8'h78; #100;
A = 8'hF7; B = 8'h79; #100;
A = 8'hF7; B = 8'h7A; #100;
A = 8'hF7; B = 8'h7B; #100;
A = 8'hF7; B = 8'h7C; #100;
A = 8'hF7; B = 8'h7D; #100;
A = 8'hF7; B = 8'h7E; #100;
A = 8'hF7; B = 8'h7F; #100;
A = 8'hF7; B = 8'h80; #100;
A = 8'hF7; B = 8'h81; #100;
A = 8'hF7; B = 8'h82; #100;
A = 8'hF7; B = 8'h83; #100;
A = 8'hF7; B = 8'h84; #100;
A = 8'hF7; B = 8'h85; #100;
A = 8'hF7; B = 8'h86; #100;
A = 8'hF7; B = 8'h87; #100;
A = 8'hF7; B = 8'h88; #100;
A = 8'hF7; B = 8'h89; #100;
A = 8'hF7; B = 8'h8A; #100;
A = 8'hF7; B = 8'h8B; #100;
A = 8'hF7; B = 8'h8C; #100;
A = 8'hF7; B = 8'h8D; #100;
A = 8'hF7; B = 8'h8E; #100;
A = 8'hF7; B = 8'h8F; #100;
A = 8'hF7; B = 8'h90; #100;
A = 8'hF7; B = 8'h91; #100;
A = 8'hF7; B = 8'h92; #100;
A = 8'hF7; B = 8'h93; #100;
A = 8'hF7; B = 8'h94; #100;
A = 8'hF7; B = 8'h95; #100;
A = 8'hF7; B = 8'h96; #100;
A = 8'hF7; B = 8'h97; #100;
A = 8'hF7; B = 8'h98; #100;
A = 8'hF7; B = 8'h99; #100;
A = 8'hF7; B = 8'h9A; #100;
A = 8'hF7; B = 8'h9B; #100;
A = 8'hF7; B = 8'h9C; #100;
A = 8'hF7; B = 8'h9D; #100;
A = 8'hF7; B = 8'h9E; #100;
A = 8'hF7; B = 8'h9F; #100;
A = 8'hF7; B = 8'hA0; #100;
A = 8'hF7; B = 8'hA1; #100;
A = 8'hF7; B = 8'hA2; #100;
A = 8'hF7; B = 8'hA3; #100;
A = 8'hF7; B = 8'hA4; #100;
A = 8'hF7; B = 8'hA5; #100;
A = 8'hF7; B = 8'hA6; #100;
A = 8'hF7; B = 8'hA7; #100;
A = 8'hF7; B = 8'hA8; #100;
A = 8'hF7; B = 8'hA9; #100;
A = 8'hF7; B = 8'hAA; #100;
A = 8'hF7; B = 8'hAB; #100;
A = 8'hF7; B = 8'hAC; #100;
A = 8'hF7; B = 8'hAD; #100;
A = 8'hF7; B = 8'hAE; #100;
A = 8'hF7; B = 8'hAF; #100;
A = 8'hF7; B = 8'hB0; #100;
A = 8'hF7; B = 8'hB1; #100;
A = 8'hF7; B = 8'hB2; #100;
A = 8'hF7; B = 8'hB3; #100;
A = 8'hF7; B = 8'hB4; #100;
A = 8'hF7; B = 8'hB5; #100;
A = 8'hF7; B = 8'hB6; #100;
A = 8'hF7; B = 8'hB7; #100;
A = 8'hF7; B = 8'hB8; #100;
A = 8'hF7; B = 8'hB9; #100;
A = 8'hF7; B = 8'hBA; #100;
A = 8'hF7; B = 8'hBB; #100;
A = 8'hF7; B = 8'hBC; #100;
A = 8'hF7; B = 8'hBD; #100;
A = 8'hF7; B = 8'hBE; #100;
A = 8'hF7; B = 8'hBF; #100;
A = 8'hF7; B = 8'hC0; #100;
A = 8'hF7; B = 8'hC1; #100;
A = 8'hF7; B = 8'hC2; #100;
A = 8'hF7; B = 8'hC3; #100;
A = 8'hF7; B = 8'hC4; #100;
A = 8'hF7; B = 8'hC5; #100;
A = 8'hF7; B = 8'hC6; #100;
A = 8'hF7; B = 8'hC7; #100;
A = 8'hF7; B = 8'hC8; #100;
A = 8'hF7; B = 8'hC9; #100;
A = 8'hF7; B = 8'hCA; #100;
A = 8'hF7; B = 8'hCB; #100;
A = 8'hF7; B = 8'hCC; #100;
A = 8'hF7; B = 8'hCD; #100;
A = 8'hF7; B = 8'hCE; #100;
A = 8'hF7; B = 8'hCF; #100;
A = 8'hF7; B = 8'hD0; #100;
A = 8'hF7; B = 8'hD1; #100;
A = 8'hF7; B = 8'hD2; #100;
A = 8'hF7; B = 8'hD3; #100;
A = 8'hF7; B = 8'hD4; #100;
A = 8'hF7; B = 8'hD5; #100;
A = 8'hF7; B = 8'hD6; #100;
A = 8'hF7; B = 8'hD7; #100;
A = 8'hF7; B = 8'hD8; #100;
A = 8'hF7; B = 8'hD9; #100;
A = 8'hF7; B = 8'hDA; #100;
A = 8'hF7; B = 8'hDB; #100;
A = 8'hF7; B = 8'hDC; #100;
A = 8'hF7; B = 8'hDD; #100;
A = 8'hF7; B = 8'hDE; #100;
A = 8'hF7; B = 8'hDF; #100;
A = 8'hF7; B = 8'hE0; #100;
A = 8'hF7; B = 8'hE1; #100;
A = 8'hF7; B = 8'hE2; #100;
A = 8'hF7; B = 8'hE3; #100;
A = 8'hF7; B = 8'hE4; #100;
A = 8'hF7; B = 8'hE5; #100;
A = 8'hF7; B = 8'hE6; #100;
A = 8'hF7; B = 8'hE7; #100;
A = 8'hF7; B = 8'hE8; #100;
A = 8'hF7; B = 8'hE9; #100;
A = 8'hF7; B = 8'hEA; #100;
A = 8'hF7; B = 8'hEB; #100;
A = 8'hF7; B = 8'hEC; #100;
A = 8'hF7; B = 8'hED; #100;
A = 8'hF7; B = 8'hEE; #100;
A = 8'hF7; B = 8'hEF; #100;
A = 8'hF7; B = 8'hF0; #100;
A = 8'hF7; B = 8'hF1; #100;
A = 8'hF7; B = 8'hF2; #100;
A = 8'hF7; B = 8'hF3; #100;
A = 8'hF7; B = 8'hF4; #100;
A = 8'hF7; B = 8'hF5; #100;
A = 8'hF7; B = 8'hF6; #100;
A = 8'hF7; B = 8'hF7; #100;
A = 8'hF7; B = 8'hF8; #100;
A = 8'hF7; B = 8'hF9; #100;
A = 8'hF7; B = 8'hFA; #100;
A = 8'hF7; B = 8'hFB; #100;
A = 8'hF7; B = 8'hFC; #100;
A = 8'hF7; B = 8'hFD; #100;
A = 8'hF7; B = 8'hFE; #100;
A = 8'hF7; B = 8'hFF; #100;
A = 8'hF8; B = 8'h0; #100;
A = 8'hF8; B = 8'h1; #100;
A = 8'hF8; B = 8'h2; #100;
A = 8'hF8; B = 8'h3; #100;
A = 8'hF8; B = 8'h4; #100;
A = 8'hF8; B = 8'h5; #100;
A = 8'hF8; B = 8'h6; #100;
A = 8'hF8; B = 8'h7; #100;
A = 8'hF8; B = 8'h8; #100;
A = 8'hF8; B = 8'h9; #100;
A = 8'hF8; B = 8'hA; #100;
A = 8'hF8; B = 8'hB; #100;
A = 8'hF8; B = 8'hC; #100;
A = 8'hF8; B = 8'hD; #100;
A = 8'hF8; B = 8'hE; #100;
A = 8'hF8; B = 8'hF; #100;
A = 8'hF8; B = 8'h10; #100;
A = 8'hF8; B = 8'h11; #100;
A = 8'hF8; B = 8'h12; #100;
A = 8'hF8; B = 8'h13; #100;
A = 8'hF8; B = 8'h14; #100;
A = 8'hF8; B = 8'h15; #100;
A = 8'hF8; B = 8'h16; #100;
A = 8'hF8; B = 8'h17; #100;
A = 8'hF8; B = 8'h18; #100;
A = 8'hF8; B = 8'h19; #100;
A = 8'hF8; B = 8'h1A; #100;
A = 8'hF8; B = 8'h1B; #100;
A = 8'hF8; B = 8'h1C; #100;
A = 8'hF8; B = 8'h1D; #100;
A = 8'hF8; B = 8'h1E; #100;
A = 8'hF8; B = 8'h1F; #100;
A = 8'hF8; B = 8'h20; #100;
A = 8'hF8; B = 8'h21; #100;
A = 8'hF8; B = 8'h22; #100;
A = 8'hF8; B = 8'h23; #100;
A = 8'hF8; B = 8'h24; #100;
A = 8'hF8; B = 8'h25; #100;
A = 8'hF8; B = 8'h26; #100;
A = 8'hF8; B = 8'h27; #100;
A = 8'hF8; B = 8'h28; #100;
A = 8'hF8; B = 8'h29; #100;
A = 8'hF8; B = 8'h2A; #100;
A = 8'hF8; B = 8'h2B; #100;
A = 8'hF8; B = 8'h2C; #100;
A = 8'hF8; B = 8'h2D; #100;
A = 8'hF8; B = 8'h2E; #100;
A = 8'hF8; B = 8'h2F; #100;
A = 8'hF8; B = 8'h30; #100;
A = 8'hF8; B = 8'h31; #100;
A = 8'hF8; B = 8'h32; #100;
A = 8'hF8; B = 8'h33; #100;
A = 8'hF8; B = 8'h34; #100;
A = 8'hF8; B = 8'h35; #100;
A = 8'hF8; B = 8'h36; #100;
A = 8'hF8; B = 8'h37; #100;
A = 8'hF8; B = 8'h38; #100;
A = 8'hF8; B = 8'h39; #100;
A = 8'hF8; B = 8'h3A; #100;
A = 8'hF8; B = 8'h3B; #100;
A = 8'hF8; B = 8'h3C; #100;
A = 8'hF8; B = 8'h3D; #100;
A = 8'hF8; B = 8'h3E; #100;
A = 8'hF8; B = 8'h3F; #100;
A = 8'hF8; B = 8'h40; #100;
A = 8'hF8; B = 8'h41; #100;
A = 8'hF8; B = 8'h42; #100;
A = 8'hF8; B = 8'h43; #100;
A = 8'hF8; B = 8'h44; #100;
A = 8'hF8; B = 8'h45; #100;
A = 8'hF8; B = 8'h46; #100;
A = 8'hF8; B = 8'h47; #100;
A = 8'hF8; B = 8'h48; #100;
A = 8'hF8; B = 8'h49; #100;
A = 8'hF8; B = 8'h4A; #100;
A = 8'hF8; B = 8'h4B; #100;
A = 8'hF8; B = 8'h4C; #100;
A = 8'hF8; B = 8'h4D; #100;
A = 8'hF8; B = 8'h4E; #100;
A = 8'hF8; B = 8'h4F; #100;
A = 8'hF8; B = 8'h50; #100;
A = 8'hF8; B = 8'h51; #100;
A = 8'hF8; B = 8'h52; #100;
A = 8'hF8; B = 8'h53; #100;
A = 8'hF8; B = 8'h54; #100;
A = 8'hF8; B = 8'h55; #100;
A = 8'hF8; B = 8'h56; #100;
A = 8'hF8; B = 8'h57; #100;
A = 8'hF8; B = 8'h58; #100;
A = 8'hF8; B = 8'h59; #100;
A = 8'hF8; B = 8'h5A; #100;
A = 8'hF8; B = 8'h5B; #100;
A = 8'hF8; B = 8'h5C; #100;
A = 8'hF8; B = 8'h5D; #100;
A = 8'hF8; B = 8'h5E; #100;
A = 8'hF8; B = 8'h5F; #100;
A = 8'hF8; B = 8'h60; #100;
A = 8'hF8; B = 8'h61; #100;
A = 8'hF8; B = 8'h62; #100;
A = 8'hF8; B = 8'h63; #100;
A = 8'hF8; B = 8'h64; #100;
A = 8'hF8; B = 8'h65; #100;
A = 8'hF8; B = 8'h66; #100;
A = 8'hF8; B = 8'h67; #100;
A = 8'hF8; B = 8'h68; #100;
A = 8'hF8; B = 8'h69; #100;
A = 8'hF8; B = 8'h6A; #100;
A = 8'hF8; B = 8'h6B; #100;
A = 8'hF8; B = 8'h6C; #100;
A = 8'hF8; B = 8'h6D; #100;
A = 8'hF8; B = 8'h6E; #100;
A = 8'hF8; B = 8'h6F; #100;
A = 8'hF8; B = 8'h70; #100;
A = 8'hF8; B = 8'h71; #100;
A = 8'hF8; B = 8'h72; #100;
A = 8'hF8; B = 8'h73; #100;
A = 8'hF8; B = 8'h74; #100;
A = 8'hF8; B = 8'h75; #100;
A = 8'hF8; B = 8'h76; #100;
A = 8'hF8; B = 8'h77; #100;
A = 8'hF8; B = 8'h78; #100;
A = 8'hF8; B = 8'h79; #100;
A = 8'hF8; B = 8'h7A; #100;
A = 8'hF8; B = 8'h7B; #100;
A = 8'hF8; B = 8'h7C; #100;
A = 8'hF8; B = 8'h7D; #100;
A = 8'hF8; B = 8'h7E; #100;
A = 8'hF8; B = 8'h7F; #100;
A = 8'hF8; B = 8'h80; #100;
A = 8'hF8; B = 8'h81; #100;
A = 8'hF8; B = 8'h82; #100;
A = 8'hF8; B = 8'h83; #100;
A = 8'hF8; B = 8'h84; #100;
A = 8'hF8; B = 8'h85; #100;
A = 8'hF8; B = 8'h86; #100;
A = 8'hF8; B = 8'h87; #100;
A = 8'hF8; B = 8'h88; #100;
A = 8'hF8; B = 8'h89; #100;
A = 8'hF8; B = 8'h8A; #100;
A = 8'hF8; B = 8'h8B; #100;
A = 8'hF8; B = 8'h8C; #100;
A = 8'hF8; B = 8'h8D; #100;
A = 8'hF8; B = 8'h8E; #100;
A = 8'hF8; B = 8'h8F; #100;
A = 8'hF8; B = 8'h90; #100;
A = 8'hF8; B = 8'h91; #100;
A = 8'hF8; B = 8'h92; #100;
A = 8'hF8; B = 8'h93; #100;
A = 8'hF8; B = 8'h94; #100;
A = 8'hF8; B = 8'h95; #100;
A = 8'hF8; B = 8'h96; #100;
A = 8'hF8; B = 8'h97; #100;
A = 8'hF8; B = 8'h98; #100;
A = 8'hF8; B = 8'h99; #100;
A = 8'hF8; B = 8'h9A; #100;
A = 8'hF8; B = 8'h9B; #100;
A = 8'hF8; B = 8'h9C; #100;
A = 8'hF8; B = 8'h9D; #100;
A = 8'hF8; B = 8'h9E; #100;
A = 8'hF8; B = 8'h9F; #100;
A = 8'hF8; B = 8'hA0; #100;
A = 8'hF8; B = 8'hA1; #100;
A = 8'hF8; B = 8'hA2; #100;
A = 8'hF8; B = 8'hA3; #100;
A = 8'hF8; B = 8'hA4; #100;
A = 8'hF8; B = 8'hA5; #100;
A = 8'hF8; B = 8'hA6; #100;
A = 8'hF8; B = 8'hA7; #100;
A = 8'hF8; B = 8'hA8; #100;
A = 8'hF8; B = 8'hA9; #100;
A = 8'hF8; B = 8'hAA; #100;
A = 8'hF8; B = 8'hAB; #100;
A = 8'hF8; B = 8'hAC; #100;
A = 8'hF8; B = 8'hAD; #100;
A = 8'hF8; B = 8'hAE; #100;
A = 8'hF8; B = 8'hAF; #100;
A = 8'hF8; B = 8'hB0; #100;
A = 8'hF8; B = 8'hB1; #100;
A = 8'hF8; B = 8'hB2; #100;
A = 8'hF8; B = 8'hB3; #100;
A = 8'hF8; B = 8'hB4; #100;
A = 8'hF8; B = 8'hB5; #100;
A = 8'hF8; B = 8'hB6; #100;
A = 8'hF8; B = 8'hB7; #100;
A = 8'hF8; B = 8'hB8; #100;
A = 8'hF8; B = 8'hB9; #100;
A = 8'hF8; B = 8'hBA; #100;
A = 8'hF8; B = 8'hBB; #100;
A = 8'hF8; B = 8'hBC; #100;
A = 8'hF8; B = 8'hBD; #100;
A = 8'hF8; B = 8'hBE; #100;
A = 8'hF8; B = 8'hBF; #100;
A = 8'hF8; B = 8'hC0; #100;
A = 8'hF8; B = 8'hC1; #100;
A = 8'hF8; B = 8'hC2; #100;
A = 8'hF8; B = 8'hC3; #100;
A = 8'hF8; B = 8'hC4; #100;
A = 8'hF8; B = 8'hC5; #100;
A = 8'hF8; B = 8'hC6; #100;
A = 8'hF8; B = 8'hC7; #100;
A = 8'hF8; B = 8'hC8; #100;
A = 8'hF8; B = 8'hC9; #100;
A = 8'hF8; B = 8'hCA; #100;
A = 8'hF8; B = 8'hCB; #100;
A = 8'hF8; B = 8'hCC; #100;
A = 8'hF8; B = 8'hCD; #100;
A = 8'hF8; B = 8'hCE; #100;
A = 8'hF8; B = 8'hCF; #100;
A = 8'hF8; B = 8'hD0; #100;
A = 8'hF8; B = 8'hD1; #100;
A = 8'hF8; B = 8'hD2; #100;
A = 8'hF8; B = 8'hD3; #100;
A = 8'hF8; B = 8'hD4; #100;
A = 8'hF8; B = 8'hD5; #100;
A = 8'hF8; B = 8'hD6; #100;
A = 8'hF8; B = 8'hD7; #100;
A = 8'hF8; B = 8'hD8; #100;
A = 8'hF8; B = 8'hD9; #100;
A = 8'hF8; B = 8'hDA; #100;
A = 8'hF8; B = 8'hDB; #100;
A = 8'hF8; B = 8'hDC; #100;
A = 8'hF8; B = 8'hDD; #100;
A = 8'hF8; B = 8'hDE; #100;
A = 8'hF8; B = 8'hDF; #100;
A = 8'hF8; B = 8'hE0; #100;
A = 8'hF8; B = 8'hE1; #100;
A = 8'hF8; B = 8'hE2; #100;
A = 8'hF8; B = 8'hE3; #100;
A = 8'hF8; B = 8'hE4; #100;
A = 8'hF8; B = 8'hE5; #100;
A = 8'hF8; B = 8'hE6; #100;
A = 8'hF8; B = 8'hE7; #100;
A = 8'hF8; B = 8'hE8; #100;
A = 8'hF8; B = 8'hE9; #100;
A = 8'hF8; B = 8'hEA; #100;
A = 8'hF8; B = 8'hEB; #100;
A = 8'hF8; B = 8'hEC; #100;
A = 8'hF8; B = 8'hED; #100;
A = 8'hF8; B = 8'hEE; #100;
A = 8'hF8; B = 8'hEF; #100;
A = 8'hF8; B = 8'hF0; #100;
A = 8'hF8; B = 8'hF1; #100;
A = 8'hF8; B = 8'hF2; #100;
A = 8'hF8; B = 8'hF3; #100;
A = 8'hF8; B = 8'hF4; #100;
A = 8'hF8; B = 8'hF5; #100;
A = 8'hF8; B = 8'hF6; #100;
A = 8'hF8; B = 8'hF7; #100;
A = 8'hF8; B = 8'hF8; #100;
A = 8'hF8; B = 8'hF9; #100;
A = 8'hF8; B = 8'hFA; #100;
A = 8'hF8; B = 8'hFB; #100;
A = 8'hF8; B = 8'hFC; #100;
A = 8'hF8; B = 8'hFD; #100;
A = 8'hF8; B = 8'hFE; #100;
A = 8'hF8; B = 8'hFF; #100;
A = 8'hF9; B = 8'h0; #100;
A = 8'hF9; B = 8'h1; #100;
A = 8'hF9; B = 8'h2; #100;
A = 8'hF9; B = 8'h3; #100;
A = 8'hF9; B = 8'h4; #100;
A = 8'hF9; B = 8'h5; #100;
A = 8'hF9; B = 8'h6; #100;
A = 8'hF9; B = 8'h7; #100;
A = 8'hF9; B = 8'h8; #100;
A = 8'hF9; B = 8'h9; #100;
A = 8'hF9; B = 8'hA; #100;
A = 8'hF9; B = 8'hB; #100;
A = 8'hF9; B = 8'hC; #100;
A = 8'hF9; B = 8'hD; #100;
A = 8'hF9; B = 8'hE; #100;
A = 8'hF9; B = 8'hF; #100;
A = 8'hF9; B = 8'h10; #100;
A = 8'hF9; B = 8'h11; #100;
A = 8'hF9; B = 8'h12; #100;
A = 8'hF9; B = 8'h13; #100;
A = 8'hF9; B = 8'h14; #100;
A = 8'hF9; B = 8'h15; #100;
A = 8'hF9; B = 8'h16; #100;
A = 8'hF9; B = 8'h17; #100;
A = 8'hF9; B = 8'h18; #100;
A = 8'hF9; B = 8'h19; #100;
A = 8'hF9; B = 8'h1A; #100;
A = 8'hF9; B = 8'h1B; #100;
A = 8'hF9; B = 8'h1C; #100;
A = 8'hF9; B = 8'h1D; #100;
A = 8'hF9; B = 8'h1E; #100;
A = 8'hF9; B = 8'h1F; #100;
A = 8'hF9; B = 8'h20; #100;
A = 8'hF9; B = 8'h21; #100;
A = 8'hF9; B = 8'h22; #100;
A = 8'hF9; B = 8'h23; #100;
A = 8'hF9; B = 8'h24; #100;
A = 8'hF9; B = 8'h25; #100;
A = 8'hF9; B = 8'h26; #100;
A = 8'hF9; B = 8'h27; #100;
A = 8'hF9; B = 8'h28; #100;
A = 8'hF9; B = 8'h29; #100;
A = 8'hF9; B = 8'h2A; #100;
A = 8'hF9; B = 8'h2B; #100;
A = 8'hF9; B = 8'h2C; #100;
A = 8'hF9; B = 8'h2D; #100;
A = 8'hF9; B = 8'h2E; #100;
A = 8'hF9; B = 8'h2F; #100;
A = 8'hF9; B = 8'h30; #100;
A = 8'hF9; B = 8'h31; #100;
A = 8'hF9; B = 8'h32; #100;
A = 8'hF9; B = 8'h33; #100;
A = 8'hF9; B = 8'h34; #100;
A = 8'hF9; B = 8'h35; #100;
A = 8'hF9; B = 8'h36; #100;
A = 8'hF9; B = 8'h37; #100;
A = 8'hF9; B = 8'h38; #100;
A = 8'hF9; B = 8'h39; #100;
A = 8'hF9; B = 8'h3A; #100;
A = 8'hF9; B = 8'h3B; #100;
A = 8'hF9; B = 8'h3C; #100;
A = 8'hF9; B = 8'h3D; #100;
A = 8'hF9; B = 8'h3E; #100;
A = 8'hF9; B = 8'h3F; #100;
A = 8'hF9; B = 8'h40; #100;
A = 8'hF9; B = 8'h41; #100;
A = 8'hF9; B = 8'h42; #100;
A = 8'hF9; B = 8'h43; #100;
A = 8'hF9; B = 8'h44; #100;
A = 8'hF9; B = 8'h45; #100;
A = 8'hF9; B = 8'h46; #100;
A = 8'hF9; B = 8'h47; #100;
A = 8'hF9; B = 8'h48; #100;
A = 8'hF9; B = 8'h49; #100;
A = 8'hF9; B = 8'h4A; #100;
A = 8'hF9; B = 8'h4B; #100;
A = 8'hF9; B = 8'h4C; #100;
A = 8'hF9; B = 8'h4D; #100;
A = 8'hF9; B = 8'h4E; #100;
A = 8'hF9; B = 8'h4F; #100;
A = 8'hF9; B = 8'h50; #100;
A = 8'hF9; B = 8'h51; #100;
A = 8'hF9; B = 8'h52; #100;
A = 8'hF9; B = 8'h53; #100;
A = 8'hF9; B = 8'h54; #100;
A = 8'hF9; B = 8'h55; #100;
A = 8'hF9; B = 8'h56; #100;
A = 8'hF9; B = 8'h57; #100;
A = 8'hF9; B = 8'h58; #100;
A = 8'hF9; B = 8'h59; #100;
A = 8'hF9; B = 8'h5A; #100;
A = 8'hF9; B = 8'h5B; #100;
A = 8'hF9; B = 8'h5C; #100;
A = 8'hF9; B = 8'h5D; #100;
A = 8'hF9; B = 8'h5E; #100;
A = 8'hF9; B = 8'h5F; #100;
A = 8'hF9; B = 8'h60; #100;
A = 8'hF9; B = 8'h61; #100;
A = 8'hF9; B = 8'h62; #100;
A = 8'hF9; B = 8'h63; #100;
A = 8'hF9; B = 8'h64; #100;
A = 8'hF9; B = 8'h65; #100;
A = 8'hF9; B = 8'h66; #100;
A = 8'hF9; B = 8'h67; #100;
A = 8'hF9; B = 8'h68; #100;
A = 8'hF9; B = 8'h69; #100;
A = 8'hF9; B = 8'h6A; #100;
A = 8'hF9; B = 8'h6B; #100;
A = 8'hF9; B = 8'h6C; #100;
A = 8'hF9; B = 8'h6D; #100;
A = 8'hF9; B = 8'h6E; #100;
A = 8'hF9; B = 8'h6F; #100;
A = 8'hF9; B = 8'h70; #100;
A = 8'hF9; B = 8'h71; #100;
A = 8'hF9; B = 8'h72; #100;
A = 8'hF9; B = 8'h73; #100;
A = 8'hF9; B = 8'h74; #100;
A = 8'hF9; B = 8'h75; #100;
A = 8'hF9; B = 8'h76; #100;
A = 8'hF9; B = 8'h77; #100;
A = 8'hF9; B = 8'h78; #100;
A = 8'hF9; B = 8'h79; #100;
A = 8'hF9; B = 8'h7A; #100;
A = 8'hF9; B = 8'h7B; #100;
A = 8'hF9; B = 8'h7C; #100;
A = 8'hF9; B = 8'h7D; #100;
A = 8'hF9; B = 8'h7E; #100;
A = 8'hF9; B = 8'h7F; #100;
A = 8'hF9; B = 8'h80; #100;
A = 8'hF9; B = 8'h81; #100;
A = 8'hF9; B = 8'h82; #100;
A = 8'hF9; B = 8'h83; #100;
A = 8'hF9; B = 8'h84; #100;
A = 8'hF9; B = 8'h85; #100;
A = 8'hF9; B = 8'h86; #100;
A = 8'hF9; B = 8'h87; #100;
A = 8'hF9; B = 8'h88; #100;
A = 8'hF9; B = 8'h89; #100;
A = 8'hF9; B = 8'h8A; #100;
A = 8'hF9; B = 8'h8B; #100;
A = 8'hF9; B = 8'h8C; #100;
A = 8'hF9; B = 8'h8D; #100;
A = 8'hF9; B = 8'h8E; #100;
A = 8'hF9; B = 8'h8F; #100;
A = 8'hF9; B = 8'h90; #100;
A = 8'hF9; B = 8'h91; #100;
A = 8'hF9; B = 8'h92; #100;
A = 8'hF9; B = 8'h93; #100;
A = 8'hF9; B = 8'h94; #100;
A = 8'hF9; B = 8'h95; #100;
A = 8'hF9; B = 8'h96; #100;
A = 8'hF9; B = 8'h97; #100;
A = 8'hF9; B = 8'h98; #100;
A = 8'hF9; B = 8'h99; #100;
A = 8'hF9; B = 8'h9A; #100;
A = 8'hF9; B = 8'h9B; #100;
A = 8'hF9; B = 8'h9C; #100;
A = 8'hF9; B = 8'h9D; #100;
A = 8'hF9; B = 8'h9E; #100;
A = 8'hF9; B = 8'h9F; #100;
A = 8'hF9; B = 8'hA0; #100;
A = 8'hF9; B = 8'hA1; #100;
A = 8'hF9; B = 8'hA2; #100;
A = 8'hF9; B = 8'hA3; #100;
A = 8'hF9; B = 8'hA4; #100;
A = 8'hF9; B = 8'hA5; #100;
A = 8'hF9; B = 8'hA6; #100;
A = 8'hF9; B = 8'hA7; #100;
A = 8'hF9; B = 8'hA8; #100;
A = 8'hF9; B = 8'hA9; #100;
A = 8'hF9; B = 8'hAA; #100;
A = 8'hF9; B = 8'hAB; #100;
A = 8'hF9; B = 8'hAC; #100;
A = 8'hF9; B = 8'hAD; #100;
A = 8'hF9; B = 8'hAE; #100;
A = 8'hF9; B = 8'hAF; #100;
A = 8'hF9; B = 8'hB0; #100;
A = 8'hF9; B = 8'hB1; #100;
A = 8'hF9; B = 8'hB2; #100;
A = 8'hF9; B = 8'hB3; #100;
A = 8'hF9; B = 8'hB4; #100;
A = 8'hF9; B = 8'hB5; #100;
A = 8'hF9; B = 8'hB6; #100;
A = 8'hF9; B = 8'hB7; #100;
A = 8'hF9; B = 8'hB8; #100;
A = 8'hF9; B = 8'hB9; #100;
A = 8'hF9; B = 8'hBA; #100;
A = 8'hF9; B = 8'hBB; #100;
A = 8'hF9; B = 8'hBC; #100;
A = 8'hF9; B = 8'hBD; #100;
A = 8'hF9; B = 8'hBE; #100;
A = 8'hF9; B = 8'hBF; #100;
A = 8'hF9; B = 8'hC0; #100;
A = 8'hF9; B = 8'hC1; #100;
A = 8'hF9; B = 8'hC2; #100;
A = 8'hF9; B = 8'hC3; #100;
A = 8'hF9; B = 8'hC4; #100;
A = 8'hF9; B = 8'hC5; #100;
A = 8'hF9; B = 8'hC6; #100;
A = 8'hF9; B = 8'hC7; #100;
A = 8'hF9; B = 8'hC8; #100;
A = 8'hF9; B = 8'hC9; #100;
A = 8'hF9; B = 8'hCA; #100;
A = 8'hF9; B = 8'hCB; #100;
A = 8'hF9; B = 8'hCC; #100;
A = 8'hF9; B = 8'hCD; #100;
A = 8'hF9; B = 8'hCE; #100;
A = 8'hF9; B = 8'hCF; #100;
A = 8'hF9; B = 8'hD0; #100;
A = 8'hF9; B = 8'hD1; #100;
A = 8'hF9; B = 8'hD2; #100;
A = 8'hF9; B = 8'hD3; #100;
A = 8'hF9; B = 8'hD4; #100;
A = 8'hF9; B = 8'hD5; #100;
A = 8'hF9; B = 8'hD6; #100;
A = 8'hF9; B = 8'hD7; #100;
A = 8'hF9; B = 8'hD8; #100;
A = 8'hF9; B = 8'hD9; #100;
A = 8'hF9; B = 8'hDA; #100;
A = 8'hF9; B = 8'hDB; #100;
A = 8'hF9; B = 8'hDC; #100;
A = 8'hF9; B = 8'hDD; #100;
A = 8'hF9; B = 8'hDE; #100;
A = 8'hF9; B = 8'hDF; #100;
A = 8'hF9; B = 8'hE0; #100;
A = 8'hF9; B = 8'hE1; #100;
A = 8'hF9; B = 8'hE2; #100;
A = 8'hF9; B = 8'hE3; #100;
A = 8'hF9; B = 8'hE4; #100;
A = 8'hF9; B = 8'hE5; #100;
A = 8'hF9; B = 8'hE6; #100;
A = 8'hF9; B = 8'hE7; #100;
A = 8'hF9; B = 8'hE8; #100;
A = 8'hF9; B = 8'hE9; #100;
A = 8'hF9; B = 8'hEA; #100;
A = 8'hF9; B = 8'hEB; #100;
A = 8'hF9; B = 8'hEC; #100;
A = 8'hF9; B = 8'hED; #100;
A = 8'hF9; B = 8'hEE; #100;
A = 8'hF9; B = 8'hEF; #100;
A = 8'hF9; B = 8'hF0; #100;
A = 8'hF9; B = 8'hF1; #100;
A = 8'hF9; B = 8'hF2; #100;
A = 8'hF9; B = 8'hF3; #100;
A = 8'hF9; B = 8'hF4; #100;
A = 8'hF9; B = 8'hF5; #100;
A = 8'hF9; B = 8'hF6; #100;
A = 8'hF9; B = 8'hF7; #100;
A = 8'hF9; B = 8'hF8; #100;
A = 8'hF9; B = 8'hF9; #100;
A = 8'hF9; B = 8'hFA; #100;
A = 8'hF9; B = 8'hFB; #100;
A = 8'hF9; B = 8'hFC; #100;
A = 8'hF9; B = 8'hFD; #100;
A = 8'hF9; B = 8'hFE; #100;
A = 8'hF9; B = 8'hFF; #100;
A = 8'hFA; B = 8'h0; #100;
A = 8'hFA; B = 8'h1; #100;
A = 8'hFA; B = 8'h2; #100;
A = 8'hFA; B = 8'h3; #100;
A = 8'hFA; B = 8'h4; #100;
A = 8'hFA; B = 8'h5; #100;
A = 8'hFA; B = 8'h6; #100;
A = 8'hFA; B = 8'h7; #100;
A = 8'hFA; B = 8'h8; #100;
A = 8'hFA; B = 8'h9; #100;
A = 8'hFA; B = 8'hA; #100;
A = 8'hFA; B = 8'hB; #100;
A = 8'hFA; B = 8'hC; #100;
A = 8'hFA; B = 8'hD; #100;
A = 8'hFA; B = 8'hE; #100;
A = 8'hFA; B = 8'hF; #100;
A = 8'hFA; B = 8'h10; #100;
A = 8'hFA; B = 8'h11; #100;
A = 8'hFA; B = 8'h12; #100;
A = 8'hFA; B = 8'h13; #100;
A = 8'hFA; B = 8'h14; #100;
A = 8'hFA; B = 8'h15; #100;
A = 8'hFA; B = 8'h16; #100;
A = 8'hFA; B = 8'h17; #100;
A = 8'hFA; B = 8'h18; #100;
A = 8'hFA; B = 8'h19; #100;
A = 8'hFA; B = 8'h1A; #100;
A = 8'hFA; B = 8'h1B; #100;
A = 8'hFA; B = 8'h1C; #100;
A = 8'hFA; B = 8'h1D; #100;
A = 8'hFA; B = 8'h1E; #100;
A = 8'hFA; B = 8'h1F; #100;
A = 8'hFA; B = 8'h20; #100;
A = 8'hFA; B = 8'h21; #100;
A = 8'hFA; B = 8'h22; #100;
A = 8'hFA; B = 8'h23; #100;
A = 8'hFA; B = 8'h24; #100;
A = 8'hFA; B = 8'h25; #100;
A = 8'hFA; B = 8'h26; #100;
A = 8'hFA; B = 8'h27; #100;
A = 8'hFA; B = 8'h28; #100;
A = 8'hFA; B = 8'h29; #100;
A = 8'hFA; B = 8'h2A; #100;
A = 8'hFA; B = 8'h2B; #100;
A = 8'hFA; B = 8'h2C; #100;
A = 8'hFA; B = 8'h2D; #100;
A = 8'hFA; B = 8'h2E; #100;
A = 8'hFA; B = 8'h2F; #100;
A = 8'hFA; B = 8'h30; #100;
A = 8'hFA; B = 8'h31; #100;
A = 8'hFA; B = 8'h32; #100;
A = 8'hFA; B = 8'h33; #100;
A = 8'hFA; B = 8'h34; #100;
A = 8'hFA; B = 8'h35; #100;
A = 8'hFA; B = 8'h36; #100;
A = 8'hFA; B = 8'h37; #100;
A = 8'hFA; B = 8'h38; #100;
A = 8'hFA; B = 8'h39; #100;
A = 8'hFA; B = 8'h3A; #100;
A = 8'hFA; B = 8'h3B; #100;
A = 8'hFA; B = 8'h3C; #100;
A = 8'hFA; B = 8'h3D; #100;
A = 8'hFA; B = 8'h3E; #100;
A = 8'hFA; B = 8'h3F; #100;
A = 8'hFA; B = 8'h40; #100;
A = 8'hFA; B = 8'h41; #100;
A = 8'hFA; B = 8'h42; #100;
A = 8'hFA; B = 8'h43; #100;
A = 8'hFA; B = 8'h44; #100;
A = 8'hFA; B = 8'h45; #100;
A = 8'hFA; B = 8'h46; #100;
A = 8'hFA; B = 8'h47; #100;
A = 8'hFA; B = 8'h48; #100;
A = 8'hFA; B = 8'h49; #100;
A = 8'hFA; B = 8'h4A; #100;
A = 8'hFA; B = 8'h4B; #100;
A = 8'hFA; B = 8'h4C; #100;
A = 8'hFA; B = 8'h4D; #100;
A = 8'hFA; B = 8'h4E; #100;
A = 8'hFA; B = 8'h4F; #100;
A = 8'hFA; B = 8'h50; #100;
A = 8'hFA; B = 8'h51; #100;
A = 8'hFA; B = 8'h52; #100;
A = 8'hFA; B = 8'h53; #100;
A = 8'hFA; B = 8'h54; #100;
A = 8'hFA; B = 8'h55; #100;
A = 8'hFA; B = 8'h56; #100;
A = 8'hFA; B = 8'h57; #100;
A = 8'hFA; B = 8'h58; #100;
A = 8'hFA; B = 8'h59; #100;
A = 8'hFA; B = 8'h5A; #100;
A = 8'hFA; B = 8'h5B; #100;
A = 8'hFA; B = 8'h5C; #100;
A = 8'hFA; B = 8'h5D; #100;
A = 8'hFA; B = 8'h5E; #100;
A = 8'hFA; B = 8'h5F; #100;
A = 8'hFA; B = 8'h60; #100;
A = 8'hFA; B = 8'h61; #100;
A = 8'hFA; B = 8'h62; #100;
A = 8'hFA; B = 8'h63; #100;
A = 8'hFA; B = 8'h64; #100;
A = 8'hFA; B = 8'h65; #100;
A = 8'hFA; B = 8'h66; #100;
A = 8'hFA; B = 8'h67; #100;
A = 8'hFA; B = 8'h68; #100;
A = 8'hFA; B = 8'h69; #100;
A = 8'hFA; B = 8'h6A; #100;
A = 8'hFA; B = 8'h6B; #100;
A = 8'hFA; B = 8'h6C; #100;
A = 8'hFA; B = 8'h6D; #100;
A = 8'hFA; B = 8'h6E; #100;
A = 8'hFA; B = 8'h6F; #100;
A = 8'hFA; B = 8'h70; #100;
A = 8'hFA; B = 8'h71; #100;
A = 8'hFA; B = 8'h72; #100;
A = 8'hFA; B = 8'h73; #100;
A = 8'hFA; B = 8'h74; #100;
A = 8'hFA; B = 8'h75; #100;
A = 8'hFA; B = 8'h76; #100;
A = 8'hFA; B = 8'h77; #100;
A = 8'hFA; B = 8'h78; #100;
A = 8'hFA; B = 8'h79; #100;
A = 8'hFA; B = 8'h7A; #100;
A = 8'hFA; B = 8'h7B; #100;
A = 8'hFA; B = 8'h7C; #100;
A = 8'hFA; B = 8'h7D; #100;
A = 8'hFA; B = 8'h7E; #100;
A = 8'hFA; B = 8'h7F; #100;
A = 8'hFA; B = 8'h80; #100;
A = 8'hFA; B = 8'h81; #100;
A = 8'hFA; B = 8'h82; #100;
A = 8'hFA; B = 8'h83; #100;
A = 8'hFA; B = 8'h84; #100;
A = 8'hFA; B = 8'h85; #100;
A = 8'hFA; B = 8'h86; #100;
A = 8'hFA; B = 8'h87; #100;
A = 8'hFA; B = 8'h88; #100;
A = 8'hFA; B = 8'h89; #100;
A = 8'hFA; B = 8'h8A; #100;
A = 8'hFA; B = 8'h8B; #100;
A = 8'hFA; B = 8'h8C; #100;
A = 8'hFA; B = 8'h8D; #100;
A = 8'hFA; B = 8'h8E; #100;
A = 8'hFA; B = 8'h8F; #100;
A = 8'hFA; B = 8'h90; #100;
A = 8'hFA; B = 8'h91; #100;
A = 8'hFA; B = 8'h92; #100;
A = 8'hFA; B = 8'h93; #100;
A = 8'hFA; B = 8'h94; #100;
A = 8'hFA; B = 8'h95; #100;
A = 8'hFA; B = 8'h96; #100;
A = 8'hFA; B = 8'h97; #100;
A = 8'hFA; B = 8'h98; #100;
A = 8'hFA; B = 8'h99; #100;
A = 8'hFA; B = 8'h9A; #100;
A = 8'hFA; B = 8'h9B; #100;
A = 8'hFA; B = 8'h9C; #100;
A = 8'hFA; B = 8'h9D; #100;
A = 8'hFA; B = 8'h9E; #100;
A = 8'hFA; B = 8'h9F; #100;
A = 8'hFA; B = 8'hA0; #100;
A = 8'hFA; B = 8'hA1; #100;
A = 8'hFA; B = 8'hA2; #100;
A = 8'hFA; B = 8'hA3; #100;
A = 8'hFA; B = 8'hA4; #100;
A = 8'hFA; B = 8'hA5; #100;
A = 8'hFA; B = 8'hA6; #100;
A = 8'hFA; B = 8'hA7; #100;
A = 8'hFA; B = 8'hA8; #100;
A = 8'hFA; B = 8'hA9; #100;
A = 8'hFA; B = 8'hAA; #100;
A = 8'hFA; B = 8'hAB; #100;
A = 8'hFA; B = 8'hAC; #100;
A = 8'hFA; B = 8'hAD; #100;
A = 8'hFA; B = 8'hAE; #100;
A = 8'hFA; B = 8'hAF; #100;
A = 8'hFA; B = 8'hB0; #100;
A = 8'hFA; B = 8'hB1; #100;
A = 8'hFA; B = 8'hB2; #100;
A = 8'hFA; B = 8'hB3; #100;
A = 8'hFA; B = 8'hB4; #100;
A = 8'hFA; B = 8'hB5; #100;
A = 8'hFA; B = 8'hB6; #100;
A = 8'hFA; B = 8'hB7; #100;
A = 8'hFA; B = 8'hB8; #100;
A = 8'hFA; B = 8'hB9; #100;
A = 8'hFA; B = 8'hBA; #100;
A = 8'hFA; B = 8'hBB; #100;
A = 8'hFA; B = 8'hBC; #100;
A = 8'hFA; B = 8'hBD; #100;
A = 8'hFA; B = 8'hBE; #100;
A = 8'hFA; B = 8'hBF; #100;
A = 8'hFA; B = 8'hC0; #100;
A = 8'hFA; B = 8'hC1; #100;
A = 8'hFA; B = 8'hC2; #100;
A = 8'hFA; B = 8'hC3; #100;
A = 8'hFA; B = 8'hC4; #100;
A = 8'hFA; B = 8'hC5; #100;
A = 8'hFA; B = 8'hC6; #100;
A = 8'hFA; B = 8'hC7; #100;
A = 8'hFA; B = 8'hC8; #100;
A = 8'hFA; B = 8'hC9; #100;
A = 8'hFA; B = 8'hCA; #100;
A = 8'hFA; B = 8'hCB; #100;
A = 8'hFA; B = 8'hCC; #100;
A = 8'hFA; B = 8'hCD; #100;
A = 8'hFA; B = 8'hCE; #100;
A = 8'hFA; B = 8'hCF; #100;
A = 8'hFA; B = 8'hD0; #100;
A = 8'hFA; B = 8'hD1; #100;
A = 8'hFA; B = 8'hD2; #100;
A = 8'hFA; B = 8'hD3; #100;
A = 8'hFA; B = 8'hD4; #100;
A = 8'hFA; B = 8'hD5; #100;
A = 8'hFA; B = 8'hD6; #100;
A = 8'hFA; B = 8'hD7; #100;
A = 8'hFA; B = 8'hD8; #100;
A = 8'hFA; B = 8'hD9; #100;
A = 8'hFA; B = 8'hDA; #100;
A = 8'hFA; B = 8'hDB; #100;
A = 8'hFA; B = 8'hDC; #100;
A = 8'hFA; B = 8'hDD; #100;
A = 8'hFA; B = 8'hDE; #100;
A = 8'hFA; B = 8'hDF; #100;
A = 8'hFA; B = 8'hE0; #100;
A = 8'hFA; B = 8'hE1; #100;
A = 8'hFA; B = 8'hE2; #100;
A = 8'hFA; B = 8'hE3; #100;
A = 8'hFA; B = 8'hE4; #100;
A = 8'hFA; B = 8'hE5; #100;
A = 8'hFA; B = 8'hE6; #100;
A = 8'hFA; B = 8'hE7; #100;
A = 8'hFA; B = 8'hE8; #100;
A = 8'hFA; B = 8'hE9; #100;
A = 8'hFA; B = 8'hEA; #100;
A = 8'hFA; B = 8'hEB; #100;
A = 8'hFA; B = 8'hEC; #100;
A = 8'hFA; B = 8'hED; #100;
A = 8'hFA; B = 8'hEE; #100;
A = 8'hFA; B = 8'hEF; #100;
A = 8'hFA; B = 8'hF0; #100;
A = 8'hFA; B = 8'hF1; #100;
A = 8'hFA; B = 8'hF2; #100;
A = 8'hFA; B = 8'hF3; #100;
A = 8'hFA; B = 8'hF4; #100;
A = 8'hFA; B = 8'hF5; #100;
A = 8'hFA; B = 8'hF6; #100;
A = 8'hFA; B = 8'hF7; #100;
A = 8'hFA; B = 8'hF8; #100;
A = 8'hFA; B = 8'hF9; #100;
A = 8'hFA; B = 8'hFA; #100;
A = 8'hFA; B = 8'hFB; #100;
A = 8'hFA; B = 8'hFC; #100;
A = 8'hFA; B = 8'hFD; #100;
A = 8'hFA; B = 8'hFE; #100;
A = 8'hFA; B = 8'hFF; #100;
A = 8'hFB; B = 8'h0; #100;
A = 8'hFB; B = 8'h1; #100;
A = 8'hFB; B = 8'h2; #100;
A = 8'hFB; B = 8'h3; #100;
A = 8'hFB; B = 8'h4; #100;
A = 8'hFB; B = 8'h5; #100;
A = 8'hFB; B = 8'h6; #100;
A = 8'hFB; B = 8'h7; #100;
A = 8'hFB; B = 8'h8; #100;
A = 8'hFB; B = 8'h9; #100;
A = 8'hFB; B = 8'hA; #100;
A = 8'hFB; B = 8'hB; #100;
A = 8'hFB; B = 8'hC; #100;
A = 8'hFB; B = 8'hD; #100;
A = 8'hFB; B = 8'hE; #100;
A = 8'hFB; B = 8'hF; #100;
A = 8'hFB; B = 8'h10; #100;
A = 8'hFB; B = 8'h11; #100;
A = 8'hFB; B = 8'h12; #100;
A = 8'hFB; B = 8'h13; #100;
A = 8'hFB; B = 8'h14; #100;
A = 8'hFB; B = 8'h15; #100;
A = 8'hFB; B = 8'h16; #100;
A = 8'hFB; B = 8'h17; #100;
A = 8'hFB; B = 8'h18; #100;
A = 8'hFB; B = 8'h19; #100;
A = 8'hFB; B = 8'h1A; #100;
A = 8'hFB; B = 8'h1B; #100;
A = 8'hFB; B = 8'h1C; #100;
A = 8'hFB; B = 8'h1D; #100;
A = 8'hFB; B = 8'h1E; #100;
A = 8'hFB; B = 8'h1F; #100;
A = 8'hFB; B = 8'h20; #100;
A = 8'hFB; B = 8'h21; #100;
A = 8'hFB; B = 8'h22; #100;
A = 8'hFB; B = 8'h23; #100;
A = 8'hFB; B = 8'h24; #100;
A = 8'hFB; B = 8'h25; #100;
A = 8'hFB; B = 8'h26; #100;
A = 8'hFB; B = 8'h27; #100;
A = 8'hFB; B = 8'h28; #100;
A = 8'hFB; B = 8'h29; #100;
A = 8'hFB; B = 8'h2A; #100;
A = 8'hFB; B = 8'h2B; #100;
A = 8'hFB; B = 8'h2C; #100;
A = 8'hFB; B = 8'h2D; #100;
A = 8'hFB; B = 8'h2E; #100;
A = 8'hFB; B = 8'h2F; #100;
A = 8'hFB; B = 8'h30; #100;
A = 8'hFB; B = 8'h31; #100;
A = 8'hFB; B = 8'h32; #100;
A = 8'hFB; B = 8'h33; #100;
A = 8'hFB; B = 8'h34; #100;
A = 8'hFB; B = 8'h35; #100;
A = 8'hFB; B = 8'h36; #100;
A = 8'hFB; B = 8'h37; #100;
A = 8'hFB; B = 8'h38; #100;
A = 8'hFB; B = 8'h39; #100;
A = 8'hFB; B = 8'h3A; #100;
A = 8'hFB; B = 8'h3B; #100;
A = 8'hFB; B = 8'h3C; #100;
A = 8'hFB; B = 8'h3D; #100;
A = 8'hFB; B = 8'h3E; #100;
A = 8'hFB; B = 8'h3F; #100;
A = 8'hFB; B = 8'h40; #100;
A = 8'hFB; B = 8'h41; #100;
A = 8'hFB; B = 8'h42; #100;
A = 8'hFB; B = 8'h43; #100;
A = 8'hFB; B = 8'h44; #100;
A = 8'hFB; B = 8'h45; #100;
A = 8'hFB; B = 8'h46; #100;
A = 8'hFB; B = 8'h47; #100;
A = 8'hFB; B = 8'h48; #100;
A = 8'hFB; B = 8'h49; #100;
A = 8'hFB; B = 8'h4A; #100;
A = 8'hFB; B = 8'h4B; #100;
A = 8'hFB; B = 8'h4C; #100;
A = 8'hFB; B = 8'h4D; #100;
A = 8'hFB; B = 8'h4E; #100;
A = 8'hFB; B = 8'h4F; #100;
A = 8'hFB; B = 8'h50; #100;
A = 8'hFB; B = 8'h51; #100;
A = 8'hFB; B = 8'h52; #100;
A = 8'hFB; B = 8'h53; #100;
A = 8'hFB; B = 8'h54; #100;
A = 8'hFB; B = 8'h55; #100;
A = 8'hFB; B = 8'h56; #100;
A = 8'hFB; B = 8'h57; #100;
A = 8'hFB; B = 8'h58; #100;
A = 8'hFB; B = 8'h59; #100;
A = 8'hFB; B = 8'h5A; #100;
A = 8'hFB; B = 8'h5B; #100;
A = 8'hFB; B = 8'h5C; #100;
A = 8'hFB; B = 8'h5D; #100;
A = 8'hFB; B = 8'h5E; #100;
A = 8'hFB; B = 8'h5F; #100;
A = 8'hFB; B = 8'h60; #100;
A = 8'hFB; B = 8'h61; #100;
A = 8'hFB; B = 8'h62; #100;
A = 8'hFB; B = 8'h63; #100;
A = 8'hFB; B = 8'h64; #100;
A = 8'hFB; B = 8'h65; #100;
A = 8'hFB; B = 8'h66; #100;
A = 8'hFB; B = 8'h67; #100;
A = 8'hFB; B = 8'h68; #100;
A = 8'hFB; B = 8'h69; #100;
A = 8'hFB; B = 8'h6A; #100;
A = 8'hFB; B = 8'h6B; #100;
A = 8'hFB; B = 8'h6C; #100;
A = 8'hFB; B = 8'h6D; #100;
A = 8'hFB; B = 8'h6E; #100;
A = 8'hFB; B = 8'h6F; #100;
A = 8'hFB; B = 8'h70; #100;
A = 8'hFB; B = 8'h71; #100;
A = 8'hFB; B = 8'h72; #100;
A = 8'hFB; B = 8'h73; #100;
A = 8'hFB; B = 8'h74; #100;
A = 8'hFB; B = 8'h75; #100;
A = 8'hFB; B = 8'h76; #100;
A = 8'hFB; B = 8'h77; #100;
A = 8'hFB; B = 8'h78; #100;
A = 8'hFB; B = 8'h79; #100;
A = 8'hFB; B = 8'h7A; #100;
A = 8'hFB; B = 8'h7B; #100;
A = 8'hFB; B = 8'h7C; #100;
A = 8'hFB; B = 8'h7D; #100;
A = 8'hFB; B = 8'h7E; #100;
A = 8'hFB; B = 8'h7F; #100;
A = 8'hFB; B = 8'h80; #100;
A = 8'hFB; B = 8'h81; #100;
A = 8'hFB; B = 8'h82; #100;
A = 8'hFB; B = 8'h83; #100;
A = 8'hFB; B = 8'h84; #100;
A = 8'hFB; B = 8'h85; #100;
A = 8'hFB; B = 8'h86; #100;
A = 8'hFB; B = 8'h87; #100;
A = 8'hFB; B = 8'h88; #100;
A = 8'hFB; B = 8'h89; #100;
A = 8'hFB; B = 8'h8A; #100;
A = 8'hFB; B = 8'h8B; #100;
A = 8'hFB; B = 8'h8C; #100;
A = 8'hFB; B = 8'h8D; #100;
A = 8'hFB; B = 8'h8E; #100;
A = 8'hFB; B = 8'h8F; #100;
A = 8'hFB; B = 8'h90; #100;
A = 8'hFB; B = 8'h91; #100;
A = 8'hFB; B = 8'h92; #100;
A = 8'hFB; B = 8'h93; #100;
A = 8'hFB; B = 8'h94; #100;
A = 8'hFB; B = 8'h95; #100;
A = 8'hFB; B = 8'h96; #100;
A = 8'hFB; B = 8'h97; #100;
A = 8'hFB; B = 8'h98; #100;
A = 8'hFB; B = 8'h99; #100;
A = 8'hFB; B = 8'h9A; #100;
A = 8'hFB; B = 8'h9B; #100;
A = 8'hFB; B = 8'h9C; #100;
A = 8'hFB; B = 8'h9D; #100;
A = 8'hFB; B = 8'h9E; #100;
A = 8'hFB; B = 8'h9F; #100;
A = 8'hFB; B = 8'hA0; #100;
A = 8'hFB; B = 8'hA1; #100;
A = 8'hFB; B = 8'hA2; #100;
A = 8'hFB; B = 8'hA3; #100;
A = 8'hFB; B = 8'hA4; #100;
A = 8'hFB; B = 8'hA5; #100;
A = 8'hFB; B = 8'hA6; #100;
A = 8'hFB; B = 8'hA7; #100;
A = 8'hFB; B = 8'hA8; #100;
A = 8'hFB; B = 8'hA9; #100;
A = 8'hFB; B = 8'hAA; #100;
A = 8'hFB; B = 8'hAB; #100;
A = 8'hFB; B = 8'hAC; #100;
A = 8'hFB; B = 8'hAD; #100;
A = 8'hFB; B = 8'hAE; #100;
A = 8'hFB; B = 8'hAF; #100;
A = 8'hFB; B = 8'hB0; #100;
A = 8'hFB; B = 8'hB1; #100;
A = 8'hFB; B = 8'hB2; #100;
A = 8'hFB; B = 8'hB3; #100;
A = 8'hFB; B = 8'hB4; #100;
A = 8'hFB; B = 8'hB5; #100;
A = 8'hFB; B = 8'hB6; #100;
A = 8'hFB; B = 8'hB7; #100;
A = 8'hFB; B = 8'hB8; #100;
A = 8'hFB; B = 8'hB9; #100;
A = 8'hFB; B = 8'hBA; #100;
A = 8'hFB; B = 8'hBB; #100;
A = 8'hFB; B = 8'hBC; #100;
A = 8'hFB; B = 8'hBD; #100;
A = 8'hFB; B = 8'hBE; #100;
A = 8'hFB; B = 8'hBF; #100;
A = 8'hFB; B = 8'hC0; #100;
A = 8'hFB; B = 8'hC1; #100;
A = 8'hFB; B = 8'hC2; #100;
A = 8'hFB; B = 8'hC3; #100;
A = 8'hFB; B = 8'hC4; #100;
A = 8'hFB; B = 8'hC5; #100;
A = 8'hFB; B = 8'hC6; #100;
A = 8'hFB; B = 8'hC7; #100;
A = 8'hFB; B = 8'hC8; #100;
A = 8'hFB; B = 8'hC9; #100;
A = 8'hFB; B = 8'hCA; #100;
A = 8'hFB; B = 8'hCB; #100;
A = 8'hFB; B = 8'hCC; #100;
A = 8'hFB; B = 8'hCD; #100;
A = 8'hFB; B = 8'hCE; #100;
A = 8'hFB; B = 8'hCF; #100;
A = 8'hFB; B = 8'hD0; #100;
A = 8'hFB; B = 8'hD1; #100;
A = 8'hFB; B = 8'hD2; #100;
A = 8'hFB; B = 8'hD3; #100;
A = 8'hFB; B = 8'hD4; #100;
A = 8'hFB; B = 8'hD5; #100;
A = 8'hFB; B = 8'hD6; #100;
A = 8'hFB; B = 8'hD7; #100;
A = 8'hFB; B = 8'hD8; #100;
A = 8'hFB; B = 8'hD9; #100;
A = 8'hFB; B = 8'hDA; #100;
A = 8'hFB; B = 8'hDB; #100;
A = 8'hFB; B = 8'hDC; #100;
A = 8'hFB; B = 8'hDD; #100;
A = 8'hFB; B = 8'hDE; #100;
A = 8'hFB; B = 8'hDF; #100;
A = 8'hFB; B = 8'hE0; #100;
A = 8'hFB; B = 8'hE1; #100;
A = 8'hFB; B = 8'hE2; #100;
A = 8'hFB; B = 8'hE3; #100;
A = 8'hFB; B = 8'hE4; #100;
A = 8'hFB; B = 8'hE5; #100;
A = 8'hFB; B = 8'hE6; #100;
A = 8'hFB; B = 8'hE7; #100;
A = 8'hFB; B = 8'hE8; #100;
A = 8'hFB; B = 8'hE9; #100;
A = 8'hFB; B = 8'hEA; #100;
A = 8'hFB; B = 8'hEB; #100;
A = 8'hFB; B = 8'hEC; #100;
A = 8'hFB; B = 8'hED; #100;
A = 8'hFB; B = 8'hEE; #100;
A = 8'hFB; B = 8'hEF; #100;
A = 8'hFB; B = 8'hF0; #100;
A = 8'hFB; B = 8'hF1; #100;
A = 8'hFB; B = 8'hF2; #100;
A = 8'hFB; B = 8'hF3; #100;
A = 8'hFB; B = 8'hF4; #100;
A = 8'hFB; B = 8'hF5; #100;
A = 8'hFB; B = 8'hF6; #100;
A = 8'hFB; B = 8'hF7; #100;
A = 8'hFB; B = 8'hF8; #100;
A = 8'hFB; B = 8'hF9; #100;
A = 8'hFB; B = 8'hFA; #100;
A = 8'hFB; B = 8'hFB; #100;
A = 8'hFB; B = 8'hFC; #100;
A = 8'hFB; B = 8'hFD; #100;
A = 8'hFB; B = 8'hFE; #100;
A = 8'hFB; B = 8'hFF; #100;
A = 8'hFC; B = 8'h0; #100;
A = 8'hFC; B = 8'h1; #100;
A = 8'hFC; B = 8'h2; #100;
A = 8'hFC; B = 8'h3; #100;
A = 8'hFC; B = 8'h4; #100;
A = 8'hFC; B = 8'h5; #100;
A = 8'hFC; B = 8'h6; #100;
A = 8'hFC; B = 8'h7; #100;
A = 8'hFC; B = 8'h8; #100;
A = 8'hFC; B = 8'h9; #100;
A = 8'hFC; B = 8'hA; #100;
A = 8'hFC; B = 8'hB; #100;
A = 8'hFC; B = 8'hC; #100;
A = 8'hFC; B = 8'hD; #100;
A = 8'hFC; B = 8'hE; #100;
A = 8'hFC; B = 8'hF; #100;
A = 8'hFC; B = 8'h10; #100;
A = 8'hFC; B = 8'h11; #100;
A = 8'hFC; B = 8'h12; #100;
A = 8'hFC; B = 8'h13; #100;
A = 8'hFC; B = 8'h14; #100;
A = 8'hFC; B = 8'h15; #100;
A = 8'hFC; B = 8'h16; #100;
A = 8'hFC; B = 8'h17; #100;
A = 8'hFC; B = 8'h18; #100;
A = 8'hFC; B = 8'h19; #100;
A = 8'hFC; B = 8'h1A; #100;
A = 8'hFC; B = 8'h1B; #100;
A = 8'hFC; B = 8'h1C; #100;
A = 8'hFC; B = 8'h1D; #100;
A = 8'hFC; B = 8'h1E; #100;
A = 8'hFC; B = 8'h1F; #100;
A = 8'hFC; B = 8'h20; #100;
A = 8'hFC; B = 8'h21; #100;
A = 8'hFC; B = 8'h22; #100;
A = 8'hFC; B = 8'h23; #100;
A = 8'hFC; B = 8'h24; #100;
A = 8'hFC; B = 8'h25; #100;
A = 8'hFC; B = 8'h26; #100;
A = 8'hFC; B = 8'h27; #100;
A = 8'hFC; B = 8'h28; #100;
A = 8'hFC; B = 8'h29; #100;
A = 8'hFC; B = 8'h2A; #100;
A = 8'hFC; B = 8'h2B; #100;
A = 8'hFC; B = 8'h2C; #100;
A = 8'hFC; B = 8'h2D; #100;
A = 8'hFC; B = 8'h2E; #100;
A = 8'hFC; B = 8'h2F; #100;
A = 8'hFC; B = 8'h30; #100;
A = 8'hFC; B = 8'h31; #100;
A = 8'hFC; B = 8'h32; #100;
A = 8'hFC; B = 8'h33; #100;
A = 8'hFC; B = 8'h34; #100;
A = 8'hFC; B = 8'h35; #100;
A = 8'hFC; B = 8'h36; #100;
A = 8'hFC; B = 8'h37; #100;
A = 8'hFC; B = 8'h38; #100;
A = 8'hFC; B = 8'h39; #100;
A = 8'hFC; B = 8'h3A; #100;
A = 8'hFC; B = 8'h3B; #100;
A = 8'hFC; B = 8'h3C; #100;
A = 8'hFC; B = 8'h3D; #100;
A = 8'hFC; B = 8'h3E; #100;
A = 8'hFC; B = 8'h3F; #100;
A = 8'hFC; B = 8'h40; #100;
A = 8'hFC; B = 8'h41; #100;
A = 8'hFC; B = 8'h42; #100;
A = 8'hFC; B = 8'h43; #100;
A = 8'hFC; B = 8'h44; #100;
A = 8'hFC; B = 8'h45; #100;
A = 8'hFC; B = 8'h46; #100;
A = 8'hFC; B = 8'h47; #100;
A = 8'hFC; B = 8'h48; #100;
A = 8'hFC; B = 8'h49; #100;
A = 8'hFC; B = 8'h4A; #100;
A = 8'hFC; B = 8'h4B; #100;
A = 8'hFC; B = 8'h4C; #100;
A = 8'hFC; B = 8'h4D; #100;
A = 8'hFC; B = 8'h4E; #100;
A = 8'hFC; B = 8'h4F; #100;
A = 8'hFC; B = 8'h50; #100;
A = 8'hFC; B = 8'h51; #100;
A = 8'hFC; B = 8'h52; #100;
A = 8'hFC; B = 8'h53; #100;
A = 8'hFC; B = 8'h54; #100;
A = 8'hFC; B = 8'h55; #100;
A = 8'hFC; B = 8'h56; #100;
A = 8'hFC; B = 8'h57; #100;
A = 8'hFC; B = 8'h58; #100;
A = 8'hFC; B = 8'h59; #100;
A = 8'hFC; B = 8'h5A; #100;
A = 8'hFC; B = 8'h5B; #100;
A = 8'hFC; B = 8'h5C; #100;
A = 8'hFC; B = 8'h5D; #100;
A = 8'hFC; B = 8'h5E; #100;
A = 8'hFC; B = 8'h5F; #100;
A = 8'hFC; B = 8'h60; #100;
A = 8'hFC; B = 8'h61; #100;
A = 8'hFC; B = 8'h62; #100;
A = 8'hFC; B = 8'h63; #100;
A = 8'hFC; B = 8'h64; #100;
A = 8'hFC; B = 8'h65; #100;
A = 8'hFC; B = 8'h66; #100;
A = 8'hFC; B = 8'h67; #100;
A = 8'hFC; B = 8'h68; #100;
A = 8'hFC; B = 8'h69; #100;
A = 8'hFC; B = 8'h6A; #100;
A = 8'hFC; B = 8'h6B; #100;
A = 8'hFC; B = 8'h6C; #100;
A = 8'hFC; B = 8'h6D; #100;
A = 8'hFC; B = 8'h6E; #100;
A = 8'hFC; B = 8'h6F; #100;
A = 8'hFC; B = 8'h70; #100;
A = 8'hFC; B = 8'h71; #100;
A = 8'hFC; B = 8'h72; #100;
A = 8'hFC; B = 8'h73; #100;
A = 8'hFC; B = 8'h74; #100;
A = 8'hFC; B = 8'h75; #100;
A = 8'hFC; B = 8'h76; #100;
A = 8'hFC; B = 8'h77; #100;
A = 8'hFC; B = 8'h78; #100;
A = 8'hFC; B = 8'h79; #100;
A = 8'hFC; B = 8'h7A; #100;
A = 8'hFC; B = 8'h7B; #100;
A = 8'hFC; B = 8'h7C; #100;
A = 8'hFC; B = 8'h7D; #100;
A = 8'hFC; B = 8'h7E; #100;
A = 8'hFC; B = 8'h7F; #100;
A = 8'hFC; B = 8'h80; #100;
A = 8'hFC; B = 8'h81; #100;
A = 8'hFC; B = 8'h82; #100;
A = 8'hFC; B = 8'h83; #100;
A = 8'hFC; B = 8'h84; #100;
A = 8'hFC; B = 8'h85; #100;
A = 8'hFC; B = 8'h86; #100;
A = 8'hFC; B = 8'h87; #100;
A = 8'hFC; B = 8'h88; #100;
A = 8'hFC; B = 8'h89; #100;
A = 8'hFC; B = 8'h8A; #100;
A = 8'hFC; B = 8'h8B; #100;
A = 8'hFC; B = 8'h8C; #100;
A = 8'hFC; B = 8'h8D; #100;
A = 8'hFC; B = 8'h8E; #100;
A = 8'hFC; B = 8'h8F; #100;
A = 8'hFC; B = 8'h90; #100;
A = 8'hFC; B = 8'h91; #100;
A = 8'hFC; B = 8'h92; #100;
A = 8'hFC; B = 8'h93; #100;
A = 8'hFC; B = 8'h94; #100;
A = 8'hFC; B = 8'h95; #100;
A = 8'hFC; B = 8'h96; #100;
A = 8'hFC; B = 8'h97; #100;
A = 8'hFC; B = 8'h98; #100;
A = 8'hFC; B = 8'h99; #100;
A = 8'hFC; B = 8'h9A; #100;
A = 8'hFC; B = 8'h9B; #100;
A = 8'hFC; B = 8'h9C; #100;
A = 8'hFC; B = 8'h9D; #100;
A = 8'hFC; B = 8'h9E; #100;
A = 8'hFC; B = 8'h9F; #100;
A = 8'hFC; B = 8'hA0; #100;
A = 8'hFC; B = 8'hA1; #100;
A = 8'hFC; B = 8'hA2; #100;
A = 8'hFC; B = 8'hA3; #100;
A = 8'hFC; B = 8'hA4; #100;
A = 8'hFC; B = 8'hA5; #100;
A = 8'hFC; B = 8'hA6; #100;
A = 8'hFC; B = 8'hA7; #100;
A = 8'hFC; B = 8'hA8; #100;
A = 8'hFC; B = 8'hA9; #100;
A = 8'hFC; B = 8'hAA; #100;
A = 8'hFC; B = 8'hAB; #100;
A = 8'hFC; B = 8'hAC; #100;
A = 8'hFC; B = 8'hAD; #100;
A = 8'hFC; B = 8'hAE; #100;
A = 8'hFC; B = 8'hAF; #100;
A = 8'hFC; B = 8'hB0; #100;
A = 8'hFC; B = 8'hB1; #100;
A = 8'hFC; B = 8'hB2; #100;
A = 8'hFC; B = 8'hB3; #100;
A = 8'hFC; B = 8'hB4; #100;
A = 8'hFC; B = 8'hB5; #100;
A = 8'hFC; B = 8'hB6; #100;
A = 8'hFC; B = 8'hB7; #100;
A = 8'hFC; B = 8'hB8; #100;
A = 8'hFC; B = 8'hB9; #100;
A = 8'hFC; B = 8'hBA; #100;
A = 8'hFC; B = 8'hBB; #100;
A = 8'hFC; B = 8'hBC; #100;
A = 8'hFC; B = 8'hBD; #100;
A = 8'hFC; B = 8'hBE; #100;
A = 8'hFC; B = 8'hBF; #100;
A = 8'hFC; B = 8'hC0; #100;
A = 8'hFC; B = 8'hC1; #100;
A = 8'hFC; B = 8'hC2; #100;
A = 8'hFC; B = 8'hC3; #100;
A = 8'hFC; B = 8'hC4; #100;
A = 8'hFC; B = 8'hC5; #100;
A = 8'hFC; B = 8'hC6; #100;
A = 8'hFC; B = 8'hC7; #100;
A = 8'hFC; B = 8'hC8; #100;
A = 8'hFC; B = 8'hC9; #100;
A = 8'hFC; B = 8'hCA; #100;
A = 8'hFC; B = 8'hCB; #100;
A = 8'hFC; B = 8'hCC; #100;
A = 8'hFC; B = 8'hCD; #100;
A = 8'hFC; B = 8'hCE; #100;
A = 8'hFC; B = 8'hCF; #100;
A = 8'hFC; B = 8'hD0; #100;
A = 8'hFC; B = 8'hD1; #100;
A = 8'hFC; B = 8'hD2; #100;
A = 8'hFC; B = 8'hD3; #100;
A = 8'hFC; B = 8'hD4; #100;
A = 8'hFC; B = 8'hD5; #100;
A = 8'hFC; B = 8'hD6; #100;
A = 8'hFC; B = 8'hD7; #100;
A = 8'hFC; B = 8'hD8; #100;
A = 8'hFC; B = 8'hD9; #100;
A = 8'hFC; B = 8'hDA; #100;
A = 8'hFC; B = 8'hDB; #100;
A = 8'hFC; B = 8'hDC; #100;
A = 8'hFC; B = 8'hDD; #100;
A = 8'hFC; B = 8'hDE; #100;
A = 8'hFC; B = 8'hDF; #100;
A = 8'hFC; B = 8'hE0; #100;
A = 8'hFC; B = 8'hE1; #100;
A = 8'hFC; B = 8'hE2; #100;
A = 8'hFC; B = 8'hE3; #100;
A = 8'hFC; B = 8'hE4; #100;
A = 8'hFC; B = 8'hE5; #100;
A = 8'hFC; B = 8'hE6; #100;
A = 8'hFC; B = 8'hE7; #100;
A = 8'hFC; B = 8'hE8; #100;
A = 8'hFC; B = 8'hE9; #100;
A = 8'hFC; B = 8'hEA; #100;
A = 8'hFC; B = 8'hEB; #100;
A = 8'hFC; B = 8'hEC; #100;
A = 8'hFC; B = 8'hED; #100;
A = 8'hFC; B = 8'hEE; #100;
A = 8'hFC; B = 8'hEF; #100;
A = 8'hFC; B = 8'hF0; #100;
A = 8'hFC; B = 8'hF1; #100;
A = 8'hFC; B = 8'hF2; #100;
A = 8'hFC; B = 8'hF3; #100;
A = 8'hFC; B = 8'hF4; #100;
A = 8'hFC; B = 8'hF5; #100;
A = 8'hFC; B = 8'hF6; #100;
A = 8'hFC; B = 8'hF7; #100;
A = 8'hFC; B = 8'hF8; #100;
A = 8'hFC; B = 8'hF9; #100;
A = 8'hFC; B = 8'hFA; #100;
A = 8'hFC; B = 8'hFB; #100;
A = 8'hFC; B = 8'hFC; #100;
A = 8'hFC; B = 8'hFD; #100;
A = 8'hFC; B = 8'hFE; #100;
A = 8'hFC; B = 8'hFF; #100;
A = 8'hFD; B = 8'h0; #100;
A = 8'hFD; B = 8'h1; #100;
A = 8'hFD; B = 8'h2; #100;
A = 8'hFD; B = 8'h3; #100;
A = 8'hFD; B = 8'h4; #100;
A = 8'hFD; B = 8'h5; #100;
A = 8'hFD; B = 8'h6; #100;
A = 8'hFD; B = 8'h7; #100;
A = 8'hFD; B = 8'h8; #100;
A = 8'hFD; B = 8'h9; #100;
A = 8'hFD; B = 8'hA; #100;
A = 8'hFD; B = 8'hB; #100;
A = 8'hFD; B = 8'hC; #100;
A = 8'hFD; B = 8'hD; #100;
A = 8'hFD; B = 8'hE; #100;
A = 8'hFD; B = 8'hF; #100;
A = 8'hFD; B = 8'h10; #100;
A = 8'hFD; B = 8'h11; #100;
A = 8'hFD; B = 8'h12; #100;
A = 8'hFD; B = 8'h13; #100;
A = 8'hFD; B = 8'h14; #100;
A = 8'hFD; B = 8'h15; #100;
A = 8'hFD; B = 8'h16; #100;
A = 8'hFD; B = 8'h17; #100;
A = 8'hFD; B = 8'h18; #100;
A = 8'hFD; B = 8'h19; #100;
A = 8'hFD; B = 8'h1A; #100;
A = 8'hFD; B = 8'h1B; #100;
A = 8'hFD; B = 8'h1C; #100;
A = 8'hFD; B = 8'h1D; #100;
A = 8'hFD; B = 8'h1E; #100;
A = 8'hFD; B = 8'h1F; #100;
A = 8'hFD; B = 8'h20; #100;
A = 8'hFD; B = 8'h21; #100;
A = 8'hFD; B = 8'h22; #100;
A = 8'hFD; B = 8'h23; #100;
A = 8'hFD; B = 8'h24; #100;
A = 8'hFD; B = 8'h25; #100;
A = 8'hFD; B = 8'h26; #100;
A = 8'hFD; B = 8'h27; #100;
A = 8'hFD; B = 8'h28; #100;
A = 8'hFD; B = 8'h29; #100;
A = 8'hFD; B = 8'h2A; #100;
A = 8'hFD; B = 8'h2B; #100;
A = 8'hFD; B = 8'h2C; #100;
A = 8'hFD; B = 8'h2D; #100;
A = 8'hFD; B = 8'h2E; #100;
A = 8'hFD; B = 8'h2F; #100;
A = 8'hFD; B = 8'h30; #100;
A = 8'hFD; B = 8'h31; #100;
A = 8'hFD; B = 8'h32; #100;
A = 8'hFD; B = 8'h33; #100;
A = 8'hFD; B = 8'h34; #100;
A = 8'hFD; B = 8'h35; #100;
A = 8'hFD; B = 8'h36; #100;
A = 8'hFD; B = 8'h37; #100;
A = 8'hFD; B = 8'h38; #100;
A = 8'hFD; B = 8'h39; #100;
A = 8'hFD; B = 8'h3A; #100;
A = 8'hFD; B = 8'h3B; #100;
A = 8'hFD; B = 8'h3C; #100;
A = 8'hFD; B = 8'h3D; #100;
A = 8'hFD; B = 8'h3E; #100;
A = 8'hFD; B = 8'h3F; #100;
A = 8'hFD; B = 8'h40; #100;
A = 8'hFD; B = 8'h41; #100;
A = 8'hFD; B = 8'h42; #100;
A = 8'hFD; B = 8'h43; #100;
A = 8'hFD; B = 8'h44; #100;
A = 8'hFD; B = 8'h45; #100;
A = 8'hFD; B = 8'h46; #100;
A = 8'hFD; B = 8'h47; #100;
A = 8'hFD; B = 8'h48; #100;
A = 8'hFD; B = 8'h49; #100;
A = 8'hFD; B = 8'h4A; #100;
A = 8'hFD; B = 8'h4B; #100;
A = 8'hFD; B = 8'h4C; #100;
A = 8'hFD; B = 8'h4D; #100;
A = 8'hFD; B = 8'h4E; #100;
A = 8'hFD; B = 8'h4F; #100;
A = 8'hFD; B = 8'h50; #100;
A = 8'hFD; B = 8'h51; #100;
A = 8'hFD; B = 8'h52; #100;
A = 8'hFD; B = 8'h53; #100;
A = 8'hFD; B = 8'h54; #100;
A = 8'hFD; B = 8'h55; #100;
A = 8'hFD; B = 8'h56; #100;
A = 8'hFD; B = 8'h57; #100;
A = 8'hFD; B = 8'h58; #100;
A = 8'hFD; B = 8'h59; #100;
A = 8'hFD; B = 8'h5A; #100;
A = 8'hFD; B = 8'h5B; #100;
A = 8'hFD; B = 8'h5C; #100;
A = 8'hFD; B = 8'h5D; #100;
A = 8'hFD; B = 8'h5E; #100;
A = 8'hFD; B = 8'h5F; #100;
A = 8'hFD; B = 8'h60; #100;
A = 8'hFD; B = 8'h61; #100;
A = 8'hFD; B = 8'h62; #100;
A = 8'hFD; B = 8'h63; #100;
A = 8'hFD; B = 8'h64; #100;
A = 8'hFD; B = 8'h65; #100;
A = 8'hFD; B = 8'h66; #100;
A = 8'hFD; B = 8'h67; #100;
A = 8'hFD; B = 8'h68; #100;
A = 8'hFD; B = 8'h69; #100;
A = 8'hFD; B = 8'h6A; #100;
A = 8'hFD; B = 8'h6B; #100;
A = 8'hFD; B = 8'h6C; #100;
A = 8'hFD; B = 8'h6D; #100;
A = 8'hFD; B = 8'h6E; #100;
A = 8'hFD; B = 8'h6F; #100;
A = 8'hFD; B = 8'h70; #100;
A = 8'hFD; B = 8'h71; #100;
A = 8'hFD; B = 8'h72; #100;
A = 8'hFD; B = 8'h73; #100;
A = 8'hFD; B = 8'h74; #100;
A = 8'hFD; B = 8'h75; #100;
A = 8'hFD; B = 8'h76; #100;
A = 8'hFD; B = 8'h77; #100;
A = 8'hFD; B = 8'h78; #100;
A = 8'hFD; B = 8'h79; #100;
A = 8'hFD; B = 8'h7A; #100;
A = 8'hFD; B = 8'h7B; #100;
A = 8'hFD; B = 8'h7C; #100;
A = 8'hFD; B = 8'h7D; #100;
A = 8'hFD; B = 8'h7E; #100;
A = 8'hFD; B = 8'h7F; #100;
A = 8'hFD; B = 8'h80; #100;
A = 8'hFD; B = 8'h81; #100;
A = 8'hFD; B = 8'h82; #100;
A = 8'hFD; B = 8'h83; #100;
A = 8'hFD; B = 8'h84; #100;
A = 8'hFD; B = 8'h85; #100;
A = 8'hFD; B = 8'h86; #100;
A = 8'hFD; B = 8'h87; #100;
A = 8'hFD; B = 8'h88; #100;
A = 8'hFD; B = 8'h89; #100;
A = 8'hFD; B = 8'h8A; #100;
A = 8'hFD; B = 8'h8B; #100;
A = 8'hFD; B = 8'h8C; #100;
A = 8'hFD; B = 8'h8D; #100;
A = 8'hFD; B = 8'h8E; #100;
A = 8'hFD; B = 8'h8F; #100;
A = 8'hFD; B = 8'h90; #100;
A = 8'hFD; B = 8'h91; #100;
A = 8'hFD; B = 8'h92; #100;
A = 8'hFD; B = 8'h93; #100;
A = 8'hFD; B = 8'h94; #100;
A = 8'hFD; B = 8'h95; #100;
A = 8'hFD; B = 8'h96; #100;
A = 8'hFD; B = 8'h97; #100;
A = 8'hFD; B = 8'h98; #100;
A = 8'hFD; B = 8'h99; #100;
A = 8'hFD; B = 8'h9A; #100;
A = 8'hFD; B = 8'h9B; #100;
A = 8'hFD; B = 8'h9C; #100;
A = 8'hFD; B = 8'h9D; #100;
A = 8'hFD; B = 8'h9E; #100;
A = 8'hFD; B = 8'h9F; #100;
A = 8'hFD; B = 8'hA0; #100;
A = 8'hFD; B = 8'hA1; #100;
A = 8'hFD; B = 8'hA2; #100;
A = 8'hFD; B = 8'hA3; #100;
A = 8'hFD; B = 8'hA4; #100;
A = 8'hFD; B = 8'hA5; #100;
A = 8'hFD; B = 8'hA6; #100;
A = 8'hFD; B = 8'hA7; #100;
A = 8'hFD; B = 8'hA8; #100;
A = 8'hFD; B = 8'hA9; #100;
A = 8'hFD; B = 8'hAA; #100;
A = 8'hFD; B = 8'hAB; #100;
A = 8'hFD; B = 8'hAC; #100;
A = 8'hFD; B = 8'hAD; #100;
A = 8'hFD; B = 8'hAE; #100;
A = 8'hFD; B = 8'hAF; #100;
A = 8'hFD; B = 8'hB0; #100;
A = 8'hFD; B = 8'hB1; #100;
A = 8'hFD; B = 8'hB2; #100;
A = 8'hFD; B = 8'hB3; #100;
A = 8'hFD; B = 8'hB4; #100;
A = 8'hFD; B = 8'hB5; #100;
A = 8'hFD; B = 8'hB6; #100;
A = 8'hFD; B = 8'hB7; #100;
A = 8'hFD; B = 8'hB8; #100;
A = 8'hFD; B = 8'hB9; #100;
A = 8'hFD; B = 8'hBA; #100;
A = 8'hFD; B = 8'hBB; #100;
A = 8'hFD; B = 8'hBC; #100;
A = 8'hFD; B = 8'hBD; #100;
A = 8'hFD; B = 8'hBE; #100;
A = 8'hFD; B = 8'hBF; #100;
A = 8'hFD; B = 8'hC0; #100;
A = 8'hFD; B = 8'hC1; #100;
A = 8'hFD; B = 8'hC2; #100;
A = 8'hFD; B = 8'hC3; #100;
A = 8'hFD; B = 8'hC4; #100;
A = 8'hFD; B = 8'hC5; #100;
A = 8'hFD; B = 8'hC6; #100;
A = 8'hFD; B = 8'hC7; #100;
A = 8'hFD; B = 8'hC8; #100;
A = 8'hFD; B = 8'hC9; #100;
A = 8'hFD; B = 8'hCA; #100;
A = 8'hFD; B = 8'hCB; #100;
A = 8'hFD; B = 8'hCC; #100;
A = 8'hFD; B = 8'hCD; #100;
A = 8'hFD; B = 8'hCE; #100;
A = 8'hFD; B = 8'hCF; #100;
A = 8'hFD; B = 8'hD0; #100;
A = 8'hFD; B = 8'hD1; #100;
A = 8'hFD; B = 8'hD2; #100;
A = 8'hFD; B = 8'hD3; #100;
A = 8'hFD; B = 8'hD4; #100;
A = 8'hFD; B = 8'hD5; #100;
A = 8'hFD; B = 8'hD6; #100;
A = 8'hFD; B = 8'hD7; #100;
A = 8'hFD; B = 8'hD8; #100;
A = 8'hFD; B = 8'hD9; #100;
A = 8'hFD; B = 8'hDA; #100;
A = 8'hFD; B = 8'hDB; #100;
A = 8'hFD; B = 8'hDC; #100;
A = 8'hFD; B = 8'hDD; #100;
A = 8'hFD; B = 8'hDE; #100;
A = 8'hFD; B = 8'hDF; #100;
A = 8'hFD; B = 8'hE0; #100;
A = 8'hFD; B = 8'hE1; #100;
A = 8'hFD; B = 8'hE2; #100;
A = 8'hFD; B = 8'hE3; #100;
A = 8'hFD; B = 8'hE4; #100;
A = 8'hFD; B = 8'hE5; #100;
A = 8'hFD; B = 8'hE6; #100;
A = 8'hFD; B = 8'hE7; #100;
A = 8'hFD; B = 8'hE8; #100;
A = 8'hFD; B = 8'hE9; #100;
A = 8'hFD; B = 8'hEA; #100;
A = 8'hFD; B = 8'hEB; #100;
A = 8'hFD; B = 8'hEC; #100;
A = 8'hFD; B = 8'hED; #100;
A = 8'hFD; B = 8'hEE; #100;
A = 8'hFD; B = 8'hEF; #100;
A = 8'hFD; B = 8'hF0; #100;
A = 8'hFD; B = 8'hF1; #100;
A = 8'hFD; B = 8'hF2; #100;
A = 8'hFD; B = 8'hF3; #100;
A = 8'hFD; B = 8'hF4; #100;
A = 8'hFD; B = 8'hF5; #100;
A = 8'hFD; B = 8'hF6; #100;
A = 8'hFD; B = 8'hF7; #100;
A = 8'hFD; B = 8'hF8; #100;
A = 8'hFD; B = 8'hF9; #100;
A = 8'hFD; B = 8'hFA; #100;
A = 8'hFD; B = 8'hFB; #100;
A = 8'hFD; B = 8'hFC; #100;
A = 8'hFD; B = 8'hFD; #100;
A = 8'hFD; B = 8'hFE; #100;
A = 8'hFD; B = 8'hFF; #100;
A = 8'hFE; B = 8'h0; #100;
A = 8'hFE; B = 8'h1; #100;
A = 8'hFE; B = 8'h2; #100;
A = 8'hFE; B = 8'h3; #100;
A = 8'hFE; B = 8'h4; #100;
A = 8'hFE; B = 8'h5; #100;
A = 8'hFE; B = 8'h6; #100;
A = 8'hFE; B = 8'h7; #100;
A = 8'hFE; B = 8'h8; #100;
A = 8'hFE; B = 8'h9; #100;
A = 8'hFE; B = 8'hA; #100;
A = 8'hFE; B = 8'hB; #100;
A = 8'hFE; B = 8'hC; #100;
A = 8'hFE; B = 8'hD; #100;
A = 8'hFE; B = 8'hE; #100;
A = 8'hFE; B = 8'hF; #100;
A = 8'hFE; B = 8'h10; #100;
A = 8'hFE; B = 8'h11; #100;
A = 8'hFE; B = 8'h12; #100;
A = 8'hFE; B = 8'h13; #100;
A = 8'hFE; B = 8'h14; #100;
A = 8'hFE; B = 8'h15; #100;
A = 8'hFE; B = 8'h16; #100;
A = 8'hFE; B = 8'h17; #100;
A = 8'hFE; B = 8'h18; #100;
A = 8'hFE; B = 8'h19; #100;
A = 8'hFE; B = 8'h1A; #100;
A = 8'hFE; B = 8'h1B; #100;
A = 8'hFE; B = 8'h1C; #100;
A = 8'hFE; B = 8'h1D; #100;
A = 8'hFE; B = 8'h1E; #100;
A = 8'hFE; B = 8'h1F; #100;
A = 8'hFE; B = 8'h20; #100;
A = 8'hFE; B = 8'h21; #100;
A = 8'hFE; B = 8'h22; #100;
A = 8'hFE; B = 8'h23; #100;
A = 8'hFE; B = 8'h24; #100;
A = 8'hFE; B = 8'h25; #100;
A = 8'hFE; B = 8'h26; #100;
A = 8'hFE; B = 8'h27; #100;
A = 8'hFE; B = 8'h28; #100;
A = 8'hFE; B = 8'h29; #100;
A = 8'hFE; B = 8'h2A; #100;
A = 8'hFE; B = 8'h2B; #100;
A = 8'hFE; B = 8'h2C; #100;
A = 8'hFE; B = 8'h2D; #100;
A = 8'hFE; B = 8'h2E; #100;
A = 8'hFE; B = 8'h2F; #100;
A = 8'hFE; B = 8'h30; #100;
A = 8'hFE; B = 8'h31; #100;
A = 8'hFE; B = 8'h32; #100;
A = 8'hFE; B = 8'h33; #100;
A = 8'hFE; B = 8'h34; #100;
A = 8'hFE; B = 8'h35; #100;
A = 8'hFE; B = 8'h36; #100;
A = 8'hFE; B = 8'h37; #100;
A = 8'hFE; B = 8'h38; #100;
A = 8'hFE; B = 8'h39; #100;
A = 8'hFE; B = 8'h3A; #100;
A = 8'hFE; B = 8'h3B; #100;
A = 8'hFE; B = 8'h3C; #100;
A = 8'hFE; B = 8'h3D; #100;
A = 8'hFE; B = 8'h3E; #100;
A = 8'hFE; B = 8'h3F; #100;
A = 8'hFE; B = 8'h40; #100;
A = 8'hFE; B = 8'h41; #100;
A = 8'hFE; B = 8'h42; #100;
A = 8'hFE; B = 8'h43; #100;
A = 8'hFE; B = 8'h44; #100;
A = 8'hFE; B = 8'h45; #100;
A = 8'hFE; B = 8'h46; #100;
A = 8'hFE; B = 8'h47; #100;
A = 8'hFE; B = 8'h48; #100;
A = 8'hFE; B = 8'h49; #100;
A = 8'hFE; B = 8'h4A; #100;
A = 8'hFE; B = 8'h4B; #100;
A = 8'hFE; B = 8'h4C; #100;
A = 8'hFE; B = 8'h4D; #100;
A = 8'hFE; B = 8'h4E; #100;
A = 8'hFE; B = 8'h4F; #100;
A = 8'hFE; B = 8'h50; #100;
A = 8'hFE; B = 8'h51; #100;
A = 8'hFE; B = 8'h52; #100;
A = 8'hFE; B = 8'h53; #100;
A = 8'hFE; B = 8'h54; #100;
A = 8'hFE; B = 8'h55; #100;
A = 8'hFE; B = 8'h56; #100;
A = 8'hFE; B = 8'h57; #100;
A = 8'hFE; B = 8'h58; #100;
A = 8'hFE; B = 8'h59; #100;
A = 8'hFE; B = 8'h5A; #100;
A = 8'hFE; B = 8'h5B; #100;
A = 8'hFE; B = 8'h5C; #100;
A = 8'hFE; B = 8'h5D; #100;
A = 8'hFE; B = 8'h5E; #100;
A = 8'hFE; B = 8'h5F; #100;
A = 8'hFE; B = 8'h60; #100;
A = 8'hFE; B = 8'h61; #100;
A = 8'hFE; B = 8'h62; #100;
A = 8'hFE; B = 8'h63; #100;
A = 8'hFE; B = 8'h64; #100;
A = 8'hFE; B = 8'h65; #100;
A = 8'hFE; B = 8'h66; #100;
A = 8'hFE; B = 8'h67; #100;
A = 8'hFE; B = 8'h68; #100;
A = 8'hFE; B = 8'h69; #100;
A = 8'hFE; B = 8'h6A; #100;
A = 8'hFE; B = 8'h6B; #100;
A = 8'hFE; B = 8'h6C; #100;
A = 8'hFE; B = 8'h6D; #100;
A = 8'hFE; B = 8'h6E; #100;
A = 8'hFE; B = 8'h6F; #100;
A = 8'hFE; B = 8'h70; #100;
A = 8'hFE; B = 8'h71; #100;
A = 8'hFE; B = 8'h72; #100;
A = 8'hFE; B = 8'h73; #100;
A = 8'hFE; B = 8'h74; #100;
A = 8'hFE; B = 8'h75; #100;
A = 8'hFE; B = 8'h76; #100;
A = 8'hFE; B = 8'h77; #100;
A = 8'hFE; B = 8'h78; #100;
A = 8'hFE; B = 8'h79; #100;
A = 8'hFE; B = 8'h7A; #100;
A = 8'hFE; B = 8'h7B; #100;
A = 8'hFE; B = 8'h7C; #100;
A = 8'hFE; B = 8'h7D; #100;
A = 8'hFE; B = 8'h7E; #100;
A = 8'hFE; B = 8'h7F; #100;
A = 8'hFE; B = 8'h80; #100;
A = 8'hFE; B = 8'h81; #100;
A = 8'hFE; B = 8'h82; #100;
A = 8'hFE; B = 8'h83; #100;
A = 8'hFE; B = 8'h84; #100;
A = 8'hFE; B = 8'h85; #100;
A = 8'hFE; B = 8'h86; #100;
A = 8'hFE; B = 8'h87; #100;
A = 8'hFE; B = 8'h88; #100;
A = 8'hFE; B = 8'h89; #100;
A = 8'hFE; B = 8'h8A; #100;
A = 8'hFE; B = 8'h8B; #100;
A = 8'hFE; B = 8'h8C; #100;
A = 8'hFE; B = 8'h8D; #100;
A = 8'hFE; B = 8'h8E; #100;
A = 8'hFE; B = 8'h8F; #100;
A = 8'hFE; B = 8'h90; #100;
A = 8'hFE; B = 8'h91; #100;
A = 8'hFE; B = 8'h92; #100;
A = 8'hFE; B = 8'h93; #100;
A = 8'hFE; B = 8'h94; #100;
A = 8'hFE; B = 8'h95; #100;
A = 8'hFE; B = 8'h96; #100;
A = 8'hFE; B = 8'h97; #100;
A = 8'hFE; B = 8'h98; #100;
A = 8'hFE; B = 8'h99; #100;
A = 8'hFE; B = 8'h9A; #100;
A = 8'hFE; B = 8'h9B; #100;
A = 8'hFE; B = 8'h9C; #100;
A = 8'hFE; B = 8'h9D; #100;
A = 8'hFE; B = 8'h9E; #100;
A = 8'hFE; B = 8'h9F; #100;
A = 8'hFE; B = 8'hA0; #100;
A = 8'hFE; B = 8'hA1; #100;
A = 8'hFE; B = 8'hA2; #100;
A = 8'hFE; B = 8'hA3; #100;
A = 8'hFE; B = 8'hA4; #100;
A = 8'hFE; B = 8'hA5; #100;
A = 8'hFE; B = 8'hA6; #100;
A = 8'hFE; B = 8'hA7; #100;
A = 8'hFE; B = 8'hA8; #100;
A = 8'hFE; B = 8'hA9; #100;
A = 8'hFE; B = 8'hAA; #100;
A = 8'hFE; B = 8'hAB; #100;
A = 8'hFE; B = 8'hAC; #100;
A = 8'hFE; B = 8'hAD; #100;
A = 8'hFE; B = 8'hAE; #100;
A = 8'hFE; B = 8'hAF; #100;
A = 8'hFE; B = 8'hB0; #100;
A = 8'hFE; B = 8'hB1; #100;
A = 8'hFE; B = 8'hB2; #100;
A = 8'hFE; B = 8'hB3; #100;
A = 8'hFE; B = 8'hB4; #100;
A = 8'hFE; B = 8'hB5; #100;
A = 8'hFE; B = 8'hB6; #100;
A = 8'hFE; B = 8'hB7; #100;
A = 8'hFE; B = 8'hB8; #100;
A = 8'hFE; B = 8'hB9; #100;
A = 8'hFE; B = 8'hBA; #100;
A = 8'hFE; B = 8'hBB; #100;
A = 8'hFE; B = 8'hBC; #100;
A = 8'hFE; B = 8'hBD; #100;
A = 8'hFE; B = 8'hBE; #100;
A = 8'hFE; B = 8'hBF; #100;
A = 8'hFE; B = 8'hC0; #100;
A = 8'hFE; B = 8'hC1; #100;
A = 8'hFE; B = 8'hC2; #100;
A = 8'hFE; B = 8'hC3; #100;
A = 8'hFE; B = 8'hC4; #100;
A = 8'hFE; B = 8'hC5; #100;
A = 8'hFE; B = 8'hC6; #100;
A = 8'hFE; B = 8'hC7; #100;
A = 8'hFE; B = 8'hC8; #100;
A = 8'hFE; B = 8'hC9; #100;
A = 8'hFE; B = 8'hCA; #100;
A = 8'hFE; B = 8'hCB; #100;
A = 8'hFE; B = 8'hCC; #100;
A = 8'hFE; B = 8'hCD; #100;
A = 8'hFE; B = 8'hCE; #100;
A = 8'hFE; B = 8'hCF; #100;
A = 8'hFE; B = 8'hD0; #100;
A = 8'hFE; B = 8'hD1; #100;
A = 8'hFE; B = 8'hD2; #100;
A = 8'hFE; B = 8'hD3; #100;
A = 8'hFE; B = 8'hD4; #100;
A = 8'hFE; B = 8'hD5; #100;
A = 8'hFE; B = 8'hD6; #100;
A = 8'hFE; B = 8'hD7; #100;
A = 8'hFE; B = 8'hD8; #100;
A = 8'hFE; B = 8'hD9; #100;
A = 8'hFE; B = 8'hDA; #100;
A = 8'hFE; B = 8'hDB; #100;
A = 8'hFE; B = 8'hDC; #100;
A = 8'hFE; B = 8'hDD; #100;
A = 8'hFE; B = 8'hDE; #100;
A = 8'hFE; B = 8'hDF; #100;
A = 8'hFE; B = 8'hE0; #100;
A = 8'hFE; B = 8'hE1; #100;
A = 8'hFE; B = 8'hE2; #100;
A = 8'hFE; B = 8'hE3; #100;
A = 8'hFE; B = 8'hE4; #100;
A = 8'hFE; B = 8'hE5; #100;
A = 8'hFE; B = 8'hE6; #100;
A = 8'hFE; B = 8'hE7; #100;
A = 8'hFE; B = 8'hE8; #100;
A = 8'hFE; B = 8'hE9; #100;
A = 8'hFE; B = 8'hEA; #100;
A = 8'hFE; B = 8'hEB; #100;
A = 8'hFE; B = 8'hEC; #100;
A = 8'hFE; B = 8'hED; #100;
A = 8'hFE; B = 8'hEE; #100;
A = 8'hFE; B = 8'hEF; #100;
A = 8'hFE; B = 8'hF0; #100;
A = 8'hFE; B = 8'hF1; #100;
A = 8'hFE; B = 8'hF2; #100;
A = 8'hFE; B = 8'hF3; #100;
A = 8'hFE; B = 8'hF4; #100;
A = 8'hFE; B = 8'hF5; #100;
A = 8'hFE; B = 8'hF6; #100;
A = 8'hFE; B = 8'hF7; #100;
A = 8'hFE; B = 8'hF8; #100;
A = 8'hFE; B = 8'hF9; #100;
A = 8'hFE; B = 8'hFA; #100;
A = 8'hFE; B = 8'hFB; #100;
A = 8'hFE; B = 8'hFC; #100;
A = 8'hFE; B = 8'hFD; #100;
A = 8'hFE; B = 8'hFE; #100;
A = 8'hFE; B = 8'hFF; #100;
A = 8'hFF; B = 8'h0; #100;
A = 8'hFF; B = 8'h1; #100;
A = 8'hFF; B = 8'h2; #100;
A = 8'hFF; B = 8'h3; #100;
A = 8'hFF; B = 8'h4; #100;
A = 8'hFF; B = 8'h5; #100;
A = 8'hFF; B = 8'h6; #100;
A = 8'hFF; B = 8'h7; #100;
A = 8'hFF; B = 8'h8; #100;
A = 8'hFF; B = 8'h9; #100;
A = 8'hFF; B = 8'hA; #100;
A = 8'hFF; B = 8'hB; #100;
A = 8'hFF; B = 8'hC; #100;
A = 8'hFF; B = 8'hD; #100;
A = 8'hFF; B = 8'hE; #100;
A = 8'hFF; B = 8'hF; #100;
A = 8'hFF; B = 8'h10; #100;
A = 8'hFF; B = 8'h11; #100;
A = 8'hFF; B = 8'h12; #100;
A = 8'hFF; B = 8'h13; #100;
A = 8'hFF; B = 8'h14; #100;
A = 8'hFF; B = 8'h15; #100;
A = 8'hFF; B = 8'h16; #100;
A = 8'hFF; B = 8'h17; #100;
A = 8'hFF; B = 8'h18; #100;
A = 8'hFF; B = 8'h19; #100;
A = 8'hFF; B = 8'h1A; #100;
A = 8'hFF; B = 8'h1B; #100;
A = 8'hFF; B = 8'h1C; #100;
A = 8'hFF; B = 8'h1D; #100;
A = 8'hFF; B = 8'h1E; #100;
A = 8'hFF; B = 8'h1F; #100;
A = 8'hFF; B = 8'h20; #100;
A = 8'hFF; B = 8'h21; #100;
A = 8'hFF; B = 8'h22; #100;
A = 8'hFF; B = 8'h23; #100;
A = 8'hFF; B = 8'h24; #100;
A = 8'hFF; B = 8'h25; #100;
A = 8'hFF; B = 8'h26; #100;
A = 8'hFF; B = 8'h27; #100;
A = 8'hFF; B = 8'h28; #100;
A = 8'hFF; B = 8'h29; #100;
A = 8'hFF; B = 8'h2A; #100;
A = 8'hFF; B = 8'h2B; #100;
A = 8'hFF; B = 8'h2C; #100;
A = 8'hFF; B = 8'h2D; #100;
A = 8'hFF; B = 8'h2E; #100;
A = 8'hFF; B = 8'h2F; #100;
A = 8'hFF; B = 8'h30; #100;
A = 8'hFF; B = 8'h31; #100;
A = 8'hFF; B = 8'h32; #100;
A = 8'hFF; B = 8'h33; #100;
A = 8'hFF; B = 8'h34; #100;
A = 8'hFF; B = 8'h35; #100;
A = 8'hFF; B = 8'h36; #100;
A = 8'hFF; B = 8'h37; #100;
A = 8'hFF; B = 8'h38; #100;
A = 8'hFF; B = 8'h39; #100;
A = 8'hFF; B = 8'h3A; #100;
A = 8'hFF; B = 8'h3B; #100;
A = 8'hFF; B = 8'h3C; #100;
A = 8'hFF; B = 8'h3D; #100;
A = 8'hFF; B = 8'h3E; #100;
A = 8'hFF; B = 8'h3F; #100;
A = 8'hFF; B = 8'h40; #100;
A = 8'hFF; B = 8'h41; #100;
A = 8'hFF; B = 8'h42; #100;
A = 8'hFF; B = 8'h43; #100;
A = 8'hFF; B = 8'h44; #100;
A = 8'hFF; B = 8'h45; #100;
A = 8'hFF; B = 8'h46; #100;
A = 8'hFF; B = 8'h47; #100;
A = 8'hFF; B = 8'h48; #100;
A = 8'hFF; B = 8'h49; #100;
A = 8'hFF; B = 8'h4A; #100;
A = 8'hFF; B = 8'h4B; #100;
A = 8'hFF; B = 8'h4C; #100;
A = 8'hFF; B = 8'h4D; #100;
A = 8'hFF; B = 8'h4E; #100;
A = 8'hFF; B = 8'h4F; #100;
A = 8'hFF; B = 8'h50; #100;
A = 8'hFF; B = 8'h51; #100;
A = 8'hFF; B = 8'h52; #100;
A = 8'hFF; B = 8'h53; #100;
A = 8'hFF; B = 8'h54; #100;
A = 8'hFF; B = 8'h55; #100;
A = 8'hFF; B = 8'h56; #100;
A = 8'hFF; B = 8'h57; #100;
A = 8'hFF; B = 8'h58; #100;
A = 8'hFF; B = 8'h59; #100;
A = 8'hFF; B = 8'h5A; #100;
A = 8'hFF; B = 8'h5B; #100;
A = 8'hFF; B = 8'h5C; #100;
A = 8'hFF; B = 8'h5D; #100;
A = 8'hFF; B = 8'h5E; #100;
A = 8'hFF; B = 8'h5F; #100;
A = 8'hFF; B = 8'h60; #100;
A = 8'hFF; B = 8'h61; #100;
A = 8'hFF; B = 8'h62; #100;
A = 8'hFF; B = 8'h63; #100;
A = 8'hFF; B = 8'h64; #100;
A = 8'hFF; B = 8'h65; #100;
A = 8'hFF; B = 8'h66; #100;
A = 8'hFF; B = 8'h67; #100;
A = 8'hFF; B = 8'h68; #100;
A = 8'hFF; B = 8'h69; #100;
A = 8'hFF; B = 8'h6A; #100;
A = 8'hFF; B = 8'h6B; #100;
A = 8'hFF; B = 8'h6C; #100;
A = 8'hFF; B = 8'h6D; #100;
A = 8'hFF; B = 8'h6E; #100;
A = 8'hFF; B = 8'h6F; #100;
A = 8'hFF; B = 8'h70; #100;
A = 8'hFF; B = 8'h71; #100;
A = 8'hFF; B = 8'h72; #100;
A = 8'hFF; B = 8'h73; #100;
A = 8'hFF; B = 8'h74; #100;
A = 8'hFF; B = 8'h75; #100;
A = 8'hFF; B = 8'h76; #100;
A = 8'hFF; B = 8'h77; #100;
A = 8'hFF; B = 8'h78; #100;
A = 8'hFF; B = 8'h79; #100;
A = 8'hFF; B = 8'h7A; #100;
A = 8'hFF; B = 8'h7B; #100;
A = 8'hFF; B = 8'h7C; #100;
A = 8'hFF; B = 8'h7D; #100;
A = 8'hFF; B = 8'h7E; #100;
A = 8'hFF; B = 8'h7F; #100;
A = 8'hFF; B = 8'h80; #100;
A = 8'hFF; B = 8'h81; #100;
A = 8'hFF; B = 8'h82; #100;
A = 8'hFF; B = 8'h83; #100;
A = 8'hFF; B = 8'h84; #100;
A = 8'hFF; B = 8'h85; #100;
A = 8'hFF; B = 8'h86; #100;
A = 8'hFF; B = 8'h87; #100;
A = 8'hFF; B = 8'h88; #100;
A = 8'hFF; B = 8'h89; #100;
A = 8'hFF; B = 8'h8A; #100;
A = 8'hFF; B = 8'h8B; #100;
A = 8'hFF; B = 8'h8C; #100;
A = 8'hFF; B = 8'h8D; #100;
A = 8'hFF; B = 8'h8E; #100;
A = 8'hFF; B = 8'h8F; #100;
A = 8'hFF; B = 8'h90; #100;
A = 8'hFF; B = 8'h91; #100;
A = 8'hFF; B = 8'h92; #100;
A = 8'hFF; B = 8'h93; #100;
A = 8'hFF; B = 8'h94; #100;
A = 8'hFF; B = 8'h95; #100;
A = 8'hFF; B = 8'h96; #100;
A = 8'hFF; B = 8'h97; #100;
A = 8'hFF; B = 8'h98; #100;
A = 8'hFF; B = 8'h99; #100;
A = 8'hFF; B = 8'h9A; #100;
A = 8'hFF; B = 8'h9B; #100;
A = 8'hFF; B = 8'h9C; #100;
A = 8'hFF; B = 8'h9D; #100;
A = 8'hFF; B = 8'h9E; #100;
A = 8'hFF; B = 8'h9F; #100;
A = 8'hFF; B = 8'hA0; #100;
A = 8'hFF; B = 8'hA1; #100;
A = 8'hFF; B = 8'hA2; #100;
A = 8'hFF; B = 8'hA3; #100;
A = 8'hFF; B = 8'hA4; #100;
A = 8'hFF; B = 8'hA5; #100;
A = 8'hFF; B = 8'hA6; #100;
A = 8'hFF; B = 8'hA7; #100;
A = 8'hFF; B = 8'hA8; #100;
A = 8'hFF; B = 8'hA9; #100;
A = 8'hFF; B = 8'hAA; #100;
A = 8'hFF; B = 8'hAB; #100;
A = 8'hFF; B = 8'hAC; #100;
A = 8'hFF; B = 8'hAD; #100;
A = 8'hFF; B = 8'hAE; #100;
A = 8'hFF; B = 8'hAF; #100;
A = 8'hFF; B = 8'hB0; #100;
A = 8'hFF; B = 8'hB1; #100;
A = 8'hFF; B = 8'hB2; #100;
A = 8'hFF; B = 8'hB3; #100;
A = 8'hFF; B = 8'hB4; #100;
A = 8'hFF; B = 8'hB5; #100;
A = 8'hFF; B = 8'hB6; #100;
A = 8'hFF; B = 8'hB7; #100;
A = 8'hFF; B = 8'hB8; #100;
A = 8'hFF; B = 8'hB9; #100;
A = 8'hFF; B = 8'hBA; #100;
A = 8'hFF; B = 8'hBB; #100;
A = 8'hFF; B = 8'hBC; #100;
A = 8'hFF; B = 8'hBD; #100;
A = 8'hFF; B = 8'hBE; #100;
A = 8'hFF; B = 8'hBF; #100;
A = 8'hFF; B = 8'hC0; #100;
A = 8'hFF; B = 8'hC1; #100;
A = 8'hFF; B = 8'hC2; #100;
A = 8'hFF; B = 8'hC3; #100;
A = 8'hFF; B = 8'hC4; #100;
A = 8'hFF; B = 8'hC5; #100;
A = 8'hFF; B = 8'hC6; #100;
A = 8'hFF; B = 8'hC7; #100;
A = 8'hFF; B = 8'hC8; #100;
A = 8'hFF; B = 8'hC9; #100;
A = 8'hFF; B = 8'hCA; #100;
A = 8'hFF; B = 8'hCB; #100;
A = 8'hFF; B = 8'hCC; #100;
A = 8'hFF; B = 8'hCD; #100;
A = 8'hFF; B = 8'hCE; #100;
A = 8'hFF; B = 8'hCF; #100;
A = 8'hFF; B = 8'hD0; #100;
A = 8'hFF; B = 8'hD1; #100;
A = 8'hFF; B = 8'hD2; #100;
A = 8'hFF; B = 8'hD3; #100;
A = 8'hFF; B = 8'hD4; #100;
A = 8'hFF; B = 8'hD5; #100;
A = 8'hFF; B = 8'hD6; #100;
A = 8'hFF; B = 8'hD7; #100;
A = 8'hFF; B = 8'hD8; #100;
A = 8'hFF; B = 8'hD9; #100;
A = 8'hFF; B = 8'hDA; #100;
A = 8'hFF; B = 8'hDB; #100;
A = 8'hFF; B = 8'hDC; #100;
A = 8'hFF; B = 8'hDD; #100;
A = 8'hFF; B = 8'hDE; #100;
A = 8'hFF; B = 8'hDF; #100;
A = 8'hFF; B = 8'hE0; #100;
A = 8'hFF; B = 8'hE1; #100;
A = 8'hFF; B = 8'hE2; #100;
A = 8'hFF; B = 8'hE3; #100;
A = 8'hFF; B = 8'hE4; #100;
A = 8'hFF; B = 8'hE5; #100;
A = 8'hFF; B = 8'hE6; #100;
A = 8'hFF; B = 8'hE7; #100;
A = 8'hFF; B = 8'hE8; #100;
A = 8'hFF; B = 8'hE9; #100;
A = 8'hFF; B = 8'hEA; #100;
A = 8'hFF; B = 8'hEB; #100;
A = 8'hFF; B = 8'hEC; #100;
A = 8'hFF; B = 8'hED; #100;
A = 8'hFF; B = 8'hEE; #100;
A = 8'hFF; B = 8'hEF; #100;
A = 8'hFF; B = 8'hF0; #100;
A = 8'hFF; B = 8'hF1; #100;
A = 8'hFF; B = 8'hF2; #100;
A = 8'hFF; B = 8'hF3; #100;
A = 8'hFF; B = 8'hF4; #100;
A = 8'hFF; B = 8'hF5; #100;
A = 8'hFF; B = 8'hF6; #100;
A = 8'hFF; B = 8'hF7; #100;
A = 8'hFF; B = 8'hF8; #100;
A = 8'hFF; B = 8'hF9; #100;
A = 8'hFF; B = 8'hFA; #100;
A = 8'hFF; B = 8'hFB; #100;
A = 8'hFF; B = 8'hFC; #100;
A = 8'hFF; B = 8'hFD; #100;
A = 8'hFF; B = 8'hFE; #100;
A = 8'hFF; B = 8'hFF; #100;

	$stop;
end


endmodule 
