*
.MODEL CMOSN NMOS (                                LEVEL   = 49
+VERSION = 3.1            TNOM    = 27             TOX     = 1.41E-8
+XJ      = 1.5E-7         NCH     = 1.7E17         VTH0    = 0.6033055
+K1      = 0.9193622      K2      = -0.1065538     K3      = 20.591979
+K3B     = -9.1011155     W0      = 4.393248E-8    NLX     = 1.426577E-9
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 0.8628177      DVT1    = 0.4045315      DVT2    = -0.5
+U0      = 455.6568715    UA      = 1E-13          UB      = 1.383698E-18
+UC      = 8.07605E-12    VSAT    = 1.97155E5      A0      = 0.5976138
+AGS     = 0.1289087      B0      = 2.029789E-6    B1      = 5E-6
+KETA    = -2.756238E-3   A1      = 2.328154E-4    A2      = 0.3
+RDSW    = 1.074553E3     PRWG    = 0.0988607      PRWB    = 7.238942E-3
+WR      = 1              WINT    = 1.965107E-7    LINT    = 8.377083E-8
+XL      = 1E-7           XW      = 0              DWG     = -8.437034E-9
+DWB     = 3.078094E-8    VOFF    = -7.633973E-5   NFACTOR = 1.1573034
+CIT     = 0              CDSC    = 2.4E-4         CDSCD   = 0
+CDSCB   = 0              ETA0    = 3.231837E-3    ETAB    = 4.803812E-3
+DSUB    = 0.0537894      PCLM    = 2.1073222      PDIBLC1 = 4.117691E-4
+PDIBLC2 = 1.173409E-3    PDIBLCB = -0.2714521     DROUT   = 2.514784E-4
+PSCBE1  = 2.167284E10    PSCBE2  = 4.309903E-9    PVAG    = 0
+DELTA   = 0.01           RSH     = 84.3           MOBMOD  = 1
+PRT     = 0              UTE     = -1.5           KT1     = -0.11
+KT1L    = 0              KT2     = 0.022          UA1     = 4.31E-9
+UB1     = -7.61E-18      UC1     = -5.6E-11       AT      = 3.3E4
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 1.82E-10       CGSO    = 1.82E-10       CGBO    = 1E-9
+CJ      = 4.175598E-4    PB      = 0.840291       MJ      = 0.4297322
+CJSW    = 3.483931E-10   PBSW    = 0.8            MJSW    = 0.2059566
+CJSWG   = 1.64E-10       PBSWG   = 0.8            MJSWG   = 0.2059566
+CF      = 0              PVTH0   = -0.0505758     PRDSW   = 281.2200286
+PK2     = -0.0697499     WKETA   = -6.123851E-3   LKETA   = -2.318372E-3    )
*
.MODEL CMOSP PMOS (                                LEVEL   = 49
+VERSION = 3.1            TNOM    = 27             TOX     = 1.41E-8
+XJ      = 1.5E-7         NCH     = 1.7E17         VTH0    = -0.9152268
+K1      = 0.553472       K2      = 7.871921E-3    K3      = 8.3456329
+K3B     = 0.8137476      W0      = 1E-8           NLX     = 1.661298E-7
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 0.6826241      DVT1    = 0.2907764      DVT2    = -0.3
+U0      = 201.3603195    UA      = 2.408572E-9    UB      = 1E-21
+UC      = -1E-10         VSAT    = 1.043844E5     A0      = 0.8625012
+AGS     = 0.097008       B0      = 5.131287E-7    B1      = 0
+KETA    = -4.865785E-3   A1      = 4.099078E-4    A2      = 0.5220155
+RDSW    = 3E3            PRWG    = -0.0260778     PRWB    = -0.0514886
+WR      = 1              WINT    = 2.224208E-7    LINT    = 1.277363E-7
+XL      = 1E-7           XW      = 0              DWG     = 1.017918E-11
+DWB     = -2.133914E-8   VOFF    = -0.0728335     NFACTOR = 1.0000003
+CIT     = 0              CDSC    = 2.4E-4         CDSCD   = 0
+CDSCB   = 0              ETA0    = 0              ETAB    = -0.0178415
+DSUB    = 0.3875471      PCLM    = 2.4913442      PDIBLC1 = 0.0335017
+PDIBLC2 = 3.071184E-3    PDIBLCB = 0.0157585      DROUT   = 0.1973195
+PSCBE1  = 1E8            PSCBE2  = 3.383681E-9    PVAG    = 0.0150059
+DELTA   = 0.01           RSH     = 107.7          MOBMOD  = 1
+PRT     = 0              UTE     = -1.5           KT1     = -0.11
+KT1L    = 0              KT2     = 0.022          UA1     = 4.31E-9
+UB1     = -7.61E-18      UC1     = -5.6E-11       AT      = 3.3E4
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 2.35E-10       CGSO    = 2.35E-10       CGBO    = 1E-9
+CJ      = 7.137225E-4    PB      = 0.8741848      MJ      = 0.4883246
+CJSW    = 2.425711E-10   PBSW    = 0.8            MJSW    = 0.2079833
+CJSWG   = 6.4E-11        PBSWG   = 0.8            MJSWG   = 0.2079833
+CF      = 0              PVTH0   = 5.98016E-3     PRDSW   = 14.8598424
+PK2     = 3.73981E-3     WKETA   = 7.275123E-3    LKETA   = 0.0298866       )
*
