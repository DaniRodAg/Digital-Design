
`timescale 1ns/1ps

module FA_16B_TB();

reg[15:0] A, B;
wire[15:0] S;
wire Cout;
wire Cin = 1'b0;

FA_16B duv
(
	.A(A),
	.B(B),
	.S(S),
	
	.Cin(Cin),
	.Cout(Cout)
);

initial
begin
A = 16'h0000; B = 16'h0000; #100;
A = 16'h0000; B = 16'h0001; #100;
A = 16'h0000; B = 16'h0002; #100;
A = 16'h0000; B = 16'h0003; #100;
A = 16'h0000; B = 16'h0004; #100;
A = 16'h0000; B = 16'h0005; #100;
A = 16'h0000; B = 16'h0006; #100;
A = 16'h0000; B = 16'h0007; #100;
A = 16'h0000; B = 16'h0008; #100;
A = 16'h0000; B = 16'h0009; #100;
A = 16'h0000; B = 16'h000A; #100;
A = 16'h0000; B = 16'h000B; #100;
A = 16'h0000; B = 16'h000C; #100;
A = 16'h0000; B = 16'h000D; #100;
A = 16'h0000; B = 16'h000E; #100;
A = 16'h0000; B = 16'h000F; #100;
A = 16'h0000; B = 16'h0010; #100;
A = 16'h0000; B = 16'h0011; #100;
A = 16'h0000; B = 16'h0012; #100;
A = 16'h0000; B = 16'h0013; #100;
A = 16'h0000; B = 16'h0014; #100;
A = 16'h0000; B = 16'h0015; #100;
A = 16'h0000; B = 16'h0016; #100;
A = 16'h0000; B = 16'h0017; #100;
A = 16'h0000; B = 16'h0018; #100;
A = 16'h0000; B = 16'h0019; #100;
A = 16'h0000; B = 16'h001A; #100;
A = 16'h0000; B = 16'h001B; #100;
A = 16'h0000; B = 16'h001C; #100;
A = 16'h0000; B = 16'h001D; #100;
A = 16'h0000; B = 16'h001E; #100;
A = 16'h0000; B = 16'h001F; #100;
A = 16'h0000; B = 16'h0020; #100;
A = 16'h0000; B = 16'h0021; #100;
A = 16'h0000; B = 16'h0022; #100;
A = 16'h0000; B = 16'h0023; #100;
A = 16'h0000; B = 16'h0024; #100;
A = 16'h0000; B = 16'h0025; #100;
A = 16'h0000; B = 16'h0026; #100;
A = 16'h0000; B = 16'h0027; #100;
A = 16'h0000; B = 16'h0028; #100;
A = 16'h0000; B = 16'h0029; #100;
A = 16'h0000; B = 16'h002A; #100;
A = 16'h0000; B = 16'h002B; #100;
A = 16'h0000; B = 16'h002C; #100;
A = 16'h0000; B = 16'h002D; #100;
A = 16'h0000; B = 16'h002E; #100;
A = 16'h0000; B = 16'h002F; #100;
A = 16'h0000; B = 16'h0030; #100;
A = 16'h0000; B = 16'h0031; #100;
A = 16'h0000; B = 16'h0032; #100;
A = 16'h0000; B = 16'h0033; #100;
A = 16'h0000; B = 16'h0034; #100;
A = 16'h0000; B = 16'h0035; #100;
A = 16'h0000; B = 16'h0036; #100;
A = 16'h0000; B = 16'h0037; #100;
A = 16'h0000; B = 16'h0038; #100;
A = 16'h0000; B = 16'h0039; #100;
A = 16'h0000; B = 16'h003A; #100;
A = 16'h0000; B = 16'h003B; #100;
A = 16'h0000; B = 16'h003C; #100;
A = 16'h0000; B = 16'h003D; #100;
A = 16'h0000; B = 16'h003E; #100;
A = 16'h0000; B = 16'h003F; #100;
A = 16'h0000; B = 16'h0040; #100;
A = 16'h0000; B = 16'h0041; #100;
A = 16'h0000; B = 16'h0042; #100;
A = 16'h000; B = 16'h0043; #100;
A = 16'h000; B = 16'h0044; #100;
A = 16'h000; B = 16'h0045; #100;
A = 16'h000; B = 16'h0046; #100;
A = 16'h000; B = 16'h0047; #100;
A = 16'h000; B = 16'h0048; #100;
A = 16'h000; B = 16'h0049; #100;
A = 16'h000; B = 16'h004A; #100;
A = 16'h000; B = 16'h004B; #100;
A = 16'h000; B = 16'h004C; #100;
A = 16'h000; B = 16'h004D; #100;
A = 16'h000; B = 16'h004E; #100;
A = 16'h000; B = 16'h004F; #100;
A = 16'h000; B = 16'h0050; #100;
A = 16'h000; B = 16'h0051; #100;
A = 16'h000; B = 16'h0052; #100;
A = 16'h000; B = 16'h0053; #100;
A = 16'h000; B = 16'h0054; #100;
A = 16'h000; B = 16'h0055; #100;
A = 16'h000; B = 16'h0056; #100;
A = 16'h000; B = 16'h0057; #100;
A = 16'h000; B = 16'h0058; #100;
A = 16'h000; B = 16'h0059; #100;
A = 16'h000; B = 16'h005A; #100;
A = 16'h000; B = 16'h005B; #100;
A = 16'h000; B = 16'h005C; #100;
A = 16'h000; B = 16'h005D; #100;
A = 16'h000; B = 16'h005E; #100;
A = 16'h000; B = 16'h005F; #100;
A = 16'h000; B = 16'h0060; #100;
A = 16'h000; B = 16'h0061; #100;
A = 16'h000; B = 16'h0062; #100;
A = 16'h000; B = 16'h0063; #100;
A = 16'h000; B = 16'h0064; #100;
A = 16'h000; B = 16'h0065; #100;
A = 16'h000; B = 16'h0066; #100;
A = 16'h000; B = 16'h0067; #100;
A = 16'h000; B = 16'h0068; #100;
A = 16'h000; B = 16'h0069; #100;
A = 16'h000; B = 16'h006A; #100;
A = 16'h000; B = 16'h006B; #100;
A = 16'h000; B = 16'h006C; #100;
A = 16'h000; B = 16'h006D; #100;
A = 16'h000; B = 16'h006E; #100;
A = 16'h000; B = 16'h006F; #100;
A = 16'h000; B = 16'h0070; #100;
A = 16'h000; B = 16'h0071; #100;
A = 16'h000; B = 16'h0072; #100;
A = 16'h000; B = 16'h0073; #100;
A = 16'h000; B = 16'h0074; #100;
A = 16'h000; B = 16'h0075; #100;
A = 16'h000; B = 16'h0076; #100;
A = 16'h000; B = 16'h0077; #100;
A = 16'h000; B = 16'h0078; #100;
A = 16'h000; B = 16'h0079; #100;
A = 16'h000; B = 16'h007A; #100;
A = 16'h000; B = 16'h007B; #100;
A = 16'h000; B = 16'h007C; #100;
A = 16'h000; B = 16'h007D; #100;
A = 16'h000; B = 16'h007E; #100;
A = 16'h000; B = 16'h007F; #100;
A = 16'h000; B = 16'h0080; #100;
A = 16'h000; B = 16'h0081; #100;
A = 16'h000; B = 16'h0082; #100;
A = 16'h000; B = 16'h0083; #100;
A = 16'h000; B = 16'h0084; #100;
A = 16'h000; B = 16'h0085; #100;
A = 16'h000; B = 16'h0086; #100;
A = 16'h000; B = 16'h0087; #100;
A = 16'h000; B = 16'h0088; #100;
A = 16'h000; B = 16'h0089; #100;
A = 16'h000; B = 16'h008A; #100;
A = 16'h000; B = 16'h008B; #100;
A = 16'h000; B = 16'h008C; #100;
A = 16'h000; B = 16'h008D; #100;
A = 16'h000; B = 16'h008E; #100;
A = 16'h000; B = 16'h008F; #100;
A = 16'h000; B = 16'h0090; #100;
A = 16'h000; B = 16'h0091; #100;
A = 16'h000; B = 16'h0092; #100;
A = 16'h000; B = 16'h0093; #100;
A = 16'h000; B = 16'h0094; #100;
A = 16'h000; B = 16'h0095; #100;
A = 16'h000; B = 16'h0096; #100;
A = 16'h000; B = 16'h0097; #100;
A = 16'h000; B = 16'h0098; #100;
A = 16'h000; B = 16'h0099; #100;
A = 16'h000; B = 16'h009A; #100;
A = 16'h000; B = 16'h009B; #100;
A = 16'h000; B = 16'h009C; #100;
A = 16'h000; B = 16'h009D; #100;
A = 16'h000; B = 16'h009E; #100;
A = 16'h000; B = 16'h009F; #100;
A = 16'h000; B = 16'h00A0; #100;
A = 16'h000; B = 16'h00A1; #100;
A = 16'h000; B = 16'h00A2; #100;
A = 16'h000; B = 16'h00A3; #100;
A = 16'h000; B = 16'h00A4; #100;
A = 16'h000; B = 16'h00A5; #100;
A = 16'h000; B = 16'h00A6; #100;
A = 16'h000; B = 16'h00A7; #100;
A = 16'h000; B = 16'h00A8; #100;
A = 16'h000; B = 16'h00A9; #100;
A = 16'h000; B = 16'h00AA; #100;
A = 16'h000; B = 16'h00AB; #100;
A = 16'h000; B = 16'h00AC; #100;
A = 16'h000; B = 16'h00AD; #100;
A = 16'h000; B = 16'h00AE; #100;
A = 16'h000; B = 16'h00AF; #100;
A = 16'h000; B = 16'h00B0; #100;
A = 16'h000; B = 16'h00B1; #100;
A = 16'h000; B = 16'h00B2; #100;
A = 16'h000; B = 16'h00B3; #100;
A = 16'h000; B = 16'h00B4; #100;
A = 16'h000; B = 16'h00B5; #100;
A = 16'h000; B = 16'h00B6; #100;
A = 16'h000; B = 16'h00B7; #100;
A = 16'h000; B = 16'h00B8; #100;
A = 16'h000; B = 16'h00B9; #100;
A = 16'h000; B = 16'h00BA; #100;
A = 16'h000; B = 16'h00BB; #100;
A = 16'h000; B = 16'h00BC; #100;
A = 16'h000; B = 16'h00BD; #100;
A = 16'h000; B = 16'h00BE; #100;
A = 16'h000; B = 16'h00BF; #100;
A = 16'h000; B = 16'h00C0; #100;
A = 16'h000; B = 16'h00C1; #100;
A = 16'h000; B = 16'h00C2; #100;
A = 16'h000; B = 16'h00C3; #100;
A = 16'h000; B = 16'h00C4; #100;
A = 16'h000; B = 16'h00C5; #100;
A = 16'h000; B = 16'h00C6; #100;
A = 16'h000; B = 16'h00C7; #100;
A = 16'h000; B = 16'h00C8; #100;
A = 16'h000; B = 16'h00C9; #100;
A = 16'h000; B = 16'h00CA; #100;
A = 16'h000; B = 16'h00CB; #100;
A = 16'h000; B = 16'h00CC; #100;
A = 16'h000; B = 16'h00CD; #100;
A = 16'h000; B = 16'h00CE; #100;
A = 16'h000; B = 16'h00CF; #100;
A = 16'h000; B = 16'h00D0; #100;
A = 16'h000; B = 16'h00D1; #100;
A = 16'h000; B = 16'h00D2; #100;
A = 16'h000; B = 16'h00D3; #100;
A = 16'h000; B = 16'h00D4; #100;
A = 16'h000; B = 16'h00D5; #100;
A = 16'h000; B = 16'h00D6; #100;
A = 16'h000; B = 16'h00D7; #100;
A = 16'h000; B = 16'h00D8; #100;
A = 16'h000; B = 16'h00D9; #100;
A = 16'h000; B = 16'h00DA; #100;
A = 16'h000; B = 16'h00DB; #100;
A = 16'h000; B = 16'h00DC; #100;
A = 16'h000; B = 16'h00DD; #100;
A = 16'h000; B = 16'h00DE; #100;
A = 16'h000; B = 16'h00DF; #100;
A = 16'h000; B = 16'h00E0; #100;
A = 16'h000; B = 16'h00E1; #100;
A = 16'h000; B = 16'h00E2; #100;
A = 16'h000; B = 16'h00E3; #100;
A = 16'h000; B = 16'h00E4; #100;
A = 16'h000; B = 16'h00E5; #100;
A = 16'h000; B = 16'h00E6; #100;
A = 16'h000; B = 16'h00E7; #100;
A = 16'h000; B = 16'h00E8; #100;
A = 16'h000; B = 16'h00E9; #100;
A = 16'h000; B = 16'h00EA; #100;
A = 16'h000; B = 16'h00EB; #100;
A = 16'h000; B = 16'h00EC; #100;
A = 16'h000; B = 16'h00ED; #100;
A = 16'h000; B = 16'h00EE; #100;
A = 16'h000; B = 16'h00EF; #100;
A = 16'h000; B = 16'h00F0; #100;
A = 16'h000; B = 16'h00F1; #100;
A = 16'h000; B = 16'h00F2; #100;
A = 16'h000; B = 16'h00F3; #100;
A = 16'h000; B = 16'h00F4; #100;
A = 16'h000; B = 16'h00F5; #100;
A = 16'h000; B = 16'h00F6; #100;
A = 16'h000; B = 16'h00F7; #100;
A = 16'h000; B = 16'h00F8; #100;
A = 16'h000; B = 16'h00F9; #100;
A = 16'h000; B = 16'h00FA; #100;
A = 16'h000; B = 16'h00FB; #100;
A = 16'h000; B = 16'h00FC; #100;
A = 16'h000; B = 16'h00FD; #100;
A = 16'h000; B = 16'h00FE; #100;
A = 16'h000; B = 16'h00FF; #100;
A = 16'h001; B = 16'h000; #100;
A = 16'h001; B = 16'h001; #100;
A = 16'h001; B = 16'h002; #100;
A = 16'h001; B = 16'h003; #100;
A = 16'h001; B = 16'h004; #100;
A = 16'h001; B = 16'h005; #100;
A = 16'h001; B = 16'h006; #100;
A = 16'h001; B = 16'h007; #100;
A = 16'h001; B = 16'h008; #100;
A = 16'h001; B = 16'h009; #100;
A = 16'h001; B = 16'h00A; #100;
A = 16'h001; B = 16'h00B; #100;
A = 16'h001; B = 16'h00C; #100;
A = 16'h001; B = 16'h00D; #100;
A = 16'h001; B = 16'h00E; #100;
A = 16'h001; B = 16'h00F; #100;
A = 16'h001; B = 16'h0010; #100;
A = 16'h001; B = 16'h0011; #100;
A = 16'h001; B = 16'h0012; #100;
A = 16'h001; B = 16'h0013; #100;
A = 16'h001; B = 16'h0014; #100;
A = 16'h001; B = 16'h0015; #100;
A = 16'h001; B = 16'h0016; #100;
A = 16'h001; B = 16'h0017; #100;
A = 16'h001; B = 16'h0018; #100;
A = 16'h001; B = 16'h0019; #100;
A = 16'h001; B = 16'h001A; #100;
A = 16'h001; B = 16'h001B; #100;
A = 16'h001; B = 16'h001C; #100;
A = 16'h001; B = 16'h001D; #100;
A = 16'h001; B = 16'h001E; #100;
A = 16'h001; B = 16'h001F; #100;
A = 16'h001; B = 16'h0020; #100;
A = 16'h001; B = 16'h0021; #100;
A = 16'h001; B = 16'h0022; #100;
A = 16'h001; B = 16'h0023; #100;
A = 16'h001; B = 16'h0024; #100;
A = 16'h001; B = 16'h0025; #100;
A = 16'h001; B = 16'h0026; #100;
A = 16'h001; B = 16'h0027; #100;
A = 16'h001; B = 16'h0028; #100;
A = 16'h001; B = 16'h0029; #100;
A = 16'h001; B = 16'h002A; #100;
A = 16'h001; B = 16'h002B; #100;
A = 16'h001; B = 16'h002C; #100;
A = 16'h001; B = 16'h002D; #100;
A = 16'h001; B = 16'h002E; #100;
A = 16'h001; B = 16'h002F; #100;
A = 16'h001; B = 16'h0030; #100;
A = 16'h001; B = 16'h0031; #100;
A = 16'h001; B = 16'h0032; #100;
A = 16'h001; B = 16'h0033; #100;
A = 16'h001; B = 16'h0034; #100;
A = 16'h001; B = 16'h0035; #100;
A = 16'h001; B = 16'h0036; #100;
A = 16'h001; B = 16'h0037; #100;
A = 16'h001; B = 16'h0038; #100;
A = 16'h001; B = 16'h0039; #100;
A = 16'h001; B = 16'h003A; #100;
A = 16'h001; B = 16'h003B; #100;
A = 16'h001; B = 16'h003C; #100;
A = 16'h001; B = 16'h003D; #100;
A = 16'h001; B = 16'h003E; #100;
A = 16'h001; B = 16'h003F; #100;
A = 16'h001; B = 16'h0040; #100;
A = 16'h001; B = 16'h0041; #100;
A = 16'h001; B = 16'h0042; #100;
A = 16'h001; B = 16'h0043; #100;
A = 16'h001; B = 16'h0044; #100;
A = 16'h001; B = 16'h0045; #100;
A = 16'h001; B = 16'h0046; #100;
A = 16'h001; B = 16'h0047; #100;
A = 16'h001; B = 16'h0048; #100;
A = 16'h001; B = 16'h0049; #100;
A = 16'h001; B = 16'h004A; #100;
A = 16'h001; B = 16'h004B; #100;
A = 16'h001; B = 16'h004C; #100;
A = 16'h001; B = 16'h004D; #100;
A = 16'h001; B = 16'h004E; #100;
A = 16'h001; B = 16'h004F; #100;
A = 16'h001; B = 16'h0050; #100;
A = 16'h001; B = 16'h0051; #100;
A = 16'h001; B = 16'h0052; #100;
A = 16'h001; B = 16'h0053; #100;
A = 16'h001; B = 16'h0054; #100;
A = 16'h001; B = 16'h0055; #100;
A = 16'h001; B = 16'h0056; #100;
A = 16'h001; B = 16'h0057; #100;
A = 16'h001; B = 16'h0058; #100;
A = 16'h001; B = 16'h0059; #100;
A = 16'h001; B = 16'h005A; #100;
A = 16'h001; B = 16'h005B; #100;
A = 16'h001; B = 16'h005C; #100;
A = 16'h001; B = 16'h005D; #100;
A = 16'h001; B = 16'h005E; #100;
A = 16'h001; B = 16'h005F; #100;
A = 16'h001; B = 16'h0060; #100;
A = 16'h001; B = 16'h0061; #100;
A = 16'h001; B = 16'h0062; #100;
A = 16'h001; B = 16'h0063; #100;
A = 16'h001; B = 16'h0064; #100;
A = 16'h001; B = 16'h0065; #100;
A = 16'h001; B = 16'h0066; #100;
A = 16'h001; B = 16'h0067; #100;
A = 16'h001; B = 16'h0068; #100;
A = 16'h001; B = 16'h0069; #100;
A = 16'h001; B = 16'h006A; #100;
A = 16'h001; B = 16'h006B; #100;
A = 16'h001; B = 16'h006C; #100;
A = 16'h001; B = 16'h006D; #100;
A = 16'h001; B = 16'h006E; #100;
A = 16'h001; B = 16'h006F; #100;
A = 16'h001; B = 16'h0070; #100;
A = 16'h001; B = 16'h0071; #100;
A = 16'h001; B = 16'h0072; #100;
A = 16'h001; B = 16'h0073; #100;
A = 16'h001; B = 16'h0074; #100;
A = 16'h001; B = 16'h0075; #100;
A = 16'h001; B = 16'h0076; #100;
A = 16'h001; B = 16'h0077; #100;
A = 16'h001; B = 16'h0078; #100;
A = 16'h001; B = 16'h0079; #100;
A = 16'h001; B = 16'h007A; #100;
A = 16'h001; B = 16'h007B; #100;
A = 16'h001; B = 16'h007C; #100;
A = 16'h001; B = 16'h007D; #100;
A = 16'h001; B = 16'h007E; #100;
A = 16'h001; B = 16'h007F; #100;
A = 16'h001; B = 16'h0080; #100;
A = 16'h001; B = 16'h0081; #100;
A = 16'h001; B = 16'h0082; #100;
A = 16'h001; B = 16'h0083; #100;
A = 16'h001; B = 16'h0084; #100;
A = 16'h001; B = 16'h0085; #100;
A = 16'h001; B = 16'h0086; #100;
A = 16'h001; B = 16'h0087; #100;
A = 16'h001; B = 16'h0088; #100;
A = 16'h001; B = 16'h0089; #100;
A = 16'h001; B = 16'h008A; #100;
A = 16'h001; B = 16'h008B; #100;
A = 16'h001; B = 16'h008C; #100;
A = 16'h001; B = 16'h008D; #100;
A = 16'h001; B = 16'h008E; #100;
A = 16'h001; B = 16'h008F; #100;
A = 16'h001; B = 16'h0090; #100;
A = 16'h001; B = 16'h0091; #100;
A = 16'h001; B = 16'h0092; #100;
A = 16'h001; B = 16'h0093; #100;
A = 16'h001; B = 16'h0094; #100;
A = 16'h001; B = 16'h0095; #100;
A = 16'h001; B = 16'h0096; #100;
A = 16'h001; B = 16'h0097; #100;
A = 16'h001; B = 16'h0098; #100;
A = 16'h001; B = 16'h0099; #100;
A = 16'h001; B = 16'h009A; #100;
A = 16'h001; B = 16'h009B; #100;
A = 16'h001; B = 16'h009C; #100;
A = 16'h001; B = 16'h009D; #100;
A = 16'h001; B = 16'h009E; #100;
A = 16'h001; B = 16'h009F; #100;
A = 16'h001; B = 16'h00A0; #100;
A = 16'h001; B = 16'h00A1; #100;
A = 16'h001; B = 16'h00A2; #100;
A = 16'h001; B = 16'h00A3; #100;
A = 16'h001; B = 16'h00A4; #100;
A = 16'h001; B = 16'h00A5; #100;
A = 16'h001; B = 16'h00A6; #100;
A = 16'h001; B = 16'h00A7; #100;
A = 16'h001; B = 16'h00A8; #100;
A = 16'h001; B = 16'h00A9; #100;
A = 16'h001; B = 16'h00AA; #100;
A = 16'h001; B = 16'h00AB; #100;
A = 16'h001; B = 16'h00AC; #100;
A = 16'h001; B = 16'h00AD; #100;
A = 16'h001; B = 16'h00AE; #100;
A = 16'h001; B = 16'h00AF; #100;
A = 16'h001; B = 16'h00B0; #100;
A = 16'h001; B = 16'h00B1; #100;
A = 16'h001; B = 16'h00B2; #100;
A = 16'h001; B = 16'h00B3; #100;
A = 16'h001; B = 16'h00B4; #100;
A = 16'h001; B = 16'h00B5; #100;
A = 16'h001; B = 16'h00B6; #100;
A = 16'h001; B = 16'h00B7; #100;
A = 16'h001; B = 16'h00B8; #100;
A = 16'h001; B = 16'h00B9; #100;
A = 16'h001; B = 16'h00BA; #100;
A = 16'h001; B = 16'h00BB; #100;
A = 16'h001; B = 16'h00BC; #100;
A = 16'h001; B = 16'h00BD; #100;
A = 16'h001; B = 16'h00BE; #100;
A = 16'h001; B = 16'h00BF; #100;
A = 16'h001; B = 16'h00C0; #100;
A = 16'h001; B = 16'h00C1; #100;
A = 16'h001; B = 16'h00C2; #100;
A = 16'h001; B = 16'h00C3; #100;
A = 16'h001; B = 16'h00C4; #100;
A = 16'h001; B = 16'h00C5; #100;
A = 16'h001; B = 16'h00C6; #100;
A = 16'h001; B = 16'h00C7; #100;
A = 16'h001; B = 16'h00C8; #100;
A = 16'h001; B = 16'h00C9; #100;
A = 16'h001; B = 16'h00CA; #100;
A = 16'h001; B = 16'h00CB; #100;
A = 16'h001; B = 16'h00CC; #100;
A = 16'h001; B = 16'h00CD; #100;
A = 16'h001; B = 16'h00CE; #100;
A = 16'h001; B = 16'h00CF; #100;
A = 16'h001; B = 16'h00D0; #100;
A = 16'h001; B = 16'h00D1; #100;
A = 16'h001; B = 16'h00D2; #100;
A = 16'h001; B = 16'h00D3; #100;
A = 16'h001; B = 16'h00D4; #100;
A = 16'h001; B = 16'h00D5; #100;
A = 16'h001; B = 16'h00D6; #100;
A = 16'h001; B = 16'h00D7; #100;
A = 16'h001; B = 16'h00D8; #100;
A = 16'h001; B = 16'h00D9; #100;
A = 16'h001; B = 16'h00DA; #100;
A = 16'h001; B = 16'h00DB; #100;
A = 16'h001; B = 16'h00DC; #100;
A = 16'h001; B = 16'h00DD; #100;
A = 16'h001; B = 16'h00DE; #100;
A = 16'h001; B = 16'h00DF; #100;
A = 16'h001; B = 16'h00E0; #100;
A = 16'h001; B = 16'h00E1; #100;
A = 16'h001; B = 16'h00E2; #100;
A = 16'h001; B = 16'h00E3; #100;
A = 16'h001; B = 16'h00E4; #100;
A = 16'h001; B = 16'h00E5; #100;
A = 16'h001; B = 16'h00E6; #100;
A = 16'h001; B = 16'h00E7; #100;
A = 16'h001; B = 16'h00E8; #100;
A = 16'h001; B = 16'h00E9; #100;
A = 16'h001; B = 16'h00EA; #100;
A = 16'h001; B = 16'h00EB; #100;
A = 16'h001; B = 16'h00EC; #100;
A = 16'h001; B = 16'h00ED; #100;
A = 16'h001; B = 16'h00EE; #100;
A = 16'h001; B = 16'h00EF; #100;
A = 16'h001; B = 16'h00F0; #100;
A = 16'h001; B = 16'h00F1; #100;
A = 16'h001; B = 16'h00F2; #100;
A = 16'h001; B = 16'h00F3; #100;
A = 16'h001; B = 16'h00F4; #100;
A = 16'h001; B = 16'h00F5; #100;
A = 16'h001; B = 16'h00F6; #100;
A = 16'h001; B = 16'h00F7; #100;
A = 16'h001; B = 16'h00F8; #100;
A = 16'h001; B = 16'h00F9; #100;
A = 16'h001; B = 16'h00FA; #100;
A = 16'h001; B = 16'h00FB; #100;
A = 16'h001; B = 16'h00FC; #100;
A = 16'h001; B = 16'h00FD; #100;
A = 16'h001; B = 16'h00FE; #100;
A = 16'h001; B = 16'h00FF; #100;
A = 16'h002; B = 16'h000; #100;
A = 16'h002; B = 16'h001; #100;
A = 16'h002; B = 16'h002; #100;
A = 16'h002; B = 16'h003; #100;
A = 16'h002; B = 16'h004; #100;
A = 16'h002; B = 16'h005; #100;
A = 16'h002; B = 16'h006; #100;
A = 16'h002; B = 16'h007; #100;
A = 16'h002; B = 16'h008; #100;
A = 16'h002; B = 16'h009; #100;
A = 16'h002; B = 16'h00A; #100;
A = 16'h002; B = 16'h00B; #100;
A = 16'h002; B = 16'h00C; #100;
A = 16'h002; B = 16'h00D; #100;
A = 16'h002; B = 16'h00E; #100;
A = 16'h002; B = 16'h00F; #100;
A = 16'h002; B = 16'h0010; #100;
A = 16'h002; B = 16'h0011; #100;
A = 16'h002; B = 16'h0012; #100;
A = 16'h002; B = 16'h0013; #100;
A = 16'h002; B = 16'h0014; #100;
A = 16'h002; B = 16'h0015; #100;
A = 16'h002; B = 16'h0016; #100;
A = 16'h002; B = 16'h0017; #100;
A = 16'h002; B = 16'h0018; #100;
A = 16'h002; B = 16'h0019; #100;
A = 16'h002; B = 16'h001A; #100;
A = 16'h002; B = 16'h001B; #100;
A = 16'h002; B = 16'h001C; #100;
A = 16'h002; B = 16'h001D; #100;
A = 16'h002; B = 16'h001E; #100;
A = 16'h002; B = 16'h001F; #100;
A = 16'h002; B = 16'h0020; #100;
A = 16'h002; B = 16'h0021; #100;
A = 16'h002; B = 16'h0022; #100;
A = 16'h002; B = 16'h0023; #100;
A = 16'h002; B = 16'h0024; #100;
A = 16'h002; B = 16'h0025; #100;
A = 16'h002; B = 16'h0026; #100;
A = 16'h002; B = 16'h0027; #100;
A = 16'h002; B = 16'h0028; #100;
A = 16'h002; B = 16'h0029; #100;
A = 16'h002; B = 16'h002A; #100;
A = 16'h002; B = 16'h002B; #100;
A = 16'h002; B = 16'h002C; #100;
A = 16'h002; B = 16'h002D; #100;
A = 16'h002; B = 16'h002E; #100;
A = 16'h002; B = 16'h002F; #100;
A = 16'h002; B = 16'h0030; #100;
A = 16'h002; B = 16'h0031; #100;
A = 16'h002; B = 16'h0032; #100;
A = 16'h002; B = 16'h0033; #100;
A = 16'h002; B = 16'h0034; #100;
A = 16'h002; B = 16'h0035; #100;
A = 16'h002; B = 16'h0036; #100;
A = 16'h002; B = 16'h0037; #100;
A = 16'h002; B = 16'h0038; #100;
A = 16'h002; B = 16'h0039; #100;
A = 16'h002; B = 16'h003A; #100;
A = 16'h002; B = 16'h003B; #100;
A = 16'h002; B = 16'h003C; #100;
A = 16'h002; B = 16'h003D; #100;
A = 16'h002; B = 16'h003E; #100;
A = 16'h002; B = 16'h003F; #100;
A = 16'h002; B = 16'h0040; #100;
A = 16'h002; B = 16'h0041; #100;
A = 16'h002; B = 16'h0042; #100;
A = 16'h002; B = 16'h0043; #100;
A = 16'h002; B = 16'h0044; #100;
A = 16'h002; B = 16'h0045; #100;
A = 16'h002; B = 16'h0046; #100;
A = 16'h002; B = 16'h0047; #100;
A = 16'h002; B = 16'h0048; #100;
A = 16'h002; B = 16'h0049; #100;
A = 16'h002; B = 16'h004A; #100;
A = 16'h002; B = 16'h004B; #100;
A = 16'h002; B = 16'h004C; #100;
A = 16'h002; B = 16'h004D; #100;
A = 16'h002; B = 16'h004E; #100;
A = 16'h002; B = 16'h004F; #100;
A = 16'h002; B = 16'h0050; #100;
A = 16'h002; B = 16'h0051; #100;
A = 16'h002; B = 16'h0052; #100;
A = 16'h002; B = 16'h0053; #100;
A = 16'h002; B = 16'h0054; #100;
A = 16'h002; B = 16'h0055; #100;
A = 16'h002; B = 16'h0056; #100;
A = 16'h002; B = 16'h0057; #100;
A = 16'h002; B = 16'h0058; #100;
A = 16'h002; B = 16'h0059; #100;
A = 16'h002; B = 16'h005A; #100;
A = 16'h002; B = 16'h005B; #100;
A = 16'h002; B = 16'h005C; #100;
A = 16'h002; B = 16'h005D; #100;
A = 16'h002; B = 16'h005E; #100;
A = 16'h002; B = 16'h005F; #100;
A = 16'h002; B = 16'h0060; #100;
A = 16'h002; B = 16'h0061; #100;
A = 16'h002; B = 16'h0062; #100;
A = 16'h002; B = 16'h0063; #100;
A = 16'h002; B = 16'h0064; #100;
A = 16'h002; B = 16'h0065; #100;
A = 16'h002; B = 16'h0066; #100;
A = 16'h002; B = 16'h0067; #100;
A = 16'h002; B = 16'h0068; #100;
A = 16'h002; B = 16'h0069; #100;
A = 16'h002; B = 16'h006A; #100;
A = 16'h002; B = 16'h006B; #100;
A = 16'h002; B = 16'h006C; #100;
A = 16'h002; B = 16'h006D; #100;
A = 16'h002; B = 16'h006E; #100;
A = 16'h002; B = 16'h006F; #100;
A = 16'h002; B = 16'h0070; #100;
A = 16'h002; B = 16'h0071; #100;
A = 16'h002; B = 16'h0072; #100;
A = 16'h002; B = 16'h0073; #100;
A = 16'h002; B = 16'h0074; #100;
A = 16'h002; B = 16'h0075; #100;
A = 16'h002; B = 16'h0076; #100;
A = 16'h002; B = 16'h0077; #100;
A = 16'h002; B = 16'h0078; #100;
A = 16'h002; B = 16'h0079; #100;
A = 16'h002; B = 16'h007A; #100;
A = 16'h002; B = 16'h007B; #100;
A = 16'h002; B = 16'h007C; #100;
A = 16'h002; B = 16'h007D; #100;
A = 16'h002; B = 16'h007E; #100;
A = 16'h002; B = 16'h007F; #100;
A = 16'h002; B = 16'h0080; #100;
A = 16'h002; B = 16'h0081; #100;
A = 16'h002; B = 16'h0082; #100;
A = 16'h002; B = 16'h0083; #100;
A = 16'h002; B = 16'h0084; #100;
A = 16'h002; B = 16'h0085; #100;
A = 16'h002; B = 16'h0086; #100;
A = 16'h002; B = 16'h0087; #100;
A = 16'h002; B = 16'h0088; #100;
A = 16'h002; B = 16'h0089; #100;
A = 16'h002; B = 16'h008A; #100;
A = 16'h002; B = 16'h008B; #100;
A = 16'h002; B = 16'h008C; #100;
A = 16'h002; B = 16'h008D; #100;
A = 16'h002; B = 16'h008E; #100;
A = 16'h002; B = 16'h008F; #100;
A = 16'h002; B = 16'h0090; #100;
A = 16'h002; B = 16'h0091; #100;
A = 16'h002; B = 16'h0092; #100;
A = 16'h002; B = 16'h0093; #100;
A = 16'h002; B = 16'h0094; #100;
A = 16'h002; B = 16'h0095; #100;
A = 16'h002; B = 16'h0096; #100;
A = 16'h002; B = 16'h0097; #100;
A = 16'h002; B = 16'h0098; #100;
A = 16'h002; B = 16'h0099; #100;
A = 16'h002; B = 16'h009A; #100;
A = 16'h002; B = 16'h009B; #100;
A = 16'h002; B = 16'h009C; #100;
A = 16'h002; B = 16'h009D; #100;
A = 16'h002; B = 16'h009E; #100;
A = 16'h002; B = 16'h009F; #100;
A = 16'h002; B = 16'h00A0; #100;
A = 16'h002; B = 16'h00A1; #100;
A = 16'h002; B = 16'h00A2; #100;
A = 16'h002; B = 16'h00A3; #100;
A = 16'h002; B = 16'h00A4; #100;
A = 16'h002; B = 16'h00A5; #100;
A = 16'h002; B = 16'h00A6; #100;
A = 16'h002; B = 16'h00A7; #100;
A = 16'h002; B = 16'h00A8; #100;
A = 16'h002; B = 16'h00A9; #100;
A = 16'h002; B = 16'h00AA; #100;
A = 16'h002; B = 16'h00AB; #100;
A = 16'h002; B = 16'h00AC; #100;
A = 16'h002; B = 16'h00AD; #100;
A = 16'h002; B = 16'h00AE; #100;
A = 16'h002; B = 16'h00AF; #100;
A = 16'h002; B = 16'h00B0; #100;
A = 16'h002; B = 16'h00B1; #100;
A = 16'h002; B = 16'h00B2; #100;
A = 16'h002; B = 16'h00B3; #100;
A = 16'h002; B = 16'h00B4; #100;
A = 16'h002; B = 16'h00B5; #100;
A = 16'h002; B = 16'h00B6; #100;
A = 16'h002; B = 16'h00B7; #100;
A = 16'h002; B = 16'h00B8; #100;
A = 16'h002; B = 16'h00B9; #100;
A = 16'h002; B = 16'h00BA; #100;
A = 16'h002; B = 16'h00BB; #100;
A = 16'h002; B = 16'h00BC; #100;
A = 16'h002; B = 16'h00BD; #100;
A = 16'h002; B = 16'h00BE; #100;
A = 16'h002; B = 16'h00BF; #100;
A = 16'h002; B = 16'h00C0; #100;
A = 16'h002; B = 16'h00C1; #100;
A = 16'h002; B = 16'h00C2; #100;
A = 16'h002; B = 16'h00C3; #100;
A = 16'h002; B = 16'h00C4; #100;
A = 16'h002; B = 16'h00C5; #100;
A = 16'h002; B = 16'h00C6; #100;
A = 16'h002; B = 16'h00C7; #100;
A = 16'h002; B = 16'h00C8; #100;
A = 16'h002; B = 16'h00C9; #100;
A = 16'h002; B = 16'h00CA; #100;
A = 16'h002; B = 16'h00CB; #100;
A = 16'h002; B = 16'h00CC; #100;
A = 16'h002; B = 16'h00CD; #100;
A = 16'h002; B = 16'h00CE; #100;
A = 16'h002; B = 16'h00CF; #100;
A = 16'h002; B = 16'h00D0; #100;
A = 16'h002; B = 16'h00D1; #100;
A = 16'h002; B = 16'h00D2; #100;
A = 16'h002; B = 16'h00D3; #100;
A = 16'h002; B = 16'h00D4; #100;
A = 16'h002; B = 16'h00D5; #100;
A = 16'h002; B = 16'h00D6; #100;
A = 16'h002; B = 16'h00D7; #100;
A = 16'h002; B = 16'h00D8; #100;
A = 16'h002; B = 16'h00D9; #100;
A = 16'h002; B = 16'h00DA; #100;
A = 16'h002; B = 16'h00DB; #100;
A = 16'h002; B = 16'h00DC; #100;
A = 16'h002; B = 16'h00DD; #100;
A = 16'h002; B = 16'h00DE; #100;
A = 16'h002; B = 16'h00DF; #100;
A = 16'h002; B = 16'h00E0; #100;
A = 16'h002; B = 16'h00E1; #100;
A = 16'h002; B = 16'h00E2; #100;
A = 16'h002; B = 16'h00E3; #100;
A = 16'h002; B = 16'h00E4; #100;
A = 16'h002; B = 16'h00E5; #100;
A = 16'h002; B = 16'h00E6; #100;
A = 16'h002; B = 16'h00E7; #100;
A = 16'h002; B = 16'h00E8; #100;
A = 16'h002; B = 16'h00E9; #100;
A = 16'h002; B = 16'h00EA; #100;
A = 16'h002; B = 16'h00EB; #100;
A = 16'h002; B = 16'h00EC; #100;
A = 16'h002; B = 16'h00ED; #100;
A = 16'h002; B = 16'h00EE; #100;
A = 16'h002; B = 16'h00EF; #100;
A = 16'h002; B = 16'h00F0; #100;
A = 16'h002; B = 16'h00F1; #100;
A = 16'h002; B = 16'h00F2; #100;
A = 16'h002; B = 16'h00F3; #100;
A = 16'h002; B = 16'h00F4; #100;
A = 16'h002; B = 16'h00F5; #100;
A = 16'h002; B = 16'h00F6; #100;
A = 16'h002; B = 16'h00F7; #100;
A = 16'h002; B = 16'h00F8; #100;
A = 16'h002; B = 16'h00F9; #100;
A = 16'h002; B = 16'h00FA; #100;
A = 16'h002; B = 16'h00FB; #100;
A = 16'h002; B = 16'h00FC; #100;
A = 16'h002; B = 16'h00FD; #100;
A = 16'h002; B = 16'h00FE; #100;
A = 16'h002; B = 16'h00FF; #100;
A = 16'h003; B = 16'h000; #100;
A = 16'h003; B = 16'h001; #100;
A = 16'h003; B = 16'h002; #100;
A = 16'h003; B = 16'h003; #100;
A = 16'h003; B = 16'h004; #100;
A = 16'h003; B = 16'h005; #100;
A = 16'h003; B = 16'h006; #100;
A = 16'h003; B = 16'h007; #100;
A = 16'h003; B = 16'h008; #100;
A = 16'h003; B = 16'h009; #100;
A = 16'h003; B = 16'h00A; #100;
A = 16'h003; B = 16'h00B; #100;
A = 16'h003; B = 16'h00C; #100;
A = 16'h003; B = 16'h00D; #100;
A = 16'h003; B = 16'h00E; #100;
A = 16'h003; B = 16'h00F; #100;
A = 16'h003; B = 16'h0010; #100;
A = 16'h003; B = 16'h0011; #100;
A = 16'h003; B = 16'h0012; #100;
A = 16'h003; B = 16'h0013; #100;
A = 16'h003; B = 16'h0014; #100;
A = 16'h003; B = 16'h0015; #100;
A = 16'h003; B = 16'h0016; #100;
A = 16'h003; B = 16'h0017; #100;
A = 16'h003; B = 16'h0018; #100;
A = 16'h003; B = 16'h0019; #100;
A = 16'h003; B = 16'h001A; #100;
A = 16'h003; B = 16'h001B; #100;
A = 16'h003; B = 16'h001C; #100;
A = 16'h003; B = 16'h001D; #100;
A = 16'h003; B = 16'h001E; #100;
A = 16'h003; B = 16'h001F; #100;
A = 16'h003; B = 16'h0020; #100;
A = 16'h003; B = 16'h0021; #100;
A = 16'h003; B = 16'h0022; #100;
A = 16'h003; B = 16'h0023; #100;
A = 16'h003; B = 16'h0024; #100;
A = 16'h003; B = 16'h0025; #100;
A = 16'h003; B = 16'h0026; #100;
A = 16'h003; B = 16'h0027; #100;
A = 16'h003; B = 16'h0028; #100;
A = 16'h003; B = 16'h0029; #100;
A = 16'h003; B = 16'h002A; #100;
A = 16'h003; B = 16'h002B; #100;
A = 16'h003; B = 16'h002C; #100;
A = 16'h003; B = 16'h002D; #100;
A = 16'h003; B = 16'h002E; #100;
A = 16'h003; B = 16'h002F; #100;
A = 16'h003; B = 16'h0030; #100;
A = 16'h003; B = 16'h0031; #100;
A = 16'h003; B = 16'h0032; #100;
A = 16'h003; B = 16'h0033; #100;
A = 16'h003; B = 16'h0034; #100;
A = 16'h003; B = 16'h0035; #100;
A = 16'h003; B = 16'h0036; #100;
A = 16'h003; B = 16'h0037; #100;
A = 16'h003; B = 16'h0038; #100;
A = 16'h003; B = 16'h0039; #100;
A = 16'h003; B = 16'h003A; #100;
A = 16'h003; B = 16'h003B; #100;
A = 16'h003; B = 16'h003C; #100;
A = 16'h003; B = 16'h003D; #100;
A = 16'h003; B = 16'h003E; #100;
A = 16'h003; B = 16'h003F; #100;
A = 16'h003; B = 16'h0040; #100;
A = 16'h003; B = 16'h0041; #100;
A = 16'h003; B = 16'h0042; #100;
A = 16'h003; B = 16'h0043; #100;
A = 16'h003; B = 16'h0044; #100;
A = 16'h003; B = 16'h0045; #100;
A = 16'h003; B = 16'h0046; #100;
A = 16'h003; B = 16'h0047; #100;
A = 16'h003; B = 16'h0048; #100;
A = 16'h003; B = 16'h0049; #100;
A = 16'h003; B = 16'h004A; #100;
A = 16'h003; B = 16'h004B; #100;
A = 16'h003; B = 16'h004C; #100;
A = 16'h003; B = 16'h004D; #100;
A = 16'h003; B = 16'h004E; #100;
A = 16'h003; B = 16'h004F; #100;
A = 16'h003; B = 16'h0050; #100;
A = 16'h003; B = 16'h0051; #100;
A = 16'h003; B = 16'h0052; #100;
A = 16'h003; B = 16'h0053; #100;
A = 16'h003; B = 16'h0054; #100;
A = 16'h003; B = 16'h0055; #100;
A = 16'h003; B = 16'h0056; #100;
A = 16'h003; B = 16'h0057; #100;
A = 16'h003; B = 16'h0058; #100;
A = 16'h003; B = 16'h0059; #100;
A = 16'h003; B = 16'h005A; #100;
A = 16'h003; B = 16'h005B; #100;
A = 16'h003; B = 16'h005C; #100;
A = 16'h003; B = 16'h005D; #100;
A = 16'h003; B = 16'h005E; #100;
A = 16'h003; B = 16'h005F; #100;
A = 16'h003; B = 16'h0060; #100;
A = 16'h003; B = 16'h0061; #100;
A = 16'h003; B = 16'h0062; #100;
A = 16'h003; B = 16'h0063; #100;
A = 16'h003; B = 16'h0064; #100;
A = 16'h003; B = 16'h0065; #100;
A = 16'h003; B = 16'h0066; #100;
A = 16'h003; B = 16'h0067; #100;
A = 16'h003; B = 16'h0068; #100;
A = 16'h003; B = 16'h0069; #100;
A = 16'h003; B = 16'h006A; #100;
A = 16'h003; B = 16'h006B; #100;
A = 16'h003; B = 16'h006C; #100;
A = 16'h003; B = 16'h006D; #100;
A = 16'h003; B = 16'h006E; #100;
A = 16'h003; B = 16'h006F; #100;
A = 16'h003; B = 16'h0070; #100;
A = 16'h003; B = 16'h0071; #100;
A = 16'h003; B = 16'h0072; #100;
A = 16'h003; B = 16'h0073; #100;
A = 16'h003; B = 16'h0074; #100;
A = 16'h003; B = 16'h0075; #100;
A = 16'h003; B = 16'h0076; #100;
A = 16'h003; B = 16'h0077; #100;
A = 16'h003; B = 16'h0078; #100;
A = 16'h003; B = 16'h0079; #100;
A = 16'h003; B = 16'h007A; #100;
A = 16'h003; B = 16'h007B; #100;
A = 16'h003; B = 16'h007C; #100;
A = 16'h003; B = 16'h007D; #100;
A = 16'h003; B = 16'h007E; #100;
A = 16'h003; B = 16'h007F; #100;
A = 16'h003; B = 16'h0080; #100;
A = 16'h003; B = 16'h0081; #100;
A = 16'h003; B = 16'h0082; #100;
A = 16'h003; B = 16'h0083; #100;
A = 16'h003; B = 16'h0084; #100;
A = 16'h003; B = 16'h0085; #100;
A = 16'h003; B = 16'h0086; #100;
A = 16'h003; B = 16'h0087; #100;
A = 16'h003; B = 16'h0088; #100;
A = 16'h003; B = 16'h0089; #100;
A = 16'h003; B = 16'h008A; #100;
A = 16'h003; B = 16'h008B; #100;
A = 16'h003; B = 16'h008C; #100;
A = 16'h003; B = 16'h008D; #100;
A = 16'h003; B = 16'h008E; #100;
A = 16'h003; B = 16'h008F; #100;
A = 16'h003; B = 16'h0090; #100;
A = 16'h003; B = 16'h0091; #100;
A = 16'h003; B = 16'h0092; #100;
A = 16'h003; B = 16'h0093; #100;
A = 16'h003; B = 16'h0094; #100;
A = 16'h003; B = 16'h0095; #100;
A = 16'h003; B = 16'h0096; #100;
A = 16'h003; B = 16'h0097; #100;
A = 16'h003; B = 16'h0098; #100;
A = 16'h003; B = 16'h0099; #100;
A = 16'h003; B = 16'h009A; #100;
A = 16'h003; B = 16'h009B; #100;
A = 16'h003; B = 16'h009C; #100;
A = 16'h003; B = 16'h009D; #100;
A = 16'h003; B = 16'h009E; #100;
A = 16'h003; B = 16'h009F; #100;
A = 16'h003; B = 16'h00A0; #100;
A = 16'h003; B = 16'h00A1; #100;
A = 16'h003; B = 16'h00A2; #100;
A = 16'h003; B = 16'h00A3; #100;
A = 16'h003; B = 16'h00A4; #100;
A = 16'h003; B = 16'h00A5; #100;
A = 16'h003; B = 16'h00A6; #100;
A = 16'h003; B = 16'h00A7; #100;
A = 16'h003; B = 16'h00A8; #100;
A = 16'h003; B = 16'h00A9; #100;
A = 16'h003; B = 16'h00AA; #100;
A = 16'h003; B = 16'h00AB; #100;
A = 16'h003; B = 16'h00AC; #100;
A = 16'h003; B = 16'h00AD; #100;
A = 16'h003; B = 16'h00AE; #100;
A = 16'h003; B = 16'h00AF; #100;
A = 16'h003; B = 16'h00B0; #100;
A = 16'h003; B = 16'h00B1; #100;
A = 16'h003; B = 16'h00B2; #100;
A = 16'h003; B = 16'h00B3; #100;
A = 16'h003; B = 16'h00B4; #100;
A = 16'h003; B = 16'h00B5; #100;
A = 16'h003; B = 16'h00B6; #100;
A = 16'h003; B = 16'h00B7; #100;
A = 16'h003; B = 16'h00B8; #100;
A = 16'h003; B = 16'h00B9; #100;
A = 16'h003; B = 16'h00BA; #100;
A = 16'h003; B = 16'h00BB; #100;
A = 16'h003; B = 16'h00BC; #100;
A = 16'h003; B = 16'h00BD; #100;
A = 16'h003; B = 16'h00BE; #100;
A = 16'h003; B = 16'h00BF; #100;
A = 16'h003; B = 16'h00C0; #100;
A = 16'h003; B = 16'h00C1; #100;
A = 16'h003; B = 16'h00C2; #100;
A = 16'h003; B = 16'h00C3; #100;
A = 16'h003; B = 16'h00C4; #100;
A = 16'h003; B = 16'h00C5; #100;
A = 16'h003; B = 16'h00C6; #100;
A = 16'h003; B = 16'h00C7; #100;
A = 16'h003; B = 16'h00C8; #100;
A = 16'h003; B = 16'h00C9; #100;
A = 16'h003; B = 16'h00CA; #100;
A = 16'h003; B = 16'h00CB; #100;
A = 16'h003; B = 16'h00CC; #100;
A = 16'h003; B = 16'h00CD; #100;
A = 16'h003; B = 16'h00CE; #100;
A = 16'h003; B = 16'h00CF; #100;
A = 16'h003; B = 16'h00D0; #100;
A = 16'h003; B = 16'h00D1; #100;
A = 16'h003; B = 16'h00D2; #100;
A = 16'h003; B = 16'h00D3; #100;
A = 16'h003; B = 16'h00D4; #100;
A = 16'h003; B = 16'h00D5; #100;
A = 16'h003; B = 16'h00D6; #100;
A = 16'h003; B = 16'h00D7; #100;
A = 16'h003; B = 16'h00D8; #100;
A = 16'h003; B = 16'h00D9; #100;
A = 16'h003; B = 16'h00DA; #100;
A = 16'h003; B = 16'h00DB; #100;
A = 16'h003; B = 16'h00DC; #100;
A = 16'h003; B = 16'h00DD; #100;
A = 16'h003; B = 16'h00DE; #100;
A = 16'h003; B = 16'h00DF; #100;
A = 16'h003; B = 16'h00E0; #100;
A = 16'h003; B = 16'h00E1; #100;
A = 16'h003; B = 16'h00E2; #100;
A = 16'h003; B = 16'h00E3; #100;
A = 16'h003; B = 16'h00E4; #100;
A = 16'h003; B = 16'h00E5; #100;
A = 16'h003; B = 16'h00E6; #100;
A = 16'h003; B = 16'h00E7; #100;
A = 16'h003; B = 16'h00E8; #100;
A = 16'h003; B = 16'h00E9; #100;
A = 16'h003; B = 16'h00EA; #100;
A = 16'h003; B = 16'h00EB; #100;
A = 16'h003; B = 16'h00EC; #100;
A = 16'h003; B = 16'h00ED; #100;
A = 16'h003; B = 16'h00EE; #100;
A = 16'h003; B = 16'h00EF; #100;
A = 16'h003; B = 16'h00F0; #100;
A = 16'h003; B = 16'h00F1; #100;
A = 16'h003; B = 16'h00F2; #100;
A = 16'h003; B = 16'h00F3; #100;
A = 16'h003; B = 16'h00F4; #100;
A = 16'h003; B = 16'h00F5; #100;
A = 16'h003; B = 16'h00F6; #100;
A = 16'h003; B = 16'h00F7; #100;
A = 16'h003; B = 16'h00F8; #100;
A = 16'h003; B = 16'h00F9; #100;
A = 16'h003; B = 16'h00FA; #100;
A = 16'h003; B = 16'h00FB; #100;
A = 16'h003; B = 16'h00FC; #100;
A = 16'h003; B = 16'h00FD; #100;
A = 16'h003; B = 16'h00FE; #100;
A = 16'h003; B = 16'h00FF; #100;
A = 16'h004; B = 16'h000; #100;
A = 16'h004; B = 16'h001; #100;
A = 16'h004; B = 16'h002; #100;
A = 16'h004; B = 16'h003; #100;
A = 16'h004; B = 16'h004; #100;
A = 16'h004; B = 16'h005; #100;
A = 16'h004; B = 16'h006; #100;
A = 16'h004; B = 16'h007; #100;
A = 16'h004; B = 16'h008; #100;
A = 16'h004; B = 16'h009; #100;
A = 16'h004; B = 16'h00A; #100;
A = 16'h004; B = 16'h00B; #100;
A = 16'h004; B = 16'h00C; #100;
A = 16'h004; B = 16'h00D; #100;
A = 16'h004; B = 16'h00E; #100;
A = 16'h004; B = 16'h00F; #100;
A = 16'h004; B = 16'h0010; #100;
A = 16'h004; B = 16'h0011; #100;
A = 16'h004; B = 16'h0012; #100;
A = 16'h004; B = 16'h0013; #100;
A = 16'h004; B = 16'h0014; #100;
A = 16'h004; B = 16'h0015; #100;
A = 16'h004; B = 16'h0016; #100;
A = 16'h004; B = 16'h0017; #100;
A = 16'h004; B = 16'h0018; #100;
A = 16'h004; B = 16'h0019; #100;
A = 16'h004; B = 16'h001A; #100;
A = 16'h004; B = 16'h001B; #100;
A = 16'h004; B = 16'h001C; #100;
A = 16'h004; B = 16'h001D; #100;
A = 16'h004; B = 16'h001E; #100;
A = 16'h004; B = 16'h001F; #100;
A = 16'h004; B = 16'h0020; #100;
A = 16'h004; B = 16'h0021; #100;
A = 16'h004; B = 16'h0022; #100;
A = 16'h004; B = 16'h0023; #100;
A = 16'h004; B = 16'h0024; #100;
A = 16'h004; B = 16'h0025; #100;
A = 16'h004; B = 16'h0026; #100;
A = 16'h004; B = 16'h0027; #100;
A = 16'h004; B = 16'h0028; #100;
A = 16'h004; B = 16'h0029; #100;
A = 16'h004; B = 16'h002A; #100;
A = 16'h004; B = 16'h002B; #100;
A = 16'h004; B = 16'h002C; #100;
A = 16'h004; B = 16'h002D; #100;
A = 16'h004; B = 16'h002E; #100;
A = 16'h004; B = 16'h002F; #100;
A = 16'h004; B = 16'h0030; #100;
A = 16'h004; B = 16'h0031; #100;
A = 16'h004; B = 16'h0032; #100;
A = 16'h004; B = 16'h0033; #100;
A = 16'h004; B = 16'h0034; #100;
A = 16'h004; B = 16'h0035; #100;
A = 16'h004; B = 16'h0036; #100;
A = 16'h004; B = 16'h0037; #100;
A = 16'h004; B = 16'h0038; #100;
A = 16'h004; B = 16'h0039; #100;
A = 16'h004; B = 16'h003A; #100;
A = 16'h004; B = 16'h003B; #100;
A = 16'h004; B = 16'h003C; #100;
A = 16'h004; B = 16'h003D; #100;
A = 16'h004; B = 16'h003E; #100;
A = 16'h004; B = 16'h003F; #100;
A = 16'h004; B = 16'h0040; #100;
A = 16'h004; B = 16'h0041; #100;
A = 16'h004; B = 16'h0042; #100;
A = 16'h004; B = 16'h0043; #100;
A = 16'h004; B = 16'h0044; #100;
A = 16'h004; B = 16'h0045; #100;
A = 16'h004; B = 16'h0046; #100;
A = 16'h004; B = 16'h0047; #100;
A = 16'h004; B = 16'h0048; #100;
A = 16'h004; B = 16'h0049; #100;
A = 16'h004; B = 16'h004A; #100;
A = 16'h004; B = 16'h004B; #100;
A = 16'h004; B = 16'h004C; #100;
A = 16'h004; B = 16'h004D; #100;
A = 16'h004; B = 16'h004E; #100;
A = 16'h004; B = 16'h004F; #100;
A = 16'h004; B = 16'h0050; #100;
A = 16'h004; B = 16'h0051; #100;
A = 16'h004; B = 16'h0052; #100;
A = 16'h004; B = 16'h0053; #100;
A = 16'h004; B = 16'h0054; #100;
A = 16'h004; B = 16'h0055; #100;
A = 16'h004; B = 16'h0056; #100;
A = 16'h004; B = 16'h0057; #100;
A = 16'h004; B = 16'h0058; #100;
A = 16'h004; B = 16'h0059; #100;
A = 16'h004; B = 16'h005A; #100;
A = 16'h004; B = 16'h005B; #100;
A = 16'h004; B = 16'h005C; #100;
A = 16'h004; B = 16'h005D; #100;
A = 16'h004; B = 16'h005E; #100;
A = 16'h004; B = 16'h005F; #100;
A = 16'h004; B = 16'h0060; #100;
A = 16'h004; B = 16'h0061; #100;
A = 16'h004; B = 16'h0062; #100;
A = 16'h004; B = 16'h0063; #100;
A = 16'h004; B = 16'h0064; #100;
A = 16'h004; B = 16'h0065; #100;
A = 16'h004; B = 16'h0066; #100;
A = 16'h004; B = 16'h0067; #100;
A = 16'h004; B = 16'h0068; #100;
A = 16'h004; B = 16'h0069; #100;
A = 16'h004; B = 16'h006A; #100;
A = 16'h004; B = 16'h006B; #100;
A = 16'h004; B = 16'h006C; #100;
A = 16'h004; B = 16'h006D; #100;
A = 16'h004; B = 16'h006E; #100;
A = 16'h004; B = 16'h006F; #100;
A = 16'h004; B = 16'h0070; #100;
A = 16'h004; B = 16'h0071; #100;
A = 16'h004; B = 16'h0072; #100;
A = 16'h004; B = 16'h0073; #100;
A = 16'h004; B = 16'h0074; #100;
A = 16'h004; B = 16'h0075; #100;
A = 16'h004; B = 16'h0076; #100;
A = 16'h004; B = 16'h0077; #100;
A = 16'h004; B = 16'h0078; #100;
A = 16'h004; B = 16'h0079; #100;
A = 16'h004; B = 16'h007A; #100;
A = 16'h004; B = 16'h007B; #100;
A = 16'h004; B = 16'h007C; #100;
A = 16'h004; B = 16'h007D; #100;
A = 16'h004; B = 16'h007E; #100;
A = 16'h004; B = 16'h007F; #100;
A = 16'h004; B = 16'h0080; #100;
A = 16'h004; B = 16'h0081; #100;
A = 16'h004; B = 16'h0082; #100;
A = 16'h004; B = 16'h0083; #100;
A = 16'h004; B = 16'h0084; #100;
A = 16'h004; B = 16'h0085; #100;
A = 16'h004; B = 16'h0086; #100;
A = 16'h004; B = 16'h0087; #100;
A = 16'h004; B = 16'h0088; #100;
A = 16'h004; B = 16'h0089; #100;
A = 16'h004; B = 16'h008A; #100;
A = 16'h004; B = 16'h008B; #100;
A = 16'h004; B = 16'h008C; #100;
A = 16'h004; B = 16'h008D; #100;
A = 16'h004; B = 16'h008E; #100;
A = 16'h004; B = 16'h008F; #100;
A = 16'h004; B = 16'h0090; #100;
A = 16'h004; B = 16'h0091; #100;
A = 16'h004; B = 16'h0092; #100;
A = 16'h004; B = 16'h0093; #100;
A = 16'h004; B = 16'h0094; #100;
A = 16'h004; B = 16'h0095; #100;
A = 16'h004; B = 16'h0096; #100;
A = 16'h004; B = 16'h0097; #100;
A = 16'h004; B = 16'h0098; #100;
A = 16'h004; B = 16'h0099; #100;
A = 16'h004; B = 16'h009A; #100;
A = 16'h004; B = 16'h009B; #100;
A = 16'h004; B = 16'h009C; #100;
A = 16'h004; B = 16'h009D; #100;
A = 16'h004; B = 16'h009E; #100;
A = 16'h004; B = 16'h009F; #100;
A = 16'h004; B = 16'h00A0; #100;
A = 16'h004; B = 16'h00A1; #100;
A = 16'h004; B = 16'h00A2; #100;
A = 16'h004; B = 16'h00A3; #100;
A = 16'h004; B = 16'h00A4; #100;
A = 16'h004; B = 16'h00A5; #100;
A = 16'h004; B = 16'h00A6; #100;
A = 16'h004; B = 16'h00A7; #100;
A = 16'h004; B = 16'h00A8; #100;
A = 16'h004; B = 16'h00A9; #100;
A = 16'h004; B = 16'h00AA; #100;
A = 16'h004; B = 16'h00AB; #100;
A = 16'h004; B = 16'h00AC; #100;
A = 16'h004; B = 16'h00AD; #100;
A = 16'h004; B = 16'h00AE; #100;
A = 16'h004; B = 16'h00AF; #100;
A = 16'h004; B = 16'h00B0; #100;
A = 16'h004; B = 16'h00B1; #100;
A = 16'h004; B = 16'h00B2; #100;
A = 16'h004; B = 16'h00B3; #100;
A = 16'h004; B = 16'h00B4; #100;
A = 16'h004; B = 16'h00B5; #100;
A = 16'h004; B = 16'h00B6; #100;
A = 16'h004; B = 16'h00B7; #100;
A = 16'h004; B = 16'h00B8; #100;
A = 16'h004; B = 16'h00B9; #100;
A = 16'h004; B = 16'h00BA; #100;
A = 16'h004; B = 16'h00BB; #100;
A = 16'h004; B = 16'h00BC; #100;
A = 16'h004; B = 16'h00BD; #100;
A = 16'h004; B = 16'h00BE; #100;
A = 16'h004; B = 16'h00BF; #100;
A = 16'h004; B = 16'h00C0; #100;
A = 16'h004; B = 16'h00C1; #100;
A = 16'h004; B = 16'h00C2; #100;
A = 16'h004; B = 16'h00C3; #100;
A = 16'h004; B = 16'h00C4; #100;
A = 16'h004; B = 16'h00C5; #100;
A = 16'h004; B = 16'h00C6; #100;
A = 16'h004; B = 16'h00C7; #100;
A = 16'h004; B = 16'h00C8; #100;
A = 16'h004; B = 16'h00C9; #100;
A = 16'h004; B = 16'h00CA; #100;
A = 16'h004; B = 16'h00CB; #100;
A = 16'h004; B = 16'h00CC; #100;
A = 16'h004; B = 16'h00CD; #100;
A = 16'h004; B = 16'h00CE; #100;
A = 16'h004; B = 16'h00CF; #100;
A = 16'h004; B = 16'h00D0; #100;
A = 16'h004; B = 16'h00D1; #100;
A = 16'h004; B = 16'h00D2; #100;
A = 16'h004; B = 16'h00D3; #100;
A = 16'h004; B = 16'h00D4; #100;
A = 16'h004; B = 16'h00D5; #100;
A = 16'h004; B = 16'h00D6; #100;
A = 16'h004; B = 16'h00D7; #100;
A = 16'h004; B = 16'h00D8; #100;
A = 16'h004; B = 16'h00D9; #100;
A = 16'h004; B = 16'h00DA; #100;
A = 16'h004; B = 16'h00DB; #100;
A = 16'h004; B = 16'h00DC; #100;
A = 16'h004; B = 16'h00DD; #100;
A = 16'h004; B = 16'h00DE; #100;
A = 16'h004; B = 16'h00DF; #100;
A = 16'h004; B = 16'h00E0; #100;
A = 16'h004; B = 16'h00E1; #100;
A = 16'h004; B = 16'h00E2; #100;
A = 16'h004; B = 16'h00E3; #100;
A = 16'h004; B = 16'h00E4; #100;
A = 16'h004; B = 16'h00E5; #100;
A = 16'h004; B = 16'h00E6; #100;
A = 16'h004; B = 16'h00E7; #100;
A = 16'h004; B = 16'h00E8; #100;
A = 16'h004; B = 16'h00E9; #100;
A = 16'h004; B = 16'h00EA; #100;
A = 16'h004; B = 16'h00EB; #100;
A = 16'h004; B = 16'h00EC; #100;
A = 16'h004; B = 16'h00ED; #100;
A = 16'h004; B = 16'h00EE; #100;
A = 16'h004; B = 16'h00EF; #100;
A = 16'h004; B = 16'h00F0; #100;
A = 16'h004; B = 16'h00F1; #100;
A = 16'h004; B = 16'h00F2; #100;
A = 16'h004; B = 16'h00F3; #100;
A = 16'h004; B = 16'h00F4; #100;
A = 16'h004; B = 16'h00F5; #100;
A = 16'h004; B = 16'h00F6; #100;
A = 16'h004; B = 16'h00F7; #100;
A = 16'h004; B = 16'h00F8; #100;
A = 16'h004; B = 16'h00F9; #100;
A = 16'h004; B = 16'h00FA; #100;
A = 16'h004; B = 16'h00FB; #100;
A = 16'h004; B = 16'h00FC; #100;
A = 16'h004; B = 16'h00FD; #100;
A = 16'h004; B = 16'h00FE; #100;
A = 16'h004; B = 16'h00FF; #100;
A = 16'h005; B = 16'h000; #100;
A = 16'h005; B = 16'h001; #100;
A = 16'h005; B = 16'h002; #100;
A = 16'h005; B = 16'h003; #100;
A = 16'h005; B = 16'h004; #100;
A = 16'h005; B = 16'h005; #100;
A = 16'h005; B = 16'h006; #100;
A = 16'h005; B = 16'h007; #100;
A = 16'h005; B = 16'h008; #100;
A = 16'h005; B = 16'h009; #100;
A = 16'h005; B = 16'h00A; #100;
A = 16'h005; B = 16'h00B; #100;
A = 16'h005; B = 16'h00C; #100;
A = 16'h005; B = 16'h00D; #100;
A = 16'h005; B = 16'h00E; #100;
A = 16'h005; B = 16'h00F; #100;
A = 16'h005; B = 16'h0010; #100;
A = 16'h005; B = 16'h0011; #100;
A = 16'h005; B = 16'h0012; #100;
A = 16'h005; B = 16'h0013; #100;
A = 16'h005; B = 16'h0014; #100;
A = 16'h005; B = 16'h0015; #100;
A = 16'h005; B = 16'h0016; #100;
A = 16'h005; B = 16'h0017; #100;
A = 16'h005; B = 16'h0018; #100;
A = 16'h005; B = 16'h0019; #100;
A = 16'h005; B = 16'h001A; #100;
A = 16'h005; B = 16'h001B; #100;
A = 16'h005; B = 16'h001C; #100;
A = 16'h005; B = 16'h001D; #100;
A = 16'h005; B = 16'h001E; #100;
A = 16'h005; B = 16'h001F; #100;
A = 16'h005; B = 16'h0020; #100;
A = 16'h005; B = 16'h0021; #100;
A = 16'h005; B = 16'h0022; #100;
A = 16'h005; B = 16'h0023; #100;
A = 16'h005; B = 16'h0024; #100;
A = 16'h005; B = 16'h0025; #100;
A = 16'h005; B = 16'h0026; #100;
A = 16'h005; B = 16'h0027; #100;
A = 16'h005; B = 16'h0028; #100;
A = 16'h005; B = 16'h0029; #100;
A = 16'h005; B = 16'h002A; #100;
A = 16'h005; B = 16'h002B; #100;
A = 16'h005; B = 16'h002C; #100;
A = 16'h005; B = 16'h002D; #100;
A = 16'h005; B = 16'h002E; #100;
A = 16'h005; B = 16'h002F; #100;
A = 16'h005; B = 16'h0030; #100;
A = 16'h005; B = 16'h0031; #100;
A = 16'h005; B = 16'h0032; #100;
A = 16'h005; B = 16'h0033; #100;
A = 16'h005; B = 16'h0034; #100;
A = 16'h005; B = 16'h0035; #100;
A = 16'h005; B = 16'h0036; #100;
A = 16'h005; B = 16'h0037; #100;
A = 16'h005; B = 16'h0038; #100;
A = 16'h005; B = 16'h0039; #100;
A = 16'h005; B = 16'h003A; #100;
A = 16'h005; B = 16'h003B; #100;
A = 16'h005; B = 16'h003C; #100;
A = 16'h005; B = 16'h003D; #100;
A = 16'h005; B = 16'h003E; #100;
A = 16'h005; B = 16'h003F; #100;
A = 16'h005; B = 16'h0040; #100;
A = 16'h005; B = 16'h0041; #100;
A = 16'h005; B = 16'h0042; #100;
A = 16'h005; B = 16'h0043; #100;
A = 16'h005; B = 16'h0044; #100;
A = 16'h005; B = 16'h0045; #100;
A = 16'h005; B = 16'h0046; #100;
A = 16'h005; B = 16'h0047; #100;
A = 16'h005; B = 16'h0048; #100;
A = 16'h005; B = 16'h0049; #100;
A = 16'h005; B = 16'h004A; #100;
A = 16'h005; B = 16'h004B; #100;
A = 16'h005; B = 16'h004C; #100;
A = 16'h005; B = 16'h004D; #100;
A = 16'h005; B = 16'h004E; #100;
A = 16'h005; B = 16'h004F; #100;
A = 16'h005; B = 16'h0050; #100;
A = 16'h005; B = 16'h0051; #100;
A = 16'h005; B = 16'h0052; #100;
A = 16'h005; B = 16'h0053; #100;
A = 16'h005; B = 16'h0054; #100;
A = 16'h005; B = 16'h0055; #100;
A = 16'h005; B = 16'h0056; #100;
A = 16'h005; B = 16'h0057; #100;
A = 16'h005; B = 16'h0058; #100;
A = 16'h005; B = 16'h0059; #100;
A = 16'h005; B = 16'h005A; #100;
A = 16'h005; B = 16'h005B; #100;
A = 16'h005; B = 16'h005C; #100;
A = 16'h005; B = 16'h005D; #100;
A = 16'h005; B = 16'h005E; #100;
A = 16'h005; B = 16'h005F; #100;
A = 16'h005; B = 16'h0060; #100;
A = 16'h005; B = 16'h0061; #100;
A = 16'h005; B = 16'h0062; #100;
A = 16'h005; B = 16'h0063; #100;
A = 16'h005; B = 16'h0064; #100;
A = 16'h005; B = 16'h0065; #100;
A = 16'h005; B = 16'h0066; #100;
A = 16'h005; B = 16'h0067; #100;
A = 16'h005; B = 16'h0068; #100;
A = 16'h005; B = 16'h0069; #100;
A = 16'h005; B = 16'h006A; #100;
A = 16'h005; B = 16'h006B; #100;
A = 16'h005; B = 16'h006C; #100;
A = 16'h005; B = 16'h006D; #100;
A = 16'h005; B = 16'h006E; #100;
A = 16'h005; B = 16'h006F; #100;
A = 16'h005; B = 16'h0070; #100;
A = 16'h005; B = 16'h0071; #100;
A = 16'h005; B = 16'h0072; #100;
A = 16'h005; B = 16'h0073; #100;
A = 16'h005; B = 16'h0074; #100;
A = 16'h005; B = 16'h0075; #100;
A = 16'h005; B = 16'h0076; #100;
A = 16'h005; B = 16'h0077; #100;
A = 16'h005; B = 16'h0078; #100;
A = 16'h005; B = 16'h0079; #100;
A = 16'h005; B = 16'h007A; #100;
A = 16'h005; B = 16'h007B; #100;
A = 16'h005; B = 16'h007C; #100;
A = 16'h005; B = 16'h007D; #100;
A = 16'h005; B = 16'h007E; #100;
A = 16'h005; B = 16'h007F; #100;
A = 16'h005; B = 16'h0080; #100;
A = 16'h005; B = 16'h0081; #100;
A = 16'h005; B = 16'h0082; #100;
A = 16'h005; B = 16'h0083; #100;
A = 16'h005; B = 16'h0084; #100;
A = 16'h005; B = 16'h0085; #100;
A = 16'h005; B = 16'h0086; #100;
A = 16'h005; B = 16'h0087; #100;
A = 16'h005; B = 16'h0088; #100;
A = 16'h005; B = 16'h0089; #100;
A = 16'h005; B = 16'h008A; #100;
A = 16'h005; B = 16'h008B; #100;
A = 16'h005; B = 16'h008C; #100;
A = 16'h005; B = 16'h008D; #100;
A = 16'h005; B = 16'h008E; #100;
A = 16'h005; B = 16'h008F; #100;
A = 16'h005; B = 16'h0090; #100;
A = 16'h005; B = 16'h0091; #100;
A = 16'h005; B = 16'h0092; #100;
A = 16'h005; B = 16'h0093; #100;
A = 16'h005; B = 16'h0094; #100;
A = 16'h005; B = 16'h0095; #100;
A = 16'h005; B = 16'h0096; #100;
A = 16'h005; B = 16'h0097; #100;
A = 16'h005; B = 16'h0098; #100;
A = 16'h005; B = 16'h0099; #100;
A = 16'h005; B = 16'h009A; #100;
A = 16'h005; B = 16'h009B; #100;
A = 16'h005; B = 16'h009C; #100;
A = 16'h005; B = 16'h009D; #100;
A = 16'h005; B = 16'h009E; #100;
A = 16'h005; B = 16'h009F; #100;
A = 16'h005; B = 16'h00A0; #100;
A = 16'h005; B = 16'h00A1; #100;
A = 16'h005; B = 16'h00A2; #100;
A = 16'h005; B = 16'h00A3; #100;
A = 16'h005; B = 16'h00A4; #100;
A = 16'h005; B = 16'h00A5; #100;
A = 16'h005; B = 16'h00A6; #100;
A = 16'h005; B = 16'h00A7; #100;
A = 16'h005; B = 16'h00A8; #100;
A = 16'h005; B = 16'h00A9; #100;
A = 16'h005; B = 16'h00AA; #100;
A = 16'h005; B = 16'h00AB; #100;
A = 16'h005; B = 16'h00AC; #100;
A = 16'h005; B = 16'h00AD; #100;
A = 16'h005; B = 16'h00AE; #100;
A = 16'h005; B = 16'h00AF; #100;
A = 16'h005; B = 16'h00B0; #100;
A = 16'h005; B = 16'h00B1; #100;
A = 16'h005; B = 16'h00B2; #100;
A = 16'h005; B = 16'h00B3; #100;
A = 16'h005; B = 16'h00B4; #100;
A = 16'h005; B = 16'h00B5; #100;
A = 16'h005; B = 16'h00B6; #100;
A = 16'h005; B = 16'h00B7; #100;
A = 16'h005; B = 16'h00B8; #100;
A = 16'h005; B = 16'h00B9; #100;
A = 16'h005; B = 16'h00BA; #100;
A = 16'h005; B = 16'h00BB; #100;
A = 16'h005; B = 16'h00BC; #100;
A = 16'h005; B = 16'h00BD; #100;
A = 16'h005; B = 16'h00BE; #100;
A = 16'h005; B = 16'h00BF; #100;
A = 16'h005; B = 16'h00C0; #100;
A = 16'h005; B = 16'h00C1; #100;
A = 16'h005; B = 16'h00C2; #100;
A = 16'h005; B = 16'h00C3; #100;
A = 16'h005; B = 16'h00C4; #100;
A = 16'h005; B = 16'h00C5; #100;
A = 16'h005; B = 16'h00C6; #100;
A = 16'h005; B = 16'h00C7; #100;
A = 16'h005; B = 16'h00C8; #100;
A = 16'h005; B = 16'h00C9; #100;
A = 16'h005; B = 16'h00CA; #100;
A = 16'h005; B = 16'h00CB; #100;
A = 16'h005; B = 16'h00CC; #100;
A = 16'h005; B = 16'h00CD; #100;
A = 16'h005; B = 16'h00CE; #100;
A = 16'h005; B = 16'h00CF; #100;
A = 16'h005; B = 16'h00D0; #100;
A = 16'h005; B = 16'h00D1; #100;
A = 16'h005; B = 16'h00D2; #100;
A = 16'h005; B = 16'h00D3; #100;
A = 16'h005; B = 16'h00D4; #100;
A = 16'h005; B = 16'h00D5; #100;
A = 16'h005; B = 16'h00D6; #100;
A = 16'h005; B = 16'h00D7; #100;
A = 16'h005; B = 16'h00D8; #100;
A = 16'h005; B = 16'h00D9; #100;
A = 16'h005; B = 16'h00DA; #100;
A = 16'h005; B = 16'h00DB; #100;
A = 16'h005; B = 16'h00DC; #100;
A = 16'h005; B = 16'h00DD; #100;
A = 16'h005; B = 16'h00DE; #100;
A = 16'h005; B = 16'h00DF; #100;
A = 16'h005; B = 16'h00E0; #100;
A = 16'h005; B = 16'h00E1; #100;
A = 16'h005; B = 16'h00E2; #100;
A = 16'h005; B = 16'h00E3; #100;
A = 16'h005; B = 16'h00E4; #100;
A = 16'h005; B = 16'h00E5; #100;
A = 16'h005; B = 16'h00E6; #100;
A = 16'h005; B = 16'h00E7; #100;
A = 16'h005; B = 16'h00E8; #100;
A = 16'h005; B = 16'h00E9; #100;
A = 16'h005; B = 16'h00EA; #100;
A = 16'h005; B = 16'h00EB; #100;
A = 16'h005; B = 16'h00EC; #100;
A = 16'h005; B = 16'h00ED; #100;
A = 16'h005; B = 16'h00EE; #100;
A = 16'h005; B = 16'h00EF; #100;
A = 16'h005; B = 16'h00F0; #100;
A = 16'h005; B = 16'h00F1; #100;
A = 16'h005; B = 16'h00F2; #100;
A = 16'h005; B = 16'h00F3; #100;
A = 16'h005; B = 16'h00F4; #100;
A = 16'h005; B = 16'h00F5; #100;
A = 16'h005; B = 16'h00F6; #100;
A = 16'h005; B = 16'h00F7; #100;
A = 16'h005; B = 16'h00F8; #100;
A = 16'h005; B = 16'h00F9; #100;
A = 16'h005; B = 16'h00FA; #100;
A = 16'h005; B = 16'h00FB; #100;
A = 16'h005; B = 16'h00FC; #100;
A = 16'h005; B = 16'h00FD; #100;
A = 16'h005; B = 16'h00FE; #100;
A = 16'h005; B = 16'h00FF; #100;
A = 16'h006; B = 16'h000; #100;
A = 16'h006; B = 16'h001; #100;
A = 16'h006; B = 16'h002; #100;
A = 16'h006; B = 16'h003; #100;
A = 16'h006; B = 16'h004; #100;
A = 16'h006; B = 16'h005; #100;
A = 16'h006; B = 16'h006; #100;
A = 16'h006; B = 16'h007; #100;
A = 16'h006; B = 16'h008; #100;
A = 16'h006; B = 16'h009; #100;
A = 16'h006; B = 16'h00A; #100;
A = 16'h006; B = 16'h00B; #100;
A = 16'h006; B = 16'h00C; #100;
A = 16'h006; B = 16'h00D; #100;
A = 16'h006; B = 16'h00E; #100;
A = 16'h006; B = 16'h00F; #100;
A = 16'h006; B = 16'h0010; #100;
A = 16'h006; B = 16'h0011; #100;
A = 16'h006; B = 16'h0012; #100;
A = 16'h006; B = 16'h0013; #100;
A = 16'h006; B = 16'h0014; #100;
A = 16'h006; B = 16'h0015; #100;
A = 16'h006; B = 16'h0016; #100;
A = 16'h006; B = 16'h0017; #100;
A = 16'h006; B = 16'h0018; #100;
A = 16'h006; B = 16'h0019; #100;
A = 16'h006; B = 16'h001A; #100;
A = 16'h006; B = 16'h001B; #100;
A = 16'h006; B = 16'h001C; #100;
A = 16'h006; B = 16'h001D; #100;
A = 16'h006; B = 16'h001E; #100;
A = 16'h006; B = 16'h001F; #100;
A = 16'h006; B = 16'h0020; #100;
A = 16'h006; B = 16'h0021; #100;
A = 16'h006; B = 16'h0022; #100;
A = 16'h006; B = 16'h0023; #100;
A = 16'h006; B = 16'h0024; #100;
A = 16'h006; B = 16'h0025; #100;
A = 16'h006; B = 16'h0026; #100;
A = 16'h006; B = 16'h0027; #100;
A = 16'h006; B = 16'h0028; #100;
A = 16'h006; B = 16'h0029; #100;
A = 16'h006; B = 16'h002A; #100;
A = 16'h006; B = 16'h002B; #100;
A = 16'h006; B = 16'h002C; #100;
A = 16'h006; B = 16'h002D; #100;
A = 16'h006; B = 16'h002E; #100;
A = 16'h006; B = 16'h002F; #100;
A = 16'h006; B = 16'h0030; #100;
A = 16'h006; B = 16'h0031; #100;
A = 16'h006; B = 16'h0032; #100;
A = 16'h006; B = 16'h0033; #100;
A = 16'h006; B = 16'h0034; #100;
A = 16'h006; B = 16'h0035; #100;
A = 16'h006; B = 16'h0036; #100;
A = 16'h006; B = 16'h0037; #100;
A = 16'h006; B = 16'h0038; #100;
A = 16'h006; B = 16'h0039; #100;
A = 16'h006; B = 16'h003A; #100;
A = 16'h006; B = 16'h003B; #100;
A = 16'h006; B = 16'h003C; #100;
A = 16'h006; B = 16'h003D; #100;
A = 16'h006; B = 16'h003E; #100;
A = 16'h006; B = 16'h003F; #100;
A = 16'h006; B = 16'h0040; #100;
A = 16'h006; B = 16'h0041; #100;
A = 16'h006; B = 16'h0042; #100;
A = 16'h006; B = 16'h0043; #100;
A = 16'h006; B = 16'h0044; #100;
A = 16'h006; B = 16'h0045; #100;
A = 16'h006; B = 16'h0046; #100;
A = 16'h006; B = 16'h0047; #100;
A = 16'h006; B = 16'h0048; #100;
A = 16'h006; B = 16'h0049; #100;
A = 16'h006; B = 16'h004A; #100;
A = 16'h006; B = 16'h004B; #100;
A = 16'h006; B = 16'h004C; #100;
A = 16'h006; B = 16'h004D; #100;
A = 16'h006; B = 16'h004E; #100;
A = 16'h006; B = 16'h004F; #100;
A = 16'h006; B = 16'h0050; #100;
A = 16'h006; B = 16'h0051; #100;
A = 16'h006; B = 16'h0052; #100;
A = 16'h006; B = 16'h0053; #100;
A = 16'h006; B = 16'h0054; #100;
A = 16'h006; B = 16'h0055; #100;
A = 16'h006; B = 16'h0056; #100;
A = 16'h006; B = 16'h0057; #100;
A = 16'h006; B = 16'h0058; #100;
A = 16'h006; B = 16'h0059; #100;
A = 16'h006; B = 16'h005A; #100;
A = 16'h006; B = 16'h005B; #100;
A = 16'h006; B = 16'h005C; #100;
A = 16'h006; B = 16'h005D; #100;
A = 16'h006; B = 16'h005E; #100;
A = 16'h006; B = 16'h005F; #100;
A = 16'h006; B = 16'h0060; #100;
A = 16'h006; B = 16'h0061; #100;
A = 16'h006; B = 16'h0062; #100;
A = 16'h006; B = 16'h0063; #100;
A = 16'h006; B = 16'h0064; #100;
A = 16'h006; B = 16'h0065; #100;
A = 16'h006; B = 16'h0066; #100;
A = 16'h006; B = 16'h0067; #100;
A = 16'h006; B = 16'h0068; #100;
A = 16'h006; B = 16'h0069; #100;
A = 16'h006; B = 16'h006A; #100;
A = 16'h006; B = 16'h006B; #100;
A = 16'h006; B = 16'h006C; #100;
A = 16'h006; B = 16'h006D; #100;
A = 16'h006; B = 16'h006E; #100;
A = 16'h006; B = 16'h006F; #100;
A = 16'h006; B = 16'h0070; #100;
A = 16'h006; B = 16'h0071; #100;
A = 16'h006; B = 16'h0072; #100;
A = 16'h006; B = 16'h0073; #100;
A = 16'h006; B = 16'h0074; #100;
A = 16'h006; B = 16'h0075; #100;
A = 16'h006; B = 16'h0076; #100;
A = 16'h006; B = 16'h0077; #100;
A = 16'h006; B = 16'h0078; #100;
A = 16'h006; B = 16'h0079; #100;
A = 16'h006; B = 16'h007A; #100;
A = 16'h006; B = 16'h007B; #100;
A = 16'h006; B = 16'h007C; #100;
A = 16'h006; B = 16'h007D; #100;
A = 16'h006; B = 16'h007E; #100;
A = 16'h006; B = 16'h007F; #100;
A = 16'h006; B = 16'h0080; #100;
A = 16'h006; B = 16'h0081; #100;
A = 16'h006; B = 16'h0082; #100;
A = 16'h006; B = 16'h0083; #100;
A = 16'h006; B = 16'h0084; #100;
A = 16'h006; B = 16'h0085; #100;
A = 16'h006; B = 16'h0086; #100;
A = 16'h006; B = 16'h0087; #100;
A = 16'h006; B = 16'h0088; #100;
A = 16'h006; B = 16'h0089; #100;
A = 16'h006; B = 16'h008A; #100;
A = 16'h006; B = 16'h008B; #100;
A = 16'h006; B = 16'h008C; #100;
A = 16'h006; B = 16'h008D; #100;
A = 16'h006; B = 16'h008E; #100;
A = 16'h006; B = 16'h008F; #100;
A = 16'h006; B = 16'h0090; #100;
A = 16'h006; B = 16'h0091; #100;
A = 16'h006; B = 16'h0092; #100;
A = 16'h006; B = 16'h0093; #100;
A = 16'h006; B = 16'h0094; #100;
A = 16'h006; B = 16'h0095; #100;
A = 16'h006; B = 16'h0096; #100;
A = 16'h006; B = 16'h0097; #100;
A = 16'h006; B = 16'h0098; #100;
A = 16'h006; B = 16'h0099; #100;
A = 16'h006; B = 16'h009A; #100;
A = 16'h006; B = 16'h009B; #100;
A = 16'h006; B = 16'h009C; #100;
A = 16'h006; B = 16'h009D; #100;
A = 16'h006; B = 16'h009E; #100;
A = 16'h006; B = 16'h009F; #100;
A = 16'h006; B = 16'h00A0; #100;
A = 16'h006; B = 16'h00A1; #100;
A = 16'h006; B = 16'h00A2; #100;
A = 16'h006; B = 16'h00A3; #100;
A = 16'h006; B = 16'h00A4; #100;
A = 16'h006; B = 16'h00A5; #100;
A = 16'h006; B = 16'h00A6; #100;
A = 16'h006; B = 16'h00A7; #100;
A = 16'h006; B = 16'h00A8; #100;
A = 16'h006; B = 16'h00A9; #100;
A = 16'h006; B = 16'h00AA; #100;
A = 16'h006; B = 16'h00AB; #100;
A = 16'h006; B = 16'h00AC; #100;
A = 16'h006; B = 16'h00AD; #100;
A = 16'h006; B = 16'h00AE; #100;
A = 16'h006; B = 16'h00AF; #100;
A = 16'h006; B = 16'h00B0; #100;
A = 16'h006; B = 16'h00B1; #100;
A = 16'h006; B = 16'h00B2; #100;
A = 16'h006; B = 16'h00B3; #100;
A = 16'h006; B = 16'h00B4; #100;
A = 16'h006; B = 16'h00B5; #100;
A = 16'h006; B = 16'h00B6; #100;
A = 16'h006; B = 16'h00B7; #100;
A = 16'h006; B = 16'h00B8; #100;
A = 16'h006; B = 16'h00B9; #100;
A = 16'h006; B = 16'h00BA; #100;
A = 16'h006; B = 16'h00BB; #100;
A = 16'h006; B = 16'h00BC; #100;
A = 16'h006; B = 16'h00BD; #100;
A = 16'h006; B = 16'h00BE; #100;
A = 16'h006; B = 16'h00BF; #100;
A = 16'h006; B = 16'h00C0; #100;
A = 16'h006; B = 16'h00C1; #100;
A = 16'h006; B = 16'h00C2; #100;
A = 16'h006; B = 16'h00C3; #100;
A = 16'h006; B = 16'h00C4; #100;
A = 16'h006; B = 16'h00C5; #100;
A = 16'h006; B = 16'h00C6; #100;
A = 16'h006; B = 16'h00C7; #100;
A = 16'h006; B = 16'h00C8; #100;
A = 16'h006; B = 16'h00C9; #100;
A = 16'h006; B = 16'h00CA; #100;
A = 16'h006; B = 16'h00CB; #100;
A = 16'h006; B = 16'h00CC; #100;
A = 16'h006; B = 16'h00CD; #100;
A = 16'h006; B = 16'h00CE; #100;
A = 16'h006; B = 16'h00CF; #100;
A = 16'h006; B = 16'h00D0; #100;
A = 16'h006; B = 16'h00D1; #100;
A = 16'h006; B = 16'h00D2; #100;
A = 16'h006; B = 16'h00D3; #100;
A = 16'h006; B = 16'h00D4; #100;
A = 16'h006; B = 16'h00D5; #100;
A = 16'h006; B = 16'h00D6; #100;
A = 16'h006; B = 16'h00D7; #100;
A = 16'h006; B = 16'h00D8; #100;
A = 16'h006; B = 16'h00D9; #100;
A = 16'h006; B = 16'h00DA; #100;
A = 16'h006; B = 16'h00DB; #100;
A = 16'h006; B = 16'h00DC; #100;
A = 16'h006; B = 16'h00DD; #100;
A = 16'h006; B = 16'h00DE; #100;
A = 16'h006; B = 16'h00DF; #100;
A = 16'h006; B = 16'h00E0; #100;
A = 16'h006; B = 16'h00E1; #100;
A = 16'h006; B = 16'h00E2; #100;
A = 16'h006; B = 16'h00E3; #100;
A = 16'h006; B = 16'h00E4; #100;
A = 16'h006; B = 16'h00E5; #100;
A = 16'h006; B = 16'h00E6; #100;
A = 16'h006; B = 16'h00E7; #100;
A = 16'h006; B = 16'h00E8; #100;
A = 16'h006; B = 16'h00E9; #100;
A = 16'h006; B = 16'h00EA; #100;
A = 16'h006; B = 16'h00EB; #100;
A = 16'h006; B = 16'h00EC; #100;
A = 16'h006; B = 16'h00ED; #100;
A = 16'h006; B = 16'h00EE; #100;
A = 16'h006; B = 16'h00EF; #100;
A = 16'h006; B = 16'h00F0; #100;
A = 16'h006; B = 16'h00F1; #100;
A = 16'h006; B = 16'h00F2; #100;
A = 16'h006; B = 16'h00F3; #100;
A = 16'h006; B = 16'h00F4; #100;
A = 16'h006; B = 16'h00F5; #100;
A = 16'h006; B = 16'h00F6; #100;
A = 16'h006; B = 16'h00F7; #100;
A = 16'h006; B = 16'h00F8; #100;
A = 16'h006; B = 16'h00F9; #100;
A = 16'h006; B = 16'h00FA; #100;
A = 16'h006; B = 16'h00FB; #100;
A = 16'h006; B = 16'h00FC; #100;
A = 16'h006; B = 16'h00FD; #100;
A = 16'h006; B = 16'h00FE; #100;
A = 16'h006; B = 16'h00FF; #100;
A = 16'h007; B = 16'h000; #100;
A = 16'h007; B = 16'h001; #100;
A = 16'h007; B = 16'h002; #100;
A = 16'h007; B = 16'h003; #100;
A = 16'h007; B = 16'h004; #100;
A = 16'h007; B = 16'h005; #100;
A = 16'h007; B = 16'h006; #100;
A = 16'h007; B = 16'h007; #100;
A = 16'h007; B = 16'h008; #100;
A = 16'h007; B = 16'h009; #100;
A = 16'h007; B = 16'h00A; #100;
A = 16'h007; B = 16'h00B; #100;
A = 16'h007; B = 16'h00C; #100;
A = 16'h007; B = 16'h00D; #100;
A = 16'h007; B = 16'h00E; #100;
A = 16'h007; B = 16'h00F; #100;
A = 16'h007; B = 16'h0010; #100;
A = 16'h007; B = 16'h0011; #100;
A = 16'h007; B = 16'h0012; #100;
A = 16'h007; B = 16'h0013; #100;
A = 16'h007; B = 16'h0014; #100;
A = 16'h007; B = 16'h0015; #100;
A = 16'h007; B = 16'h0016; #100;
A = 16'h007; B = 16'h0017; #100;
A = 16'h007; B = 16'h0018; #100;
A = 16'h007; B = 16'h0019; #100;
A = 16'h007; B = 16'h001A; #100;
A = 16'h007; B = 16'h001B; #100;
A = 16'h007; B = 16'h001C; #100;
A = 16'h007; B = 16'h001D; #100;
A = 16'h007; B = 16'h001E; #100;
A = 16'h007; B = 16'h001F; #100;
A = 16'h007; B = 16'h0020; #100;
A = 16'h007; B = 16'h0021; #100;
A = 16'h007; B = 16'h0022; #100;
A = 16'h007; B = 16'h0023; #100;
A = 16'h007; B = 16'h0024; #100;
A = 16'h007; B = 16'h0025; #100;
A = 16'h007; B = 16'h0026; #100;
A = 16'h007; B = 16'h0027; #100;
A = 16'h007; B = 16'h0028; #100;
A = 16'h007; B = 16'h0029; #100;
A = 16'h007; B = 16'h002A; #100;
A = 16'h007; B = 16'h002B; #100;
A = 16'h007; B = 16'h002C; #100;
A = 16'h007; B = 16'h002D; #100;
A = 16'h007; B = 16'h002E; #100;
A = 16'h007; B = 16'h002F; #100;
A = 16'h007; B = 16'h0030; #100;
A = 16'h007; B = 16'h0031; #100;
A = 16'h007; B = 16'h0032; #100;
A = 16'h007; B = 16'h0033; #100;
A = 16'h007; B = 16'h0034; #100;
A = 16'h007; B = 16'h0035; #100;
A = 16'h007; B = 16'h0036; #100;
A = 16'h007; B = 16'h0037; #100;
A = 16'h007; B = 16'h0038; #100;
A = 16'h007; B = 16'h0039; #100;
A = 16'h007; B = 16'h003A; #100;
A = 16'h007; B = 16'h003B; #100;
A = 16'h007; B = 16'h003C; #100;
A = 16'h007; B = 16'h003D; #100;
A = 16'h007; B = 16'h003E; #100;
A = 16'h007; B = 16'h003F; #100;
A = 16'h007; B = 16'h0040; #100;
A = 16'h007; B = 16'h0041; #100;
A = 16'h007; B = 16'h0042; #100;
A = 16'h007; B = 16'h0043; #100;
A = 16'h007; B = 16'h0044; #100;
A = 16'h007; B = 16'h0045; #100;
A = 16'h007; B = 16'h0046; #100;
A = 16'h007; B = 16'h0047; #100;
A = 16'h007; B = 16'h0048; #100;
A = 16'h007; B = 16'h0049; #100;
A = 16'h007; B = 16'h004A; #100;
A = 16'h007; B = 16'h004B; #100;
A = 16'h007; B = 16'h004C; #100;
A = 16'h007; B = 16'h004D; #100;
A = 16'h007; B = 16'h004E; #100;
A = 16'h007; B = 16'h004F; #100;
A = 16'h007; B = 16'h0050; #100;
A = 16'h007; B = 16'h0051; #100;
A = 16'h007; B = 16'h0052; #100;
A = 16'h007; B = 16'h0053; #100;
A = 16'h007; B = 16'h0054; #100;
A = 16'h007; B = 16'h0055; #100;
A = 16'h007; B = 16'h0056; #100;
A = 16'h007; B = 16'h0057; #100;
A = 16'h007; B = 16'h0058; #100;
A = 16'h007; B = 16'h0059; #100;
A = 16'h007; B = 16'h005A; #100;
A = 16'h007; B = 16'h005B; #100;
A = 16'h007; B = 16'h005C; #100;
A = 16'h007; B = 16'h005D; #100;
A = 16'h007; B = 16'h005E; #100;
A = 16'h007; B = 16'h005F; #100;
A = 16'h007; B = 16'h0060; #100;
A = 16'h007; B = 16'h0061; #100;
A = 16'h007; B = 16'h0062; #100;
A = 16'h007; B = 16'h0063; #100;
A = 16'h007; B = 16'h0064; #100;
A = 16'h007; B = 16'h0065; #100;
A = 16'h007; B = 16'h0066; #100;
A = 16'h007; B = 16'h0067; #100;
A = 16'h007; B = 16'h0068; #100;
A = 16'h007; B = 16'h0069; #100;
A = 16'h007; B = 16'h006A; #100;
A = 16'h007; B = 16'h006B; #100;
A = 16'h007; B = 16'h006C; #100;
A = 16'h007; B = 16'h006D; #100;
A = 16'h007; B = 16'h006E; #100;
A = 16'h007; B = 16'h006F; #100;
A = 16'h007; B = 16'h0070; #100;
A = 16'h007; B = 16'h0071; #100;
A = 16'h007; B = 16'h0072; #100;
A = 16'h007; B = 16'h0073; #100;
A = 16'h007; B = 16'h0074; #100;
A = 16'h007; B = 16'h0075; #100;
A = 16'h007; B = 16'h0076; #100;
A = 16'h007; B = 16'h0077; #100;
A = 16'h007; B = 16'h0078; #100;
A = 16'h007; B = 16'h0079; #100;
A = 16'h007; B = 16'h007A; #100;
A = 16'h007; B = 16'h007B; #100;
A = 16'h007; B = 16'h007C; #100;
A = 16'h007; B = 16'h007D; #100;
A = 16'h007; B = 16'h007E; #100;
A = 16'h007; B = 16'h007F; #100;
A = 16'h007; B = 16'h0080; #100;
A = 16'h007; B = 16'h0081; #100;
A = 16'h007; B = 16'h0082; #100;
A = 16'h007; B = 16'h0083; #100;
A = 16'h007; B = 16'h0084; #100;
A = 16'h007; B = 16'h0085; #100;
A = 16'h007; B = 16'h0086; #100;
A = 16'h007; B = 16'h0087; #100;
A = 16'h007; B = 16'h0088; #100;
A = 16'h007; B = 16'h0089; #100;
A = 16'h007; B = 16'h008A; #100;
A = 16'h007; B = 16'h008B; #100;
A = 16'h007; B = 16'h008C; #100;
A = 16'h007; B = 16'h008D; #100;
A = 16'h007; B = 16'h008E; #100;
A = 16'h007; B = 16'h008F; #100;
A = 16'h007; B = 16'h0090; #100;
A = 16'h007; B = 16'h0091; #100;
A = 16'h007; B = 16'h0092; #100;
A = 16'h007; B = 16'h0093; #100;
A = 16'h007; B = 16'h0094; #100;
A = 16'h007; B = 16'h0095; #100;
A = 16'h007; B = 16'h0096; #100;
A = 16'h007; B = 16'h0097; #100;
A = 16'h007; B = 16'h0098; #100;
A = 16'h007; B = 16'h0099; #100;
A = 16'h007; B = 16'h009A; #100;
A = 16'h007; B = 16'h009B; #100;
A = 16'h007; B = 16'h009C; #100;
A = 16'h007; B = 16'h009D; #100;
A = 16'h007; B = 16'h009E; #100;
A = 16'h007; B = 16'h009F; #100;
A = 16'h007; B = 16'h00A0; #100;
A = 16'h007; B = 16'h00A1; #100;
A = 16'h007; B = 16'h00A2; #100;
A = 16'h007; B = 16'h00A3; #100;
A = 16'h007; B = 16'h00A4; #100;
A = 16'h007; B = 16'h00A5; #100;
A = 16'h007; B = 16'h00A6; #100;
A = 16'h007; B = 16'h00A7; #100;
A = 16'h007; B = 16'h00A8; #100;
A = 16'h007; B = 16'h00A9; #100;
A = 16'h007; B = 16'h00AA; #100;
A = 16'h007; B = 16'h00AB; #100;
A = 16'h007; B = 16'h00AC; #100;
A = 16'h007; B = 16'h00AD; #100;
A = 16'h007; B = 16'h00AE; #100;
A = 16'h007; B = 16'h00AF; #100;
A = 16'h007; B = 16'h00B0; #100;
A = 16'h007; B = 16'h00B1; #100;
A = 16'h007; B = 16'h00B2; #100;
A = 16'h007; B = 16'h00B3; #100;
A = 16'h007; B = 16'h00B4; #100;
A = 16'h007; B = 16'h00B5; #100;
A = 16'h007; B = 16'h00B6; #100;
A = 16'h007; B = 16'h00B7; #100;
A = 16'h007; B = 16'h00B8; #100;
A = 16'h007; B = 16'h00B9; #100;
A = 16'h007; B = 16'h00BA; #100;
A = 16'h007; B = 16'h00BB; #100;
A = 16'h007; B = 16'h00BC; #100;
A = 16'h007; B = 16'h00BD; #100;
A = 16'h007; B = 16'h00BE; #100;
A = 16'h007; B = 16'h00BF; #100;
A = 16'h007; B = 16'h00C0; #100;
A = 16'h007; B = 16'h00C1; #100;
A = 16'h007; B = 16'h00C2; #100;
A = 16'h007; B = 16'h00C3; #100;
A = 16'h007; B = 16'h00C4; #100;
A = 16'h007; B = 16'h00C5; #100;
A = 16'h007; B = 16'h00C6; #100;
A = 16'h007; B = 16'h00C7; #100;
A = 16'h007; B = 16'h00C8; #100;
A = 16'h007; B = 16'h00C9; #100;
A = 16'h007; B = 16'h00CA; #100;
A = 16'h007; B = 16'h00CB; #100;
A = 16'h007; B = 16'h00CC; #100;
A = 16'h007; B = 16'h00CD; #100;
A = 16'h007; B = 16'h00CE; #100;
A = 16'h007; B = 16'h00CF; #100;
A = 16'h007; B = 16'h00D0; #100;
A = 16'h007; B = 16'h00D1; #100;
A = 16'h007; B = 16'h00D2; #100;
A = 16'h007; B = 16'h00D3; #100;
A = 16'h007; B = 16'h00D4; #100;
A = 16'h007; B = 16'h00D5; #100;
A = 16'h007; B = 16'h00D6; #100;
A = 16'h007; B = 16'h00D7; #100;
A = 16'h007; B = 16'h00D8; #100;
A = 16'h007; B = 16'h00D9; #100;
A = 16'h007; B = 16'h00DA; #100;
A = 16'h007; B = 16'h00DB; #100;
A = 16'h007; B = 16'h00DC; #100;
A = 16'h007; B = 16'h00DD; #100;
A = 16'h007; B = 16'h00DE; #100;
A = 16'h007; B = 16'h00DF; #100;
A = 16'h007; B = 16'h00E0; #100;
A = 16'h007; B = 16'h00E1; #100;
A = 16'h007; B = 16'h00E2; #100;
A = 16'h007; B = 16'h00E3; #100;
A = 16'h007; B = 16'h00E4; #100;
A = 16'h007; B = 16'h00E5; #100;
A = 16'h007; B = 16'h00E6; #100;
A = 16'h007; B = 16'h00E7; #100;
A = 16'h007; B = 16'h00E8; #100;
A = 16'h007; B = 16'h00E9; #100;
A = 16'h007; B = 16'h00EA; #100;
A = 16'h007; B = 16'h00EB; #100;
A = 16'h007; B = 16'h00EC; #100;
A = 16'h007; B = 16'h00ED; #100;
A = 16'h007; B = 16'h00EE; #100;
A = 16'h007; B = 16'h00EF; #100;
A = 16'h007; B = 16'h00F0; #100;
A = 16'h007; B = 16'h00F1; #100;
A = 16'h007; B = 16'h00F2; #100;
A = 16'h007; B = 16'h00F3; #100;
A = 16'h007; B = 16'h00F4; #100;
A = 16'h007; B = 16'h00F5; #100;
A = 16'h007; B = 16'h00F6; #100;
A = 16'h007; B = 16'h00F7; #100;
A = 16'h007; B = 16'h00F8; #100;
A = 16'h007; B = 16'h00F9; #100;
A = 16'h007; B = 16'h00FA; #100;
A = 16'h007; B = 16'h00FB; #100;
A = 16'h007; B = 16'h00FC; #100;
A = 16'h007; B = 16'h00FD; #100;
A = 16'h007; B = 16'h00FE; #100;
A = 16'h007; B = 16'h00FF; #100;
A = 16'h008; B = 16'h000; #100;
A = 16'h008; B = 16'h001; #100;
A = 16'h008; B = 16'h002; #100;
A = 16'h008; B = 16'h003; #100;
A = 16'h008; B = 16'h004; #100;
A = 16'h008; B = 16'h005; #100;
A = 16'h008; B = 16'h006; #100;
A = 16'h008; B = 16'h007; #100;
A = 16'h008; B = 16'h008; #100;
A = 16'h008; B = 16'h009; #100;
A = 16'h008; B = 16'h00A; #100;
A = 16'h008; B = 16'h00B; #100;
A = 16'h008; B = 16'h00C; #100;
A = 16'h008; B = 16'h00D; #100;
A = 16'h008; B = 16'h00E; #100;
A = 16'h008; B = 16'h00F; #100;
A = 16'h008; B = 16'h0010; #100;
A = 16'h008; B = 16'h0011; #100;
A = 16'h008; B = 16'h0012; #100;
A = 16'h008; B = 16'h0013; #100;
A = 16'h008; B = 16'h0014; #100;
A = 16'h008; B = 16'h0015; #100;
A = 16'h008; B = 16'h0016; #100;
A = 16'h008; B = 16'h0017; #100;
A = 16'h008; B = 16'h0018; #100;
A = 16'h008; B = 16'h0019; #100;
A = 16'h008; B = 16'h001A; #100;
A = 16'h008; B = 16'h001B; #100;
A = 16'h008; B = 16'h001C; #100;
A = 16'h008; B = 16'h001D; #100;
A = 16'h008; B = 16'h001E; #100;
A = 16'h008; B = 16'h001F; #100;
A = 16'h008; B = 16'h0020; #100;
A = 16'h008; B = 16'h0021; #100;
A = 16'h008; B = 16'h0022; #100;
A = 16'h008; B = 16'h0023; #100;
A = 16'h008; B = 16'h0024; #100;
A = 16'h008; B = 16'h0025; #100;
A = 16'h008; B = 16'h0026; #100;
A = 16'h008; B = 16'h0027; #100;
A = 16'h008; B = 16'h0028; #100;
A = 16'h008; B = 16'h0029; #100;
A = 16'h008; B = 16'h002A; #100;
A = 16'h008; B = 16'h002B; #100;
A = 16'h008; B = 16'h002C; #100;
A = 16'h008; B = 16'h002D; #100;
A = 16'h008; B = 16'h002E; #100;
A = 16'h008; B = 16'h002F; #100;
A = 16'h008; B = 16'h0030; #100;
A = 16'h008; B = 16'h0031; #100;
A = 16'h008; B = 16'h0032; #100;
A = 16'h008; B = 16'h0033; #100;
A = 16'h008; B = 16'h0034; #100;
A = 16'h008; B = 16'h0035; #100;
A = 16'h008; B = 16'h0036; #100;
A = 16'h008; B = 16'h0037; #100;
A = 16'h008; B = 16'h0038; #100;
A = 16'h008; B = 16'h0039; #100;
A = 16'h008; B = 16'h003A; #100;
A = 16'h008; B = 16'h003B; #100;
A = 16'h008; B = 16'h003C; #100;
A = 16'h008; B = 16'h003D; #100;
A = 16'h008; B = 16'h003E; #100;
A = 16'h008; B = 16'h003F; #100;
A = 16'h008; B = 16'h0040; #100;
A = 16'h008; B = 16'h0041; #100;
A = 16'h008; B = 16'h0042; #100;
A = 16'h008; B = 16'h0043; #100;
A = 16'h008; B = 16'h0044; #100;
A = 16'h008; B = 16'h0045; #100;
A = 16'h008; B = 16'h0046; #100;
A = 16'h008; B = 16'h0047; #100;
A = 16'h008; B = 16'h0048; #100;
A = 16'h008; B = 16'h0049; #100;
A = 16'h008; B = 16'h004A; #100;
A = 16'h008; B = 16'h004B; #100;
A = 16'h008; B = 16'h004C; #100;
A = 16'h008; B = 16'h004D; #100;
A = 16'h008; B = 16'h004E; #100;
A = 16'h008; B = 16'h004F; #100;
A = 16'h008; B = 16'h0050; #100;
A = 16'h008; B = 16'h0051; #100;
A = 16'h008; B = 16'h0052; #100;
A = 16'h008; B = 16'h0053; #100;
A = 16'h008; B = 16'h0054; #100;
A = 16'h008; B = 16'h0055; #100;
A = 16'h008; B = 16'h0056; #100;
A = 16'h008; B = 16'h0057; #100;
A = 16'h008; B = 16'h0058; #100;
A = 16'h008; B = 16'h0059; #100;
A = 16'h008; B = 16'h005A; #100;
A = 16'h008; B = 16'h005B; #100;
A = 16'h008; B = 16'h005C; #100;
A = 16'h008; B = 16'h005D; #100;
A = 16'h008; B = 16'h005E; #100;
A = 16'h008; B = 16'h005F; #100;
A = 16'h008; B = 16'h0060; #100;
A = 16'h008; B = 16'h0061; #100;
A = 16'h008; B = 16'h0062; #100;
A = 16'h008; B = 16'h0063; #100;
A = 16'h008; B = 16'h0064; #100;
A = 16'h008; B = 16'h0065; #100;
A = 16'h008; B = 16'h0066; #100;
A = 16'h008; B = 16'h0067; #100;
A = 16'h008; B = 16'h0068; #100;
A = 16'h008; B = 16'h0069; #100;
A = 16'h008; B = 16'h006A; #100;
A = 16'h008; B = 16'h006B; #100;
A = 16'h008; B = 16'h006C; #100;
A = 16'h008; B = 16'h006D; #100;
A = 16'h008; B = 16'h006E; #100;
A = 16'h008; B = 16'h006F; #100;
A = 16'h008; B = 16'h0070; #100;
A = 16'h008; B = 16'h0071; #100;
A = 16'h008; B = 16'h0072; #100;
A = 16'h008; B = 16'h0073; #100;
A = 16'h008; B = 16'h0074; #100;
A = 16'h008; B = 16'h0075; #100;
A = 16'h008; B = 16'h0076; #100;
A = 16'h008; B = 16'h0077; #100;
A = 16'h008; B = 16'h0078; #100;
A = 16'h008; B = 16'h0079; #100;
A = 16'h008; B = 16'h007A; #100;
A = 16'h008; B = 16'h007B; #100;
A = 16'h008; B = 16'h007C; #100;
A = 16'h008; B = 16'h007D; #100;
A = 16'h008; B = 16'h007E; #100;
A = 16'h008; B = 16'h007F; #100;
A = 16'h008; B = 16'h0080; #100;
A = 16'h008; B = 16'h0081; #100;
A = 16'h008; B = 16'h0082; #100;
A = 16'h008; B = 16'h0083; #100;
A = 16'h008; B = 16'h0084; #100;
A = 16'h008; B = 16'h0085; #100;
A = 16'h008; B = 16'h0086; #100;
A = 16'h008; B = 16'h0087; #100;
A = 16'h008; B = 16'h0088; #100;
A = 16'h008; B = 16'h0089; #100;
A = 16'h008; B = 16'h008A; #100;
A = 16'h008; B = 16'h008B; #100;
A = 16'h008; B = 16'h008C; #100;
A = 16'h008; B = 16'h008D; #100;
A = 16'h008; B = 16'h008E; #100;
A = 16'h008; B = 16'h008F; #100;
A = 16'h008; B = 16'h0090; #100;
A = 16'h008; B = 16'h0091; #100;
A = 16'h008; B = 16'h0092; #100;
A = 16'h008; B = 16'h0093; #100;
A = 16'h008; B = 16'h0094; #100;
A = 16'h008; B = 16'h0095; #100;
A = 16'h008; B = 16'h0096; #100;
A = 16'h008; B = 16'h0097; #100;
A = 16'h008; B = 16'h0098; #100;
A = 16'h008; B = 16'h0099; #100;
A = 16'h008; B = 16'h009A; #100;
A = 16'h008; B = 16'h009B; #100;
A = 16'h008; B = 16'h009C; #100;
A = 16'h008; B = 16'h009D; #100;
A = 16'h008; B = 16'h009E; #100;
A = 16'h008; B = 16'h009F; #100;
A = 16'h008; B = 16'h00A0; #100;
A = 16'h008; B = 16'h00A1; #100;
A = 16'h008; B = 16'h00A2; #100;
A = 16'h008; B = 16'h00A3; #100;
A = 16'h008; B = 16'h00A4; #100;
A = 16'h008; B = 16'h00A5; #100;
A = 16'h008; B = 16'h00A6; #100;
A = 16'h008; B = 16'h00A7; #100;
A = 16'h008; B = 16'h00A8; #100;
A = 16'h008; B = 16'h00A9; #100;
A = 16'h008; B = 16'h00AA; #100;
A = 16'h008; B = 16'h00AB; #100;
A = 16'h008; B = 16'h00AC; #100;
A = 16'h008; B = 16'h00AD; #100;
A = 16'h008; B = 16'h00AE; #100;
A = 16'h008; B = 16'h00AF; #100;
A = 16'h008; B = 16'h00B0; #100;
A = 16'h008; B = 16'h00B1; #100;
A = 16'h008; B = 16'h00B2; #100;
A = 16'h008; B = 16'h00B3; #100;
A = 16'h008; B = 16'h00B4; #100;
A = 16'h008; B = 16'h00B5; #100;
A = 16'h008; B = 16'h00B6; #100;
A = 16'h008; B = 16'h00B7; #100;
A = 16'h008; B = 16'h00B8; #100;
A = 16'h008; B = 16'h00B9; #100;
A = 16'h008; B = 16'h00BA; #100;
A = 16'h008; B = 16'h00BB; #100;
A = 16'h008; B = 16'h00BC; #100;
A = 16'h008; B = 16'h00BD; #100;
A = 16'h008; B = 16'h00BE; #100;
A = 16'h008; B = 16'h00BF; #100;
A = 16'h008; B = 16'h00C0; #100;
A = 16'h008; B = 16'h00C1; #100;
A = 16'h008; B = 16'h00C2; #100;
A = 16'h008; B = 16'h00C3; #100;
A = 16'h008; B = 16'h00C4; #100;
A = 16'h008; B = 16'h00C5; #100;
A = 16'h008; B = 16'h00C6; #100;
A = 16'h008; B = 16'h00C7; #100;
A = 16'h008; B = 16'h00C8; #100;
A = 16'h008; B = 16'h00C9; #100;
A = 16'h008; B = 16'h00CA; #100;
A = 16'h008; B = 16'h00CB; #100;
A = 16'h008; B = 16'h00CC; #100;
A = 16'h008; B = 16'h00CD; #100;
A = 16'h008; B = 16'h00CE; #100;
A = 16'h008; B = 16'h00CF; #100;
A = 16'h008; B = 16'h00D0; #100;
A = 16'h008; B = 16'h00D1; #100;
A = 16'h008; B = 16'h00D2; #100;
A = 16'h008; B = 16'h00D3; #100;
A = 16'h008; B = 16'h00D4; #100;
A = 16'h008; B = 16'h00D5; #100;
A = 16'h008; B = 16'h00D6; #100;
A = 16'h008; B = 16'h00D7; #100;
A = 16'h008; B = 16'h00D8; #100;
A = 16'h008; B = 16'h00D9; #100;
A = 16'h008; B = 16'h00DA; #100;
A = 16'h008; B = 16'h00DB; #100;
A = 16'h008; B = 16'h00DC; #100;
A = 16'h008; B = 16'h00DD; #100;
A = 16'h008; B = 16'h00DE; #100;
A = 16'h008; B = 16'h00DF; #100;
A = 16'h008; B = 16'h00E0; #100;
A = 16'h008; B = 16'h00E1; #100;
A = 16'h008; B = 16'h00E2; #100;
A = 16'h008; B = 16'h00E3; #100;
A = 16'h008; B = 16'h00E4; #100;
A = 16'h008; B = 16'h00E5; #100;
A = 16'h008; B = 16'h00E6; #100;
A = 16'h008; B = 16'h00E7; #100;
A = 16'h008; B = 16'h00E8; #100;
A = 16'h008; B = 16'h00E9; #100;
A = 16'h008; B = 16'h00EA; #100;
A = 16'h008; B = 16'h00EB; #100;
A = 16'h008; B = 16'h00EC; #100;
A = 16'h008; B = 16'h00ED; #100;
A = 16'h008; B = 16'h00EE; #100;
A = 16'h008; B = 16'h00EF; #100;
A = 16'h008; B = 16'h00F0; #100;
A = 16'h008; B = 16'h00F1; #100;
A = 16'h008; B = 16'h00F2; #100;
A = 16'h008; B = 16'h00F3; #100;
A = 16'h008; B = 16'h00F4; #100;
A = 16'h008; B = 16'h00F5; #100;
A = 16'h008; B = 16'h00F6; #100;
A = 16'h008; B = 16'h00F7; #100;
A = 16'h008; B = 16'h00F8; #100;
A = 16'h008; B = 16'h00F9; #100;
A = 16'h008; B = 16'h00FA; #100;
A = 16'h008; B = 16'h00FB; #100;
A = 16'h008; B = 16'h00FC; #100;
A = 16'h008; B = 16'h00FD; #100;
A = 16'h008; B = 16'h00FE; #100;
A = 16'h008; B = 16'h00FF; #100;
A = 16'h009; B = 16'h000; #100;
A = 16'h009; B = 16'h001; #100;
A = 16'h009; B = 16'h002; #100;
A = 16'h009; B = 16'h003; #100;
A = 16'h009; B = 16'h004; #100;
A = 16'h009; B = 16'h005; #100;
A = 16'h009; B = 16'h006; #100;
A = 16'h009; B = 16'h007; #100;
A = 16'h009; B = 16'h008; #100;
A = 16'h009; B = 16'h009; #100;
A = 16'h009; B = 16'h00A; #100;
A = 16'h009; B = 16'h00B; #100;
A = 16'h009; B = 16'h00C; #100;
A = 16'h009; B = 16'h00D; #100;
A = 16'h009; B = 16'h00E; #100;
A = 16'h009; B = 16'h00F; #100;
A = 16'h009; B = 16'h0010; #100;
A = 16'h009; B = 16'h0011; #100;
A = 16'h009; B = 16'h0012; #100;
A = 16'h009; B = 16'h0013; #100;
A = 16'h009; B = 16'h0014; #100;
A = 16'h009; B = 16'h0015; #100;
A = 16'h009; B = 16'h0016; #100;
A = 16'h009; B = 16'h0017; #100;
A = 16'h009; B = 16'h0018; #100;
A = 16'h009; B = 16'h0019; #100;
A = 16'h009; B = 16'h001A; #100;
A = 16'h009; B = 16'h001B; #100;
A = 16'h009; B = 16'h001C; #100;
A = 16'h009; B = 16'h001D; #100;
A = 16'h009; B = 16'h001E; #100;
A = 16'h009; B = 16'h001F; #100;
A = 16'h009; B = 16'h0020; #100;
A = 16'h009; B = 16'h0021; #100;
A = 16'h009; B = 16'h0022; #100;
A = 16'h009; B = 16'h0023; #100;
A = 16'h009; B = 16'h0024; #100;
A = 16'h009; B = 16'h0025; #100;
A = 16'h009; B = 16'h0026; #100;
A = 16'h009; B = 16'h0027; #100;
A = 16'h009; B = 16'h0028; #100;
A = 16'h009; B = 16'h0029; #100;
A = 16'h009; B = 16'h002A; #100;
A = 16'h009; B = 16'h002B; #100;
A = 16'h009; B = 16'h002C; #100;
A = 16'h009; B = 16'h002D; #100;
A = 16'h009; B = 16'h002E; #100;
A = 16'h009; B = 16'h002F; #100;
A = 16'h009; B = 16'h0030; #100;
A = 16'h009; B = 16'h0031; #100;
A = 16'h009; B = 16'h0032; #100;
A = 16'h009; B = 16'h0033; #100;
A = 16'h009; B = 16'h0034; #100;
A = 16'h009; B = 16'h0035; #100;
A = 16'h009; B = 16'h0036; #100;
A = 16'h009; B = 16'h0037; #100;
A = 16'h009; B = 16'h0038; #100;
A = 16'h009; B = 16'h0039; #100;
A = 16'h009; B = 16'h003A; #100;
A = 16'h009; B = 16'h003B; #100;
A = 16'h009; B = 16'h003C; #100;
A = 16'h009; B = 16'h003D; #100;
A = 16'h009; B = 16'h003E; #100;
A = 16'h009; B = 16'h003F; #100;
A = 16'h009; B = 16'h0040; #100;
A = 16'h009; B = 16'h0041; #100;
A = 16'h009; B = 16'h0042; #100;
A = 16'h009; B = 16'h0043; #100;
A = 16'h009; B = 16'h0044; #100;
A = 16'h009; B = 16'h0045; #100;
A = 16'h009; B = 16'h0046; #100;
A = 16'h009; B = 16'h0047; #100;
A = 16'h009; B = 16'h0048; #100;
A = 16'h009; B = 16'h0049; #100;
A = 16'h009; B = 16'h004A; #100;
A = 16'h009; B = 16'h004B; #100;
A = 16'h009; B = 16'h004C; #100;
A = 16'h009; B = 16'h004D; #100;
A = 16'h009; B = 16'h004E; #100;
A = 16'h009; B = 16'h004F; #100;
A = 16'h009; B = 16'h0050; #100;
A = 16'h009; B = 16'h0051; #100;
A = 16'h009; B = 16'h0052; #100;
A = 16'h009; B = 16'h0053; #100;
A = 16'h009; B = 16'h0054; #100;
A = 16'h009; B = 16'h0055; #100;
A = 16'h009; B = 16'h0056; #100;
A = 16'h009; B = 16'h0057; #100;
A = 16'h009; B = 16'h0058; #100;
A = 16'h009; B = 16'h0059; #100;
A = 16'h009; B = 16'h005A; #100;
A = 16'h009; B = 16'h005B; #100;
A = 16'h009; B = 16'h005C; #100;
A = 16'h009; B = 16'h005D; #100;
A = 16'h009; B = 16'h005E; #100;
A = 16'h009; B = 16'h005F; #100;
A = 16'h009; B = 16'h0060; #100;
A = 16'h009; B = 16'h0061; #100;
A = 16'h009; B = 16'h0062; #100;
A = 16'h009; B = 16'h0063; #100;
A = 16'h009; B = 16'h0064; #100;
A = 16'h009; B = 16'h0065; #100;
A = 16'h009; B = 16'h0066; #100;
A = 16'h009; B = 16'h0067; #100;
A = 16'h009; B = 16'h0068; #100;
A = 16'h009; B = 16'h0069; #100;
A = 16'h009; B = 16'h006A; #100;
A = 16'h009; B = 16'h006B; #100;
A = 16'h009; B = 16'h006C; #100;
A = 16'h009; B = 16'h006D; #100;
A = 16'h009; B = 16'h006E; #100;
A = 16'h009; B = 16'h006F; #100;
A = 16'h009; B = 16'h0070; #100;
A = 16'h009; B = 16'h0071; #100;
A = 16'h009; B = 16'h0072; #100;
A = 16'h009; B = 16'h0073; #100;
A = 16'h009; B = 16'h0074; #100;
A = 16'h009; B = 16'h0075; #100;
A = 16'h009; B = 16'h0076; #100;
A = 16'h009; B = 16'h0077; #100;
A = 16'h009; B = 16'h0078; #100;
A = 16'h009; B = 16'h0079; #100;
A = 16'h009; B = 16'h007A; #100;
A = 16'h009; B = 16'h007B; #100;
A = 16'h009; B = 16'h007C; #100;
A = 16'h009; B = 16'h007D; #100;
A = 16'h009; B = 16'h007E; #100;
A = 16'h009; B = 16'h007F; #100;
A = 16'h009; B = 16'h0080; #100;
A = 16'h009; B = 16'h0081; #100;
A = 16'h009; B = 16'h0082; #100;
A = 16'h009; B = 16'h0083; #100;
A = 16'h009; B = 16'h0084; #100;
A = 16'h009; B = 16'h0085; #100;
A = 16'h009; B = 16'h0086; #100;
A = 16'h009; B = 16'h0087; #100;
A = 16'h009; B = 16'h0088; #100;
A = 16'h009; B = 16'h0089; #100;
A = 16'h009; B = 16'h008A; #100;
A = 16'h009; B = 16'h008B; #100;
A = 16'h009; B = 16'h008C; #100;
A = 16'h009; B = 16'h008D; #100;
A = 16'h009; B = 16'h008E; #100;
A = 16'h009; B = 16'h008F; #100;
A = 16'h009; B = 16'h0090; #100;
A = 16'h009; B = 16'h0091; #100;
A = 16'h009; B = 16'h0092; #100;
A = 16'h009; B = 16'h0093; #100;
A = 16'h009; B = 16'h0094; #100;
A = 16'h009; B = 16'h0095; #100;
A = 16'h009; B = 16'h0096; #100;
A = 16'h009; B = 16'h0097; #100;
A = 16'h009; B = 16'h0098; #100;
A = 16'h009; B = 16'h0099; #100;
A = 16'h009; B = 16'h009A; #100;
A = 16'h009; B = 16'h009B; #100;
A = 16'h009; B = 16'h009C; #100;
A = 16'h009; B = 16'h009D; #100;
A = 16'h009; B = 16'h009E; #100;
A = 16'h009; B = 16'h009F; #100;
A = 16'h009; B = 16'h00A0; #100;
A = 16'h009; B = 16'h00A1; #100;
A = 16'h009; B = 16'h00A2; #100;
A = 16'h009; B = 16'h00A3; #100;
A = 16'h009; B = 16'h00A4; #100;
A = 16'h009; B = 16'h00A5; #100;
A = 16'h009; B = 16'h00A6; #100;
A = 16'h009; B = 16'h00A7; #100;
A = 16'h009; B = 16'h00A8; #100;
A = 16'h009; B = 16'h00A9; #100;
A = 16'h009; B = 16'h00AA; #100;
A = 16'h009; B = 16'h00AB; #100;
A = 16'h009; B = 16'h00AC; #100;
A = 16'h009; B = 16'h00AD; #100;
A = 16'h009; B = 16'h00AE; #100;
A = 16'h009; B = 16'h00AF; #100;
A = 16'h009; B = 16'h00B0; #100;
A = 16'h009; B = 16'h00B1; #100;
A = 16'h009; B = 16'h00B2; #100;
A = 16'h009; B = 16'h00B3; #100;
A = 16'h009; B = 16'h00B4; #100;
A = 16'h009; B = 16'h00B5; #100;
A = 16'h009; B = 16'h00B6; #100;
A = 16'h009; B = 16'h00B7; #100;
A = 16'h009; B = 16'h00B8; #100;
A = 16'h009; B = 16'h00B9; #100;
A = 16'h009; B = 16'h00BA; #100;
A = 16'h009; B = 16'h00BB; #100;
A = 16'h009; B = 16'h00BC; #100;
A = 16'h009; B = 16'h00BD; #100;
A = 16'h009; B = 16'h00BE; #100;
A = 16'h009; B = 16'h00BF; #100;
A = 16'h009; B = 16'h00C0; #100;
A = 16'h009; B = 16'h00C1; #100;
A = 16'h009; B = 16'h00C2; #100;
A = 16'h009; B = 16'h00C3; #100;
A = 16'h009; B = 16'h00C4; #100;
A = 16'h009; B = 16'h00C5; #100;
A = 16'h009; B = 16'h00C6; #100;
A = 16'h009; B = 16'h00C7; #100;
A = 16'h009; B = 16'h00C8; #100;
A = 16'h009; B = 16'h00C9; #100;
A = 16'h009; B = 16'h00CA; #100;
A = 16'h009; B = 16'h00CB; #100;
A = 16'h009; B = 16'h00CC; #100;
A = 16'h009; B = 16'h00CD; #100;
A = 16'h009; B = 16'h00CE; #100;
A = 16'h009; B = 16'h00CF; #100;
A = 16'h009; B = 16'h00D0; #100;
A = 16'h009; B = 16'h00D1; #100;
A = 16'h009; B = 16'h00D2; #100;
A = 16'h009; B = 16'h00D3; #100;
A = 16'h009; B = 16'h00D4; #100;
A = 16'h009; B = 16'h00D5; #100;
A = 16'h009; B = 16'h00D6; #100;
A = 16'h009; B = 16'h00D7; #100;
A = 16'h009; B = 16'h00D8; #100;
A = 16'h009; B = 16'h00D9; #100;
A = 16'h009; B = 16'h00DA; #100;
A = 16'h009; B = 16'h00DB; #100;
A = 16'h009; B = 16'h00DC; #100;
A = 16'h009; B = 16'h00DD; #100;
A = 16'h009; B = 16'h00DE; #100;
A = 16'h009; B = 16'h00DF; #100;
A = 16'h009; B = 16'h00E0; #100;
A = 16'h009; B = 16'h00E1; #100;
A = 16'h009; B = 16'h00E2; #100;
A = 16'h009; B = 16'h00E3; #100;
A = 16'h009; B = 16'h00E4; #100;
A = 16'h009; B = 16'h00E5; #100;
A = 16'h009; B = 16'h00E6; #100;
A = 16'h009; B = 16'h00E7; #100;
A = 16'h009; B = 16'h00E8; #100;
A = 16'h009; B = 16'h00E9; #100;
A = 16'h009; B = 16'h00EA; #100;
A = 16'h009; B = 16'h00EB; #100;
A = 16'h009; B = 16'h00EC; #100;
A = 16'h009; B = 16'h00ED; #100;
A = 16'h009; B = 16'h00EE; #100;
A = 16'h009; B = 16'h00EF; #100;
A = 16'h009; B = 16'h00F0; #100;
A = 16'h009; B = 16'h00F1; #100;
A = 16'h009; B = 16'h00F2; #100;
A = 16'h009; B = 16'h00F3; #100;
A = 16'h009; B = 16'h00F4; #100;
A = 16'h009; B = 16'h00F5; #100;
A = 16'h009; B = 16'h00F6; #100;
A = 16'h009; B = 16'h00F7; #100;
A = 16'h009; B = 16'h00F8; #100;
A = 16'h009; B = 16'h00F9; #100;
A = 16'h009; B = 16'h00FA; #100;
A = 16'h009; B = 16'h00FB; #100;
A = 16'h009; B = 16'h00FC; #100;
A = 16'h009; B = 16'h00FD; #100;
A = 16'h009; B = 16'h00FE; #100;
A = 16'h009; B = 16'h00FF; #100;
A = 16'h00A; B = 16'h000; #100;
A = 16'h00A; B = 16'h001; #100;
A = 16'h00A; B = 16'h002; #100;
A = 16'h00A; B = 16'h003; #100;
A = 16'h00A; B = 16'h004; #100;
A = 16'h00A; B = 16'h005; #100;
A = 16'h00A; B = 16'h006; #100;
A = 16'h00A; B = 16'h007; #100;
A = 16'h00A; B = 16'h008; #100;
A = 16'h00A; B = 16'h009; #100;
A = 16'h00A; B = 16'h00A; #100;
A = 16'h00A; B = 16'h00B; #100;
A = 16'h00A; B = 16'h00C; #100;
A = 16'h00A; B = 16'h00D; #100;
A = 16'h00A; B = 16'h00E; #100;
A = 16'h00A; B = 16'h00F; #100;
A = 16'h00A; B = 16'h0010; #100;
A = 16'h00A; B = 16'h0011; #100;
A = 16'h00A; B = 16'h0012; #100;
A = 16'h00A; B = 16'h0013; #100;
A = 16'h00A; B = 16'h0014; #100;
A = 16'h00A; B = 16'h0015; #100;
A = 16'h00A; B = 16'h0016; #100;
A = 16'h00A; B = 16'h0017; #100;
A = 16'h00A; B = 16'h0018; #100;
A = 16'h00A; B = 16'h0019; #100;
A = 16'h00A; B = 16'h001A; #100;
A = 16'h00A; B = 16'h001B; #100;
A = 16'h00A; B = 16'h001C; #100;
A = 16'h00A; B = 16'h001D; #100;
A = 16'h00A; B = 16'h001E; #100;
A = 16'h00A; B = 16'h001F; #100;
A = 16'h00A; B = 16'h0020; #100;
A = 16'h00A; B = 16'h0021; #100;
A = 16'h00A; B = 16'h0022; #100;
A = 16'h00A; B = 16'h0023; #100;
A = 16'h00A; B = 16'h0024; #100;
A = 16'h00A; B = 16'h0025; #100;
A = 16'h00A; B = 16'h0026; #100;
A = 16'h00A; B = 16'h0027; #100;
A = 16'h00A; B = 16'h0028; #100;
A = 16'h00A; B = 16'h0029; #100;
A = 16'h00A; B = 16'h002A; #100;
A = 16'h00A; B = 16'h002B; #100;
A = 16'h00A; B = 16'h002C; #100;
A = 16'h00A; B = 16'h002D; #100;
A = 16'h00A; B = 16'h002E; #100;
A = 16'h00A; B = 16'h002F; #100;
A = 16'h00A; B = 16'h0030; #100;
A = 16'h00A; B = 16'h0031; #100;
A = 16'h00A; B = 16'h0032; #100;
A = 16'h00A; B = 16'h0033; #100;
A = 16'h00A; B = 16'h0034; #100;
A = 16'h00A; B = 16'h0035; #100;
A = 16'h00A; B = 16'h0036; #100;
A = 16'h00A; B = 16'h0037; #100;
A = 16'h00A; B = 16'h0038; #100;
A = 16'h00A; B = 16'h0039; #100;
A = 16'h00A; B = 16'h003A; #100;
A = 16'h00A; B = 16'h003B; #100;
A = 16'h00A; B = 16'h003C; #100;
A = 16'h00A; B = 16'h003D; #100;
A = 16'h00A; B = 16'h003E; #100;
A = 16'h00A; B = 16'h003F; #100;
A = 16'h00A; B = 16'h0040; #100;
A = 16'h00A; B = 16'h0041; #100;
A = 16'h00A; B = 16'h0042; #100;
A = 16'h00A; B = 16'h0043; #100;
A = 16'h00A; B = 16'h0044; #100;
A = 16'h00A; B = 16'h0045; #100;
A = 16'h00A; B = 16'h0046; #100;
A = 16'h00A; B = 16'h0047; #100;
A = 16'h00A; B = 16'h0048; #100;
A = 16'h00A; B = 16'h0049; #100;
A = 16'h00A; B = 16'h004A; #100;
A = 16'h00A; B = 16'h004B; #100;
A = 16'h00A; B = 16'h004C; #100;
A = 16'h00A; B = 16'h004D; #100;
A = 16'h00A; B = 16'h004E; #100;
A = 16'h00A; B = 16'h004F; #100;
A = 16'h00A; B = 16'h0050; #100;
A = 16'h00A; B = 16'h0051; #100;
A = 16'h00A; B = 16'h0052; #100;
A = 16'h00A; B = 16'h0053; #100;
A = 16'h00A; B = 16'h0054; #100;
A = 16'h00A; B = 16'h0055; #100;
A = 16'h00A; B = 16'h0056; #100;
A = 16'h00A; B = 16'h0057; #100;
A = 16'h00A; B = 16'h0058; #100;
A = 16'h00A; B = 16'h0059; #100;
A = 16'h00A; B = 16'h005A; #100;
A = 16'h00A; B = 16'h005B; #100;
A = 16'h00A; B = 16'h005C; #100;
A = 16'h00A; B = 16'h005D; #100;
A = 16'h00A; B = 16'h005E; #100;
A = 16'h00A; B = 16'h005F; #100;
A = 16'h00A; B = 16'h0060; #100;
A = 16'h00A; B = 16'h0061; #100;
A = 16'h00A; B = 16'h0062; #100;
A = 16'h00A; B = 16'h0063; #100;
A = 16'h00A; B = 16'h0064; #100;
A = 16'h00A; B = 16'h0065; #100;
A = 16'h00A; B = 16'h0066; #100;
A = 16'h00A; B = 16'h0067; #100;
A = 16'h00A; B = 16'h0068; #100;
A = 16'h00A; B = 16'h0069; #100;
A = 16'h00A; B = 16'h006A; #100;
A = 16'h00A; B = 16'h006B; #100;
A = 16'h00A; B = 16'h006C; #100;
A = 16'h00A; B = 16'h006D; #100;
A = 16'h00A; B = 16'h006E; #100;
A = 16'h00A; B = 16'h006F; #100;
A = 16'h00A; B = 16'h0070; #100;
A = 16'h00A; B = 16'h0071; #100;
A = 16'h00A; B = 16'h0072; #100;
A = 16'h00A; B = 16'h0073; #100;
A = 16'h00A; B = 16'h0074; #100;
A = 16'h00A; B = 16'h0075; #100;
A = 16'h00A; B = 16'h0076; #100;
A = 16'h00A; B = 16'h0077; #100;
A = 16'h00A; B = 16'h0078; #100;
A = 16'h00A; B = 16'h0079; #100;
A = 16'h00A; B = 16'h007A; #100;
A = 16'h00A; B = 16'h007B; #100;
A = 16'h00A; B = 16'h007C; #100;
A = 16'h00A; B = 16'h007D; #100;
A = 16'h00A; B = 16'h007E; #100;
A = 16'h00A; B = 16'h007F; #100;
A = 16'h00A; B = 16'h0080; #100;
A = 16'h00A; B = 16'h0081; #100;
A = 16'h00A; B = 16'h0082; #100;
A = 16'h00A; B = 16'h0083; #100;
A = 16'h00A; B = 16'h0084; #100;
A = 16'h00A; B = 16'h0085; #100;
A = 16'h00A; B = 16'h0086; #100;
A = 16'h00A; B = 16'h0087; #100;
A = 16'h00A; B = 16'h0088; #100;
A = 16'h00A; B = 16'h0089; #100;
A = 16'h00A; B = 16'h008A; #100;
A = 16'h00A; B = 16'h008B; #100;
A = 16'h00A; B = 16'h008C; #100;
A = 16'h00A; B = 16'h008D; #100;
A = 16'h00A; B = 16'h008E; #100;
A = 16'h00A; B = 16'h008F; #100;
A = 16'h00A; B = 16'h0090; #100;
A = 16'h00A; B = 16'h0091; #100;
A = 16'h00A; B = 16'h0092; #100;
A = 16'h00A; B = 16'h0093; #100;
A = 16'h00A; B = 16'h0094; #100;
A = 16'h00A; B = 16'h0095; #100;
A = 16'h00A; B = 16'h0096; #100;
A = 16'h00A; B = 16'h0097; #100;
A = 16'h00A; B = 16'h0098; #100;
A = 16'h00A; B = 16'h0099; #100;
A = 16'h00A; B = 16'h009A; #100;
A = 16'h00A; B = 16'h009B; #100;
A = 16'h00A; B = 16'h009C; #100;
A = 16'h00A; B = 16'h009D; #100;
A = 16'h00A; B = 16'h009E; #100;
A = 16'h00A; B = 16'h009F; #100;
A = 16'h00A; B = 16'h00A0; #100;
A = 16'h00A; B = 16'h00A1; #100;
A = 16'h00A; B = 16'h00A2; #100;
A = 16'h00A; B = 16'h00A3; #100;
A = 16'h00A; B = 16'h00A4; #100;
A = 16'h00A; B = 16'h00A5; #100;
A = 16'h00A; B = 16'h00A6; #100;
A = 16'h00A; B = 16'h00A7; #100;
A = 16'h00A; B = 16'h00A8; #100;
A = 16'h00A; B = 16'h00A9; #100;
A = 16'h00A; B = 16'h00AA; #100;
A = 16'h00A; B = 16'h00AB; #100;
A = 16'h00A; B = 16'h00AC; #100;
A = 16'h00A; B = 16'h00AD; #100;
A = 16'h00A; B = 16'h00AE; #100;
A = 16'h00A; B = 16'h00AF; #100;
A = 16'h00A; B = 16'h00B0; #100;
A = 16'h00A; B = 16'h00B1; #100;
A = 16'h00A; B = 16'h00B2; #100;
A = 16'h00A; B = 16'h00B3; #100;
A = 16'h00A; B = 16'h00B4; #100;
A = 16'h00A; B = 16'h00B5; #100;
A = 16'h00A; B = 16'h00B6; #100;
A = 16'h00A; B = 16'h00B7; #100;
A = 16'h00A; B = 16'h00B8; #100;
A = 16'h00A; B = 16'h00B9; #100;
A = 16'h00A; B = 16'h00BA; #100;
A = 16'h00A; B = 16'h00BB; #100;
A = 16'h00A; B = 16'h00BC; #100;
A = 16'h00A; B = 16'h00BD; #100;
A = 16'h00A; B = 16'h00BE; #100;
A = 16'h00A; B = 16'h00BF; #100;
A = 16'h00A; B = 16'h00C0; #100;
A = 16'h00A; B = 16'h00C1; #100;
A = 16'h00A; B = 16'h00C2; #100;
A = 16'h00A; B = 16'h00C3; #100;
A = 16'h00A; B = 16'h00C4; #100;
A = 16'h00A; B = 16'h00C5; #100;
A = 16'h00A; B = 16'h00C6; #100;
A = 16'h00A; B = 16'h00C7; #100;
A = 16'h00A; B = 16'h00C8; #100;
A = 16'h00A; B = 16'h00C9; #100;
A = 16'h00A; B = 16'h00CA; #100;
A = 16'h00A; B = 16'h00CB; #100;
A = 16'h00A; B = 16'h00CC; #100;
A = 16'h00A; B = 16'h00CD; #100;
A = 16'h00A; B = 16'h00CE; #100;
A = 16'h00A; B = 16'h00CF; #100;
A = 16'h00A; B = 16'h00D0; #100;
A = 16'h00A; B = 16'h00D1; #100;
A = 16'h00A; B = 16'h00D2; #100;
A = 16'h00A; B = 16'h00D3; #100;
A = 16'h00A; B = 16'h00D4; #100;
A = 16'h00A; B = 16'h00D5; #100;
A = 16'h00A; B = 16'h00D6; #100;
A = 16'h00A; B = 16'h00D7; #100;
A = 16'h00A; B = 16'h00D8; #100;
A = 16'h00A; B = 16'h00D9; #100;
A = 16'h00A; B = 16'h00DA; #100;
A = 16'h00A; B = 16'h00DB; #100;
A = 16'h00A; B = 16'h00DC; #100;
A = 16'h00A; B = 16'h00DD; #100;
A = 16'h00A; B = 16'h00DE; #100;
A = 16'h00A; B = 16'h00DF; #100;
A = 16'h00A; B = 16'h00E0; #100;
A = 16'h00A; B = 16'h00E1; #100;
A = 16'h00A; B = 16'h00E2; #100;
A = 16'h00A; B = 16'h00E3; #100;
A = 16'h00A; B = 16'h00E4; #100;
A = 16'h00A; B = 16'h00E5; #100;
A = 16'h00A; B = 16'h00E6; #100;
A = 16'h00A; B = 16'h00E7; #100;
A = 16'h00A; B = 16'h00E8; #100;
A = 16'h00A; B = 16'h00E9; #100;
A = 16'h00A; B = 16'h00EA; #100;
A = 16'h00A; B = 16'h00EB; #100;
A = 16'h00A; B = 16'h00EC; #100;
A = 16'h00A; B = 16'h00ED; #100;
A = 16'h00A; B = 16'h00EE; #100;
A = 16'h00A; B = 16'h00EF; #100;
A = 16'h00A; B = 16'h00F0; #100;
A = 16'h00A; B = 16'h00F1; #100;
A = 16'h00A; B = 16'h00F2; #100;
A = 16'h00A; B = 16'h00F3; #100;
A = 16'h00A; B = 16'h00F4; #100;
A = 16'h00A; B = 16'h00F5; #100;
A = 16'h00A; B = 16'h00F6; #100;
A = 16'h00A; B = 16'h00F7; #100;
A = 16'h00A; B = 16'h00F8; #100;
A = 16'h00A; B = 16'h00F9; #100;
A = 16'h00A; B = 16'h00FA; #100;
A = 16'h00A; B = 16'h00FB; #100;
A = 16'h00A; B = 16'h00FC; #100;
A = 16'h00A; B = 16'h00FD; #100;
A = 16'h00A; B = 16'h00FE; #100;
A = 16'h00A; B = 16'h00FF; #100;
A = 16'h00B; B = 16'h000; #100;
A = 16'h00B; B = 16'h001; #100;
A = 16'h00B; B = 16'h002; #100;
A = 16'h00B; B = 16'h003; #100;
A = 16'h00B; B = 16'h004; #100;
A = 16'h00B; B = 16'h005; #100;
A = 16'h00B; B = 16'h006; #100;
A = 16'h00B; B = 16'h007; #100;
A = 16'h00B; B = 16'h008; #100;
A = 16'h00B; B = 16'h009; #100;
A = 16'h00B; B = 16'h00A; #100;
A = 16'h00B; B = 16'h00B; #100;
A = 16'h00B; B = 16'h00C; #100;
A = 16'h00B; B = 16'h00D; #100;
A = 16'h00B; B = 16'h00E; #100;
A = 16'h00B; B = 16'h00F; #100;
A = 16'h00B; B = 16'h0010; #100;
A = 16'h00B; B = 16'h0011; #100;
A = 16'h00B; B = 16'h0012; #100;
A = 16'h00B; B = 16'h0013; #100;
A = 16'h00B; B = 16'h0014; #100;
A = 16'h00B; B = 16'h0015; #100;
A = 16'h00B; B = 16'h0016; #100;
A = 16'h00B; B = 16'h0017; #100;
A = 16'h00B; B = 16'h0018; #100;
A = 16'h00B; B = 16'h0019; #100;
A = 16'h00B; B = 16'h001A; #100;
A = 16'h00B; B = 16'h001B; #100;
A = 16'h00B; B = 16'h001C; #100;
A = 16'h00B; B = 16'h001D; #100;
A = 16'h00B; B = 16'h001E; #100;
A = 16'h00B; B = 16'h001F; #100;
A = 16'h00B; B = 16'h0020; #100;
A = 16'h00B; B = 16'h0021; #100;
A = 16'h00B; B = 16'h0022; #100;
A = 16'h00B; B = 16'h0023; #100;
A = 16'h00B; B = 16'h0024; #100;
A = 16'h00B; B = 16'h0025; #100;
A = 16'h00B; B = 16'h0026; #100;
A = 16'h00B; B = 16'h0027; #100;
A = 16'h00B; B = 16'h0028; #100;
A = 16'h00B; B = 16'h0029; #100;
A = 16'h00B; B = 16'h002A; #100;
A = 16'h00B; B = 16'h002B; #100;
A = 16'h00B; B = 16'h002C; #100;
A = 16'h00B; B = 16'h002D; #100;
A = 16'h00B; B = 16'h002E; #100;
A = 16'h00B; B = 16'h002F; #100;
A = 16'h00B; B = 16'h0030; #100;
A = 16'h00B; B = 16'h0031; #100;
A = 16'h00B; B = 16'h0032; #100;
A = 16'h00B; B = 16'h0033; #100;
A = 16'h00B; B = 16'h0034; #100;
A = 16'h00B; B = 16'h0035; #100;
A = 16'h00B; B = 16'h0036; #100;
A = 16'h00B; B = 16'h0037; #100;
A = 16'h00B; B = 16'h0038; #100;
A = 16'h00B; B = 16'h0039; #100;
A = 16'h00B; B = 16'h003A; #100;
A = 16'h00B; B = 16'h003B; #100;
A = 16'h00B; B = 16'h003C; #100;
A = 16'h00B; B = 16'h003D; #100;
A = 16'h00B; B = 16'h003E; #100;
A = 16'h00B; B = 16'h003F; #100;
A = 16'h00B; B = 16'h0040; #100;
A = 16'h00B; B = 16'h0041; #100;
A = 16'h00B; B = 16'h0042; #100;
A = 16'h00B; B = 16'h0043; #100;
A = 16'h00B; B = 16'h0044; #100;
A = 16'h00B; B = 16'h0045; #100;
A = 16'h00B; B = 16'h0046; #100;
A = 16'h00B; B = 16'h0047; #100;
A = 16'h00B; B = 16'h0048; #100;
A = 16'h00B; B = 16'h0049; #100;
A = 16'h00B; B = 16'h004A; #100;
A = 16'h00B; B = 16'h004B; #100;
A = 16'h00B; B = 16'h004C; #100;
A = 16'h00B; B = 16'h004D; #100;
A = 16'h00B; B = 16'h004E; #100;
A = 16'h00B; B = 16'h004F; #100;
A = 16'h00B; B = 16'h0050; #100;
A = 16'h00B; B = 16'h0051; #100;
A = 16'h00B; B = 16'h0052; #100;
A = 16'h00B; B = 16'h0053; #100;
A = 16'h00B; B = 16'h0054; #100;
A = 16'h00B; B = 16'h0055; #100;
A = 16'h00B; B = 16'h0056; #100;
A = 16'h00B; B = 16'h0057; #100;
A = 16'h00B; B = 16'h0058; #100;
A = 16'h00B; B = 16'h0059; #100;
A = 16'h00B; B = 16'h005A; #100;
A = 16'h00B; B = 16'h005B; #100;
A = 16'h00B; B = 16'h005C; #100;
A = 16'h00B; B = 16'h005D; #100;
A = 16'h00B; B = 16'h005E; #100;
A = 16'h00B; B = 16'h005F; #100;
A = 16'h00B; B = 16'h0060; #100;
A = 16'h00B; B = 16'h0061; #100;
A = 16'h00B; B = 16'h0062; #100;
A = 16'h00B; B = 16'h0063; #100;
A = 16'h00B; B = 16'h0064; #100;
A = 16'h00B; B = 16'h0065; #100;
A = 16'h00B; B = 16'h0066; #100;
A = 16'h00B; B = 16'h0067; #100;
A = 16'h00B; B = 16'h0068; #100;
A = 16'h00B; B = 16'h0069; #100;
A = 16'h00B; B = 16'h006A; #100;
A = 16'h00B; B = 16'h006B; #100;
A = 16'h00B; B = 16'h006C; #100;
A = 16'h00B; B = 16'h006D; #100;
A = 16'h00B; B = 16'h006E; #100;
A = 16'h00B; B = 16'h006F; #100;
A = 16'h00B; B = 16'h0070; #100;
A = 16'h00B; B = 16'h0071; #100;
A = 16'h00B; B = 16'h0072; #100;
A = 16'h00B; B = 16'h0073; #100;
A = 16'h00B; B = 16'h0074; #100;
A = 16'h00B; B = 16'h0075; #100;
A = 16'h00B; B = 16'h0076; #100;
A = 16'h00B; B = 16'h0077; #100;
A = 16'h00B; B = 16'h0078; #100;
A = 16'h00B; B = 16'h0079; #100;
A = 16'h00B; B = 16'h007A; #100;
A = 16'h00B; B = 16'h007B; #100;
A = 16'h00B; B = 16'h007C; #100;
A = 16'h00B; B = 16'h007D; #100;
A = 16'h00B; B = 16'h007E; #100;
A = 16'h00B; B = 16'h007F; #100;
A = 16'h00B; B = 16'h0080; #100;
A = 16'h00B; B = 16'h0081; #100;
A = 16'h00B; B = 16'h0082; #100;
A = 16'h00B; B = 16'h0083; #100;
A = 16'h00B; B = 16'h0084; #100;
A = 16'h00B; B = 16'h0085; #100;
A = 16'h00B; B = 16'h0086; #100;
A = 16'h00B; B = 16'h0087; #100;
A = 16'h00B; B = 16'h0088; #100;
A = 16'h00B; B = 16'h0089; #100;
A = 16'h00B; B = 16'h008A; #100;
A = 16'h00B; B = 16'h008B; #100;
A = 16'h00B; B = 16'h008C; #100;
A = 16'h00B; B = 16'h008D; #100;
A = 16'h00B; B = 16'h008E; #100;
A = 16'h00B; B = 16'h008F; #100;
A = 16'h00B; B = 16'h0090; #100;
A = 16'h00B; B = 16'h0091; #100;
A = 16'h00B; B = 16'h0092; #100;
A = 16'h00B; B = 16'h0093; #100;
A = 16'h00B; B = 16'h0094; #100;
A = 16'h00B; B = 16'h0095; #100;
A = 16'h00B; B = 16'h0096; #100;
A = 16'h00B; B = 16'h0097; #100;
A = 16'h00B; B = 16'h0098; #100;
A = 16'h00B; B = 16'h0099; #100;
A = 16'h00B; B = 16'h009A; #100;
A = 16'h00B; B = 16'h009B; #100;
A = 16'h00B; B = 16'h009C; #100;
A = 16'h00B; B = 16'h009D; #100;
A = 16'h00B; B = 16'h009E; #100;
A = 16'h00B; B = 16'h009F; #100;
A = 16'h00B; B = 16'h00A0; #100;
A = 16'h00B; B = 16'h00A1; #100;
A = 16'h00B; B = 16'h00A2; #100;
A = 16'h00B; B = 16'h00A3; #100;
A = 16'h00B; B = 16'h00A4; #100;
A = 16'h00B; B = 16'h00A5; #100;
A = 16'h00B; B = 16'h00A6; #100;
A = 16'h00B; B = 16'h00A7; #100;
A = 16'h00B; B = 16'h00A8; #100;
A = 16'h00B; B = 16'h00A9; #100;
A = 16'h00B; B = 16'h00AA; #100;
A = 16'h00B; B = 16'h00AB; #100;
A = 16'h00B; B = 16'h00AC; #100;
A = 16'h00B; B = 16'h00AD; #100;
A = 16'h00B; B = 16'h00AE; #100;
A = 16'h00B; B = 16'h00AF; #100;
A = 16'h00B; B = 16'h00B0; #100;
A = 16'h00B; B = 16'h00B1; #100;
A = 16'h00B; B = 16'h00B2; #100;
A = 16'h00B; B = 16'h00B3; #100;
A = 16'h00B; B = 16'h00B4; #100;
A = 16'h00B; B = 16'h00B5; #100;
A = 16'h00B; B = 16'h00B6; #100;
A = 16'h00B; B = 16'h00B7; #100;
A = 16'h00B; B = 16'h00B8; #100;
A = 16'h00B; B = 16'h00B9; #100;
A = 16'h00B; B = 16'h00BA; #100;
A = 16'h00B; B = 16'h00BB; #100;
A = 16'h00B; B = 16'h00BC; #100;
A = 16'h00B; B = 16'h00BD; #100;
A = 16'h00B; B = 16'h00BE; #100;
A = 16'h00B; B = 16'h00BF; #100;
A = 16'h00B; B = 16'h00C0; #100;
A = 16'h00B; B = 16'h00C1; #100;
A = 16'h00B; B = 16'h00C2; #100;
A = 16'h00B; B = 16'h00C3; #100;
A = 16'h00B; B = 16'h00C4; #100;
A = 16'h00B; B = 16'h00C5; #100;
A = 16'h00B; B = 16'h00C6; #100;
A = 16'h00B; B = 16'h00C7; #100;
A = 16'h00B; B = 16'h00C8; #100;
A = 16'h00B; B = 16'h00C9; #100;
A = 16'h00B; B = 16'h00CA; #100;
A = 16'h00B; B = 16'h00CB; #100;
A = 16'h00B; B = 16'h00CC; #100;
A = 16'h00B; B = 16'h00CD; #100;
A = 16'h00B; B = 16'h00CE; #100;
A = 16'h00B; B = 16'h00CF; #100;
A = 16'h00B; B = 16'h00D0; #100;
A = 16'h00B; B = 16'h00D1; #100;
A = 16'h00B; B = 16'h00D2; #100;
A = 16'h00B; B = 16'h00D3; #100;
A = 16'h00B; B = 16'h00D4; #100;
A = 16'h00B; B = 16'h00D5; #100;
A = 16'h00B; B = 16'h00D6; #100;
A = 16'h00B; B = 16'h00D7; #100;
A = 16'h00B; B = 16'h00D8; #100;
A = 16'h00B; B = 16'h00D9; #100;
A = 16'h00B; B = 16'h00DA; #100;
A = 16'h00B; B = 16'h00DB; #100;
A = 16'h00B; B = 16'h00DC; #100;
A = 16'h00B; B = 16'h00DD; #100;
A = 16'h00B; B = 16'h00DE; #100;
A = 16'h00B; B = 16'h00DF; #100;
A = 16'h00B; B = 16'h00E0; #100;
A = 16'h00B; B = 16'h00E1; #100;
A = 16'h00B; B = 16'h00E2; #100;
A = 16'h00B; B = 16'h00E3; #100;
A = 16'h00B; B = 16'h00E4; #100;
A = 16'h00B; B = 16'h00E5; #100;
A = 16'h00B; B = 16'h00E6; #100;
A = 16'h00B; B = 16'h00E7; #100;
A = 16'h00B; B = 16'h00E8; #100;
A = 16'h00B; B = 16'h00E9; #100;
A = 16'h00B; B = 16'h00EA; #100;
A = 16'h00B; B = 16'h00EB; #100;
A = 16'h00B; B = 16'h00EC; #100;
A = 16'h00B; B = 16'h00ED; #100;
A = 16'h00B; B = 16'h00EE; #100;
A = 16'h00B; B = 16'h00EF; #100;
A = 16'h00B; B = 16'h00F0; #100;
A = 16'h00B; B = 16'h00F1; #100;
A = 16'h00B; B = 16'h00F2; #100;
A = 16'h00B; B = 16'h00F3; #100;
A = 16'h00B; B = 16'h00F4; #100;
A = 16'h00B; B = 16'h00F5; #100;
A = 16'h00B; B = 16'h00F6; #100;
A = 16'h00B; B = 16'h00F7; #100;
A = 16'h00B; B = 16'h00F8; #100;
A = 16'h00B; B = 16'h00F9; #100;
A = 16'h00B; B = 16'h00FA; #100;
A = 16'h00B; B = 16'h00FB; #100;
A = 16'h00B; B = 16'h00FC; #100;
A = 16'h00B; B = 16'h00FD; #100;
A = 16'h00B; B = 16'h00FE; #100;
A = 16'h00B; B = 16'h00FF; #100;
A = 16'h00C; B = 16'h000; #100;
A = 16'h00C; B = 16'h001; #100;
A = 16'h00C; B = 16'h002; #100;
A = 16'h00C; B = 16'h003; #100;
A = 16'h00C; B = 16'h004; #100;
A = 16'h00C; B = 16'h005; #100;
A = 16'h00C; B = 16'h006; #100;
A = 16'h00C; B = 16'h007; #100;
A = 16'h00C; B = 16'h008; #100;
A = 16'h00C; B = 16'h009; #100;
A = 16'h00C; B = 16'h00A; #100;
A = 16'h00C; B = 16'h00B; #100;
A = 16'h00C; B = 16'h00C; #100;
A = 16'h00C; B = 16'h00D; #100;
A = 16'h00C; B = 16'h00E; #100;
A = 16'h00C; B = 16'h00F; #100;
A = 16'h00C; B = 16'h0010; #100;
A = 16'h00C; B = 16'h0011; #100;
A = 16'h00C; B = 16'h0012; #100;
A = 16'h00C; B = 16'h0013; #100;
A = 16'h00C; B = 16'h0014; #100;
A = 16'h00C; B = 16'h0015; #100;
A = 16'h00C; B = 16'h0016; #100;
A = 16'h00C; B = 16'h0017; #100;
A = 16'h00C; B = 16'h0018; #100;
A = 16'h00C; B = 16'h0019; #100;
A = 16'h00C; B = 16'h001A; #100;
A = 16'h00C; B = 16'h001B; #100;
A = 16'h00C; B = 16'h001C; #100;
A = 16'h00C; B = 16'h001D; #100;
A = 16'h00C; B = 16'h001E; #100;
A = 16'h00C; B = 16'h001F; #100;
A = 16'h00C; B = 16'h0020; #100;
A = 16'h00C; B = 16'h0021; #100;
A = 16'h00C; B = 16'h0022; #100;
A = 16'h00C; B = 16'h0023; #100;
A = 16'h00C; B = 16'h0024; #100;
A = 16'h00C; B = 16'h0025; #100;
A = 16'h00C; B = 16'h0026; #100;
A = 16'h00C; B = 16'h0027; #100;
A = 16'h00C; B = 16'h0028; #100;
A = 16'h00C; B = 16'h0029; #100;
A = 16'h00C; B = 16'h002A; #100;
A = 16'h00C; B = 16'h002B; #100;
A = 16'h00C; B = 16'h002C; #100;
A = 16'h00C; B = 16'h002D; #100;
A = 16'h00C; B = 16'h002E; #100;
A = 16'h00C; B = 16'h002F; #100;
A = 16'h00C; B = 16'h0030; #100;
A = 16'h00C; B = 16'h0031; #100;
A = 16'h00C; B = 16'h0032; #100;
A = 16'h00C; B = 16'h0033; #100;
A = 16'h00C; B = 16'h0034; #100;
A = 16'h00C; B = 16'h0035; #100;
A = 16'h00C; B = 16'h0036; #100;
A = 16'h00C; B = 16'h0037; #100;
A = 16'h00C; B = 16'h0038; #100;
A = 16'h00C; B = 16'h0039; #100;
A = 16'h00C; B = 16'h003A; #100;
A = 16'h00C; B = 16'h003B; #100;
A = 16'h00C; B = 16'h003C; #100;
A = 16'h00C; B = 16'h003D; #100;
A = 16'h00C; B = 16'h003E; #100;
A = 16'h00C; B = 16'h003F; #100;
A = 16'h00C; B = 16'h0040; #100;
A = 16'h00C; B = 16'h0041; #100;
A = 16'h00C; B = 16'h0042; #100;
A = 16'h00C; B = 16'h0043; #100;
A = 16'h00C; B = 16'h0044; #100;
A = 16'h00C; B = 16'h0045; #100;
A = 16'h00C; B = 16'h0046; #100;
A = 16'h00C; B = 16'h0047; #100;
A = 16'h00C; B = 16'h0048; #100;
A = 16'h00C; B = 16'h0049; #100;
A = 16'h00C; B = 16'h004A; #100;
A = 16'h00C; B = 16'h004B; #100;
A = 16'h00C; B = 16'h004C; #100;
A = 16'h00C; B = 16'h004D; #100;
A = 16'h00C; B = 16'h004E; #100;
A = 16'h00C; B = 16'h004F; #100;
A = 16'h00C; B = 16'h0050; #100;
A = 16'h00C; B = 16'h0051; #100;
A = 16'h00C; B = 16'h0052; #100;
A = 16'h00C; B = 16'h0053; #100;
A = 16'h00C; B = 16'h0054; #100;
A = 16'h00C; B = 16'h0055; #100;
A = 16'h00C; B = 16'h0056; #100;
A = 16'h00C; B = 16'h0057; #100;
A = 16'h00C; B = 16'h0058; #100;
A = 16'h00C; B = 16'h0059; #100;
A = 16'h00C; B = 16'h005A; #100;
A = 16'h00C; B = 16'h005B; #100;
A = 16'h00C; B = 16'h005C; #100;
A = 16'h00C; B = 16'h005D; #100;
A = 16'h00C; B = 16'h005E; #100;
A = 16'h00C; B = 16'h005F; #100;
A = 16'h00C; B = 16'h0060; #100;
A = 16'h00C; B = 16'h0061; #100;
A = 16'h00C; B = 16'h0062; #100;
A = 16'h00C; B = 16'h0063; #100;
A = 16'h00C; B = 16'h0064; #100;
A = 16'h00C; B = 16'h0065; #100;
A = 16'h00C; B = 16'h0066; #100;
A = 16'h00C; B = 16'h0067; #100;
A = 16'h00C; B = 16'h0068; #100;
A = 16'h00C; B = 16'h0069; #100;
A = 16'h00C; B = 16'h006A; #100;
A = 16'h00C; B = 16'h006B; #100;
A = 16'h00C; B = 16'h006C; #100;
A = 16'h00C; B = 16'h006D; #100;
A = 16'h00C; B = 16'h006E; #100;
A = 16'h00C; B = 16'h006F; #100;
A = 16'h00C; B = 16'h0070; #100;
A = 16'h00C; B = 16'h0071; #100;
A = 16'h00C; B = 16'h0072; #100;
A = 16'h00C; B = 16'h0073; #100;
A = 16'h00C; B = 16'h0074; #100;
A = 16'h00C; B = 16'h0075; #100;
A = 16'h00C; B = 16'h0076; #100;
A = 16'h00C; B = 16'h0077; #100;
A = 16'h00C; B = 16'h0078; #100;
A = 16'h00C; B = 16'h0079; #100;
A = 16'h00C; B = 16'h007A; #100;
A = 16'h00C; B = 16'h007B; #100;
A = 16'h00C; B = 16'h007C; #100;
A = 16'h00C; B = 16'h007D; #100;
A = 16'h00C; B = 16'h007E; #100;
A = 16'h00C; B = 16'h007F; #100;
A = 16'h00C; B = 16'h0080; #100;
A = 16'h00C; B = 16'h0081; #100;
A = 16'h00C; B = 16'h0082; #100;
A = 16'h00C; B = 16'h0083; #100;
A = 16'h00C; B = 16'h0084; #100;
A = 16'h00C; B = 16'h0085; #100;
A = 16'h00C; B = 16'h0086; #100;
A = 16'h00C; B = 16'h0087; #100;
A = 16'h00C; B = 16'h0088; #100;
A = 16'h00C; B = 16'h0089; #100;
A = 16'h00C; B = 16'h008A; #100;
A = 16'h00C; B = 16'h008B; #100;
A = 16'h00C; B = 16'h008C; #100;
A = 16'h00C; B = 16'h008D; #100;
A = 16'h00C; B = 16'h008E; #100;
A = 16'h00C; B = 16'h008F; #100;
A = 16'h00C; B = 16'h0090; #100;
A = 16'h00C; B = 16'h0091; #100;
A = 16'h00C; B = 16'h0092; #100;
A = 16'h00C; B = 16'h0093; #100;
A = 16'h00C; B = 16'h0094; #100;
A = 16'h00C; B = 16'h0095; #100;
A = 16'h00C; B = 16'h0096; #100;
A = 16'h00C; B = 16'h0097; #100;
A = 16'h00C; B = 16'h0098; #100;
A = 16'h00C; B = 16'h0099; #100;
A = 16'h00C; B = 16'h009A; #100;
A = 16'h00C; B = 16'h009B; #100;
A = 16'h00C; B = 16'h009C; #100;
A = 16'h00C; B = 16'h009D; #100;
A = 16'h00C; B = 16'h009E; #100;
A = 16'h00C; B = 16'h009F; #100;
A = 16'h00C; B = 16'h00A0; #100;
A = 16'h00C; B = 16'h00A1; #100;
A = 16'h00C; B = 16'h00A2; #100;
A = 16'h00C; B = 16'h00A3; #100;
A = 16'h00C; B = 16'h00A4; #100;
A = 16'h00C; B = 16'h00A5; #100;
A = 16'h00C; B = 16'h00A6; #100;
A = 16'h00C; B = 16'h00A7; #100;
A = 16'h00C; B = 16'h00A8; #100;
A = 16'h00C; B = 16'h00A9; #100;
A = 16'h00C; B = 16'h00AA; #100;
A = 16'h00C; B = 16'h00AB; #100;
A = 16'h00C; B = 16'h00AC; #100;
A = 16'h00C; B = 16'h00AD; #100;
A = 16'h00C; B = 16'h00AE; #100;
A = 16'h00C; B = 16'h00AF; #100;
A = 16'h00C; B = 16'h00B0; #100;
A = 16'h00C; B = 16'h00B1; #100;
A = 16'h00C; B = 16'h00B2; #100;
A = 16'h00C; B = 16'h00B3; #100;
A = 16'h00C; B = 16'h00B4; #100;
A = 16'h00C; B = 16'h00B5; #100;
A = 16'h00C; B = 16'h00B6; #100;
A = 16'h00C; B = 16'h00B7; #100;
A = 16'h00C; B = 16'h00B8; #100;
A = 16'h00C; B = 16'h00B9; #100;
A = 16'h00C; B = 16'h00BA; #100;
A = 16'h00C; B = 16'h00BB; #100;
A = 16'h00C; B = 16'h00BC; #100;
A = 16'h00C; B = 16'h00BD; #100;
A = 16'h00C; B = 16'h00BE; #100;
A = 16'h00C; B = 16'h00BF; #100;
A = 16'h00C; B = 16'h00C0; #100;
A = 16'h00C; B = 16'h00C1; #100;
A = 16'h00C; B = 16'h00C2; #100;
A = 16'h00C; B = 16'h00C3; #100;
A = 16'h00C; B = 16'h00C4; #100;
A = 16'h00C; B = 16'h00C5; #100;
A = 16'h00C; B = 16'h00C6; #100;
A = 16'h00C; B = 16'h00C7; #100;
A = 16'h00C; B = 16'h00C8; #100;
A = 16'h00C; B = 16'h00C9; #100;
A = 16'h00C; B = 16'h00CA; #100;
A = 16'h00C; B = 16'h00CB; #100;
A = 16'h00C; B = 16'h00CC; #100;
A = 16'h00C; B = 16'h00CD; #100;
A = 16'h00C; B = 16'h00CE; #100;
A = 16'h00C; B = 16'h00CF; #100;
A = 16'h00C; B = 16'h00D0; #100;
A = 16'h00C; B = 16'h00D1; #100;
A = 16'h00C; B = 16'h00D2; #100;
A = 16'h00C; B = 16'h00D3; #100;
A = 16'h00C; B = 16'h00D4; #100;
A = 16'h00C; B = 16'h00D5; #100;
A = 16'h00C; B = 16'h00D6; #100;
A = 16'h00C; B = 16'h00D7; #100;
A = 16'h00C; B = 16'h00D8; #100;
A = 16'h00C; B = 16'h00D9; #100;
A = 16'h00C; B = 16'h00DA; #100;
A = 16'h00C; B = 16'h00DB; #100;
A = 16'h00C; B = 16'h00DC; #100;
A = 16'h00C; B = 16'h00DD; #100;
A = 16'h00C; B = 16'h00DE; #100;
A = 16'h00C; B = 16'h00DF; #100;
A = 16'h00C; B = 16'h00E0; #100;
A = 16'h00C; B = 16'h00E1; #100;
A = 16'h00C; B = 16'h00E2; #100;
A = 16'h00C; B = 16'h00E3; #100;
A = 16'h00C; B = 16'h00E4; #100;
A = 16'h00C; B = 16'h00E5; #100;
A = 16'h00C; B = 16'h00E6; #100;
A = 16'h00C; B = 16'h00E7; #100;
A = 16'h00C; B = 16'h00E8; #100;
A = 16'h00C; B = 16'h00E9; #100;
A = 16'h00C; B = 16'h00EA; #100;
A = 16'h00C; B = 16'h00EB; #100;
A = 16'h00C; B = 16'h00EC; #100;
A = 16'h00C; B = 16'h00ED; #100;
A = 16'h00C; B = 16'h00EE; #100;
A = 16'h00C; B = 16'h00EF; #100;
A = 16'h00C; B = 16'h00F0; #100;
A = 16'h00C; B = 16'h00F1; #100;
A = 16'h00C; B = 16'h00F2; #100;
A = 16'h00C; B = 16'h00F3; #100;
A = 16'h00C; B = 16'h00F4; #100;
A = 16'h00C; B = 16'h00F5; #100;
A = 16'h00C; B = 16'h00F6; #100;
A = 16'h00C; B = 16'h00F7; #100;
A = 16'h00C; B = 16'h00F8; #100;
A = 16'h00C; B = 16'h00F9; #100;
A = 16'h00C; B = 16'h00FA; #100;
A = 16'h00C; B = 16'h00FB; #100;
A = 16'h00C; B = 16'h00FC; #100;
A = 16'h00C; B = 16'h00FD; #100;
A = 16'h00C; B = 16'h00FE; #100;
A = 16'h00C; B = 16'h00FF; #100;
A = 16'h00D; B = 16'h000; #100;
A = 16'h00D; B = 16'h001; #100;
A = 16'h00D; B = 16'h002; #100;
A = 16'h00D; B = 16'h003; #100;
A = 16'h00D; B = 16'h004; #100;
A = 16'h00D; B = 16'h005; #100;
A = 16'h00D; B = 16'h006; #100;
A = 16'h00D; B = 16'h007; #100;
A = 16'h00D; B = 16'h008; #100;
A = 16'h00D; B = 16'h009; #100;
A = 16'h00D; B = 16'h00A; #100;
A = 16'h00D; B = 16'h00B; #100;
A = 16'h00D; B = 16'h00C; #100;
A = 16'h00D; B = 16'h00D; #100;
A = 16'h00D; B = 16'h00E; #100;
A = 16'h00D; B = 16'h00F; #100;
A = 16'h00D; B = 16'h0010; #100;
A = 16'h00D; B = 16'h0011; #100;
A = 16'h00D; B = 16'h0012; #100;
A = 16'h00D; B = 16'h0013; #100;
A = 16'h00D; B = 16'h0014; #100;
A = 16'h00D; B = 16'h0015; #100;
A = 16'h00D; B = 16'h0016; #100;
A = 16'h00D; B = 16'h0017; #100;
A = 16'h00D; B = 16'h0018; #100;
A = 16'h00D; B = 16'h0019; #100;
A = 16'h00D; B = 16'h001A; #100;
A = 16'h00D; B = 16'h001B; #100;
A = 16'h00D; B = 16'h001C; #100;
A = 16'h00D; B = 16'h001D; #100;
A = 16'h00D; B = 16'h001E; #100;
A = 16'h00D; B = 16'h001F; #100;
A = 16'h00D; B = 16'h0020; #100;
A = 16'h00D; B = 16'h0021; #100;
A = 16'h00D; B = 16'h0022; #100;
A = 16'h00D; B = 16'h0023; #100;
A = 16'h00D; B = 16'h0024; #100;
A = 16'h00D; B = 16'h0025; #100;
A = 16'h00D; B = 16'h0026; #100;
A = 16'h00D; B = 16'h0027; #100;
A = 16'h00D; B = 16'h0028; #100;
A = 16'h00D; B = 16'h0029; #100;
A = 16'h00D; B = 16'h002A; #100;
A = 16'h00D; B = 16'h002B; #100;
A = 16'h00D; B = 16'h002C; #100;
A = 16'h00D; B = 16'h002D; #100;
A = 16'h00D; B = 16'h002E; #100;
A = 16'h00D; B = 16'h002F; #100;
A = 16'h00D; B = 16'h0030; #100;
A = 16'h00D; B = 16'h0031; #100;
A = 16'h00D; B = 16'h0032; #100;
A = 16'h00D; B = 16'h0033; #100;
A = 16'h00D; B = 16'h0034; #100;
A = 16'h00D; B = 16'h0035; #100;
A = 16'h00D; B = 16'h0036; #100;
A = 16'h00D; B = 16'h0037; #100;
A = 16'h00D; B = 16'h0038; #100;
A = 16'h00D; B = 16'h0039; #100;
A = 16'h00D; B = 16'h003A; #100;
A = 16'h00D; B = 16'h003B; #100;
A = 16'h00D; B = 16'h003C; #100;
A = 16'h00D; B = 16'h003D; #100;
A = 16'h00D; B = 16'h003E; #100;
A = 16'h00D; B = 16'h003F; #100;
A = 16'h00D; B = 16'h0040; #100;
A = 16'h00D; B = 16'h0041; #100;
A = 16'h00D; B = 16'h0042; #100;
A = 16'h00D; B = 16'h0043; #100;
A = 16'h00D; B = 16'h0044; #100;
A = 16'h00D; B = 16'h0045; #100;
A = 16'h00D; B = 16'h0046; #100;
A = 16'h00D; B = 16'h0047; #100;
A = 16'h00D; B = 16'h0048; #100;
A = 16'h00D; B = 16'h0049; #100;
A = 16'h00D; B = 16'h004A; #100;
A = 16'h00D; B = 16'h004B; #100;
A = 16'h00D; B = 16'h004C; #100;
A = 16'h00D; B = 16'h004D; #100;
A = 16'h00D; B = 16'h004E; #100;
A = 16'h00D; B = 16'h004F; #100;
A = 16'h00D; B = 16'h0050; #100;
A = 16'h00D; B = 16'h0051; #100;
A = 16'h00D; B = 16'h0052; #100;
A = 16'h00D; B = 16'h0053; #100;
A = 16'h00D; B = 16'h0054; #100;
A = 16'h00D; B = 16'h0055; #100;
A = 16'h00D; B = 16'h0056; #100;
A = 16'h00D; B = 16'h0057; #100;
A = 16'h00D; B = 16'h0058; #100;
A = 16'h00D; B = 16'h0059; #100;
A = 16'h00D; B = 16'h005A; #100;
A = 16'h00D; B = 16'h005B; #100;
A = 16'h00D; B = 16'h005C; #100;
A = 16'h00D; B = 16'h005D; #100;
A = 16'h00D; B = 16'h005E; #100;
A = 16'h00D; B = 16'h005F; #100;
A = 16'h00D; B = 16'h0060; #100;
A = 16'h00D; B = 16'h0061; #100;
A = 16'h00D; B = 16'h0062; #100;
A = 16'h00D; B = 16'h0063; #100;
A = 16'h00D; B = 16'h0064; #100;
A = 16'h00D; B = 16'h0065; #100;
A = 16'h00D; B = 16'h0066; #100;
A = 16'h00D; B = 16'h0067; #100;
A = 16'h00D; B = 16'h0068; #100;
A = 16'h00D; B = 16'h0069; #100;
A = 16'h00D; B = 16'h006A; #100;
A = 16'h00D; B = 16'h006B; #100;
A = 16'h00D; B = 16'h006C; #100;
A = 16'h00D; B = 16'h006D; #100;
A = 16'h00D; B = 16'h006E; #100;
A = 16'h00D; B = 16'h006F; #100;
A = 16'h00D; B = 16'h0070; #100;
A = 16'h00D; B = 16'h0071; #100;
A = 16'h00D; B = 16'h0072; #100;
A = 16'h00D; B = 16'h0073; #100;
A = 16'h00D; B = 16'h0074; #100;
A = 16'h00D; B = 16'h0075; #100;
A = 16'h00D; B = 16'h0076; #100;
A = 16'h00D; B = 16'h0077; #100;
A = 16'h00D; B = 16'h0078; #100;
A = 16'h00D; B = 16'h0079; #100;
A = 16'h00D; B = 16'h007A; #100;
A = 16'h00D; B = 16'h007B; #100;
A = 16'h00D; B = 16'h007C; #100;
A = 16'h00D; B = 16'h007D; #100;
A = 16'h00D; B = 16'h007E; #100;
A = 16'h00D; B = 16'h007F; #100;
A = 16'h00D; B = 16'h0080; #100;
A = 16'h00D; B = 16'h0081; #100;
A = 16'h00D; B = 16'h0082; #100;
A = 16'h00D; B = 16'h0083; #100;
A = 16'h00D; B = 16'h0084; #100;
A = 16'h00D; B = 16'h0085; #100;
A = 16'h00D; B = 16'h0086; #100;
A = 16'h00D; B = 16'h0087; #100;
A = 16'h00D; B = 16'h0088; #100;
A = 16'h00D; B = 16'h0089; #100;
A = 16'h00D; B = 16'h008A; #100;
A = 16'h00D; B = 16'h008B; #100;
A = 16'h00D; B = 16'h008C; #100;
A = 16'h00D; B = 16'h008D; #100;
A = 16'h00D; B = 16'h008E; #100;
A = 16'h00D; B = 16'h008F; #100;
A = 16'h00D; B = 16'h0090; #100;
A = 16'h00D; B = 16'h0091; #100;
A = 16'h00D; B = 16'h0092; #100;
A = 16'h00D; B = 16'h0093; #100;
A = 16'h00D; B = 16'h0094; #100;
A = 16'h00D; B = 16'h0095; #100;
A = 16'h00D; B = 16'h0096; #100;
A = 16'h00D; B = 16'h0097; #100;
A = 16'h00D; B = 16'h0098; #100;
A = 16'h00D; B = 16'h0099; #100;
A = 16'h00D; B = 16'h009A; #100;
A = 16'h00D; B = 16'h009B; #100;
A = 16'h00D; B = 16'h009C; #100;
A = 16'h00D; B = 16'h009D; #100;
A = 16'h00D; B = 16'h009E; #100;
A = 16'h00D; B = 16'h009F; #100;
A = 16'h00D; B = 16'h00A0; #100;
A = 16'h00D; B = 16'h00A1; #100;
A = 16'h00D; B = 16'h00A2; #100;
A = 16'h00D; B = 16'h00A3; #100;
A = 16'h00D; B = 16'h00A4; #100;
A = 16'h00D; B = 16'h00A5; #100;
A = 16'h00D; B = 16'h00A6; #100;
A = 16'h00D; B = 16'h00A7; #100;
A = 16'h00D; B = 16'h00A8; #100;
A = 16'h00D; B = 16'h00A9; #100;
A = 16'h00D; B = 16'h00AA; #100;
A = 16'h00D; B = 16'h00AB; #100;
A = 16'h00D; B = 16'h00AC; #100;
A = 16'h00D; B = 16'h00AD; #100;
A = 16'h00D; B = 16'h00AE; #100;
A = 16'h00D; B = 16'h00AF; #100;
A = 16'h00D; B = 16'h00B0; #100;
A = 16'h00D; B = 16'h00B1; #100;
A = 16'h00D; B = 16'h00B2; #100;
A = 16'h00D; B = 16'h00B3; #100;
A = 16'h00D; B = 16'h00B4; #100;
A = 16'h00D; B = 16'h00B5; #100;
A = 16'h00D; B = 16'h00B6; #100;
A = 16'h00D; B = 16'h00B7; #100;
A = 16'h00D; B = 16'h00B8; #100;
A = 16'h00D; B = 16'h00B9; #100;
A = 16'h00D; B = 16'h00BA; #100;
A = 16'h00D; B = 16'h00BB; #100;
A = 16'h00D; B = 16'h00BC; #100;
A = 16'h00D; B = 16'h00BD; #100;
A = 16'h00D; B = 16'h00BE; #100;
A = 16'h00D; B = 16'h00BF; #100;
A = 16'h00D; B = 16'h00C0; #100;
A = 16'h00D; B = 16'h00C1; #100;
A = 16'h00D; B = 16'h00C2; #100;
A = 16'h00D; B = 16'h00C3; #100;
A = 16'h00D; B = 16'h00C4; #100;
A = 16'h00D; B = 16'h00C5; #100;
A = 16'h00D; B = 16'h00C6; #100;
A = 16'h00D; B = 16'h00C7; #100;
A = 16'h00D; B = 16'h00C8; #100;
A = 16'h00D; B = 16'h00C9; #100;
A = 16'h00D; B = 16'h00CA; #100;
A = 16'h00D; B = 16'h00CB; #100;
A = 16'h00D; B = 16'h00CC; #100;
A = 16'h00D; B = 16'h00CD; #100;
A = 16'h00D; B = 16'h00CE; #100;
A = 16'h00D; B = 16'h00CF; #100;
A = 16'h00D; B = 16'h00D0; #100;
A = 16'h00D; B = 16'h00D1; #100;
A = 16'h00D; B = 16'h00D2; #100;
A = 16'h00D; B = 16'h00D3; #100;
A = 16'h00D; B = 16'h00D4; #100;
A = 16'h00D; B = 16'h00D5; #100;
A = 16'h00D; B = 16'h00D6; #100;
A = 16'h00D; B = 16'h00D7; #100;
A = 16'h00D; B = 16'h00D8; #100;
A = 16'h00D; B = 16'h00D9; #100;
A = 16'h00D; B = 16'h00DA; #100;
A = 16'h00D; B = 16'h00DB; #100;
A = 16'h00D; B = 16'h00DC; #100;
A = 16'h00D; B = 16'h00DD; #100;
A = 16'h00D; B = 16'h00DE; #100;
A = 16'h00D; B = 16'h00DF; #100;
A = 16'h00D; B = 16'h00E0; #100;
A = 16'h00D; B = 16'h00E1; #100;
A = 16'h00D; B = 16'h00E2; #100;
A = 16'h00D; B = 16'h00E3; #100;
A = 16'h00D; B = 16'h00E4; #100;
A = 16'h00D; B = 16'h00E5; #100;
A = 16'h00D; B = 16'h00E6; #100;
A = 16'h00D; B = 16'h00E7; #100;
A = 16'h00D; B = 16'h00E8; #100;
A = 16'h00D; B = 16'h00E9; #100;
A = 16'h00D; B = 16'h00EA; #100;
A = 16'h00D; B = 16'h00EB; #100;
A = 16'h00D; B = 16'h00EC; #100;
A = 16'h00D; B = 16'h00ED; #100;
A = 16'h00D; B = 16'h00EE; #100;
A = 16'h00D; B = 16'h00EF; #100;
A = 16'h00D; B = 16'h00F0; #100;
A = 16'h00D; B = 16'h00F1; #100;
A = 16'h00D; B = 16'h00F2; #100;
A = 16'h00D; B = 16'h00F3; #100;
A = 16'h00D; B = 16'h00F4; #100;
A = 16'h00D; B = 16'h00F5; #100;
A = 16'h00D; B = 16'h00F6; #100;
A = 16'h00D; B = 16'h00F7; #100;
A = 16'h00D; B = 16'h00F8; #100;
A = 16'h00D; B = 16'h00F9; #100;
A = 16'h00D; B = 16'h00FA; #100;
A = 16'h00D; B = 16'h00FB; #100;
A = 16'h00D; B = 16'h00FC; #100;
A = 16'h00D; B = 16'h00FD; #100;
A = 16'h00D; B = 16'h00FE; #100;
A = 16'h00D; B = 16'h00FF; #100;
A = 16'h00E; B = 16'h000; #100;
A = 16'h00E; B = 16'h001; #100;
A = 16'h00E; B = 16'h002; #100;
A = 16'h00E; B = 16'h003; #100;
A = 16'h00E; B = 16'h004; #100;
A = 16'h00E; B = 16'h005; #100;
A = 16'h00E; B = 16'h006; #100;
A = 16'h00E; B = 16'h007; #100;
A = 16'h00E; B = 16'h008; #100;
A = 16'h00E; B = 16'h009; #100;
A = 16'h00E; B = 16'h00A; #100;
A = 16'h00E; B = 16'h00B; #100;
A = 16'h00E; B = 16'h00C; #100;
A = 16'h00E; B = 16'h00D; #100;
A = 16'h00E; B = 16'h00E; #100;
A = 16'h00E; B = 16'h00F; #100;
A = 16'h00E; B = 16'h0010; #100;
A = 16'h00E; B = 16'h0011; #100;
A = 16'h00E; B = 16'h0012; #100;
A = 16'h00E; B = 16'h0013; #100;
A = 16'h00E; B = 16'h0014; #100;
A = 16'h00E; B = 16'h0015; #100;
A = 16'h00E; B = 16'h0016; #100;
A = 16'h00E; B = 16'h0017; #100;
A = 16'h00E; B = 16'h0018; #100;
A = 16'h00E; B = 16'h0019; #100;
A = 16'h00E; B = 16'h001A; #100;
A = 16'h00E; B = 16'h001B; #100;
A = 16'h00E; B = 16'h001C; #100;
A = 16'h00E; B = 16'h001D; #100;
A = 16'h00E; B = 16'h001E; #100;
A = 16'h00E; B = 16'h001F; #100;
A = 16'h00E; B = 16'h0020; #100;
A = 16'h00E; B = 16'h0021; #100;
A = 16'h00E; B = 16'h0022; #100;
A = 16'h00E; B = 16'h0023; #100;
A = 16'h00E; B = 16'h0024; #100;
A = 16'h00E; B = 16'h0025; #100;
A = 16'h00E; B = 16'h0026; #100;
A = 16'h00E; B = 16'h0027; #100;
A = 16'h00E; B = 16'h0028; #100;
A = 16'h00E; B = 16'h0029; #100;
A = 16'h00E; B = 16'h002A; #100;
A = 16'h00E; B = 16'h002B; #100;
A = 16'h00E; B = 16'h002C; #100;
A = 16'h00E; B = 16'h002D; #100;
A = 16'h00E; B = 16'h002E; #100;
A = 16'h00E; B = 16'h002F; #100;
A = 16'h00E; B = 16'h0030; #100;
A = 16'h00E; B = 16'h0031; #100;
A = 16'h00E; B = 16'h0032; #100;
A = 16'h00E; B = 16'h0033; #100;
A = 16'h00E; B = 16'h0034; #100;
A = 16'h00E; B = 16'h0035; #100;
A = 16'h00E; B = 16'h0036; #100;
A = 16'h00E; B = 16'h0037; #100;
A = 16'h00E; B = 16'h0038; #100;
A = 16'h00E; B = 16'h0039; #100;
A = 16'h00E; B = 16'h003A; #100;
A = 16'h00E; B = 16'h003B; #100;
A = 16'h00E; B = 16'h003C; #100;
A = 16'h00E; B = 16'h003D; #100;
A = 16'h00E; B = 16'h003E; #100;
A = 16'h00E; B = 16'h003F; #100;
A = 16'h00E; B = 16'h0040; #100;
A = 16'h00E; B = 16'h0041; #100;
A = 16'h00E; B = 16'h0042; #100;
A = 16'h00E; B = 16'h0043; #100;
A = 16'h00E; B = 16'h0044; #100;
A = 16'h00E; B = 16'h0045; #100;
A = 16'h00E; B = 16'h0046; #100;
A = 16'h00E; B = 16'h0047; #100;
A = 16'h00E; B = 16'h0048; #100;
A = 16'h00E; B = 16'h0049; #100;
A = 16'h00E; B = 16'h004A; #100;
A = 16'h00E; B = 16'h004B; #100;
A = 16'h00E; B = 16'h004C; #100;
A = 16'h00E; B = 16'h004D; #100;
A = 16'h00E; B = 16'h004E; #100;
A = 16'h00E; B = 16'h004F; #100;
A = 16'h00E; B = 16'h0050; #100;
A = 16'h00E; B = 16'h0051; #100;
A = 16'h00E; B = 16'h0052; #100;
A = 16'h00E; B = 16'h0053; #100;
A = 16'h00E; B = 16'h0054; #100;
A = 16'h00E; B = 16'h0055; #100;
A = 16'h00E; B = 16'h0056; #100;
A = 16'h00E; B = 16'h0057; #100;
A = 16'h00E; B = 16'h0058; #100;
A = 16'h00E; B = 16'h0059; #100;
A = 16'h00E; B = 16'h005A; #100;
A = 16'h00E; B = 16'h005B; #100;
A = 16'h00E; B = 16'h005C; #100;
A = 16'h00E; B = 16'h005D; #100;
A = 16'h00E; B = 16'h005E; #100;
A = 16'h00E; B = 16'h005F; #100;
A = 16'h00E; B = 16'h0060; #100;
A = 16'h00E; B = 16'h0061; #100;
A = 16'h00E; B = 16'h0062; #100;
A = 16'h00E; B = 16'h0063; #100;
A = 16'h00E; B = 16'h0064; #100;
A = 16'h00E; B = 16'h0065; #100;
A = 16'h00E; B = 16'h0066; #100;
A = 16'h00E; B = 16'h0067; #100;
A = 16'h00E; B = 16'h0068; #100;
A = 16'h00E; B = 16'h0069; #100;
A = 16'h00E; B = 16'h006A; #100;
A = 16'h00E; B = 16'h006B; #100;
A = 16'h00E; B = 16'h006C; #100;
A = 16'h00E; B = 16'h006D; #100;
A = 16'h00E; B = 16'h006E; #100;
A = 16'h00E; B = 16'h006F; #100;
A = 16'h00E; B = 16'h0070; #100;
A = 16'h00E; B = 16'h0071; #100;
A = 16'h00E; B = 16'h0072; #100;
A = 16'h00E; B = 16'h0073; #100;
A = 16'h00E; B = 16'h0074; #100;
A = 16'h00E; B = 16'h0075; #100;
A = 16'h00E; B = 16'h0076; #100;
A = 16'h00E; B = 16'h0077; #100;
A = 16'h00E; B = 16'h0078; #100;
A = 16'h00E; B = 16'h0079; #100;
A = 16'h00E; B = 16'h007A; #100;
A = 16'h00E; B = 16'h007B; #100;
A = 16'h00E; B = 16'h007C; #100;
A = 16'h00E; B = 16'h007D; #100;
A = 16'h00E; B = 16'h007E; #100;
A = 16'h00E; B = 16'h007F; #100;
A = 16'h00E; B = 16'h0080; #100;
A = 16'h00E; B = 16'h0081; #100;
A = 16'h00E; B = 16'h0082; #100;
A = 16'h00E; B = 16'h0083; #100;
A = 16'h00E; B = 16'h0084; #100;
A = 16'h00E; B = 16'h0085; #100;
A = 16'h00E; B = 16'h0086; #100;
A = 16'h00E; B = 16'h0087; #100;
A = 16'h00E; B = 16'h0088; #100;
A = 16'h00E; B = 16'h0089; #100;
A = 16'h00E; B = 16'h008A; #100;
A = 16'h00E; B = 16'h008B; #100;
A = 16'h00E; B = 16'h008C; #100;
A = 16'h00E; B = 16'h008D; #100;
A = 16'h00E; B = 16'h008E; #100;
A = 16'h00E; B = 16'h008F; #100;
A = 16'h00E; B = 16'h0090; #100;
A = 16'h00E; B = 16'h0091; #100;
A = 16'h00E; B = 16'h0092; #100;
A = 16'h00E; B = 16'h0093; #100;
A = 16'h00E; B = 16'h0094; #100;
A = 16'h00E; B = 16'h0095; #100;
A = 16'h00E; B = 16'h0096; #100;
A = 16'h00E; B = 16'h0097; #100;
A = 16'h00E; B = 16'h0098; #100;
A = 16'h00E; B = 16'h0099; #100;
A = 16'h00E; B = 16'h009A; #100;
A = 16'h00E; B = 16'h009B; #100;
A = 16'h00E; B = 16'h009C; #100;
A = 16'h00E; B = 16'h009D; #100;
A = 16'h00E; B = 16'h009E; #100;
A = 16'h00E; B = 16'h009F; #100;
A = 16'h00E; B = 16'h00A0; #100;
A = 16'h00E; B = 16'h00A1; #100;
A = 16'h00E; B = 16'h00A2; #100;
A = 16'h00E; B = 16'h00A3; #100;
A = 16'h00E; B = 16'h00A4; #100;
A = 16'h00E; B = 16'h00A5; #100;
A = 16'h00E; B = 16'h00A6; #100;
A = 16'h00E; B = 16'h00A7; #100;
A = 16'h00E; B = 16'h00A8; #100;
A = 16'h00E; B = 16'h00A9; #100;
A = 16'h00E; B = 16'h00AA; #100;
A = 16'h00E; B = 16'h00AB; #100;
A = 16'h00E; B = 16'h00AC; #100;
A = 16'h00E; B = 16'h00AD; #100;
A = 16'h00E; B = 16'h00AE; #100;
A = 16'h00E; B = 16'h00AF; #100;
A = 16'h00E; B = 16'h00B0; #100;
A = 16'h00E; B = 16'h00B1; #100;
A = 16'h00E; B = 16'h00B2; #100;
A = 16'h00E; B = 16'h00B3; #100;
A = 16'h00E; B = 16'h00B4; #100;
A = 16'h00E; B = 16'h00B5; #100;
A = 16'h00E; B = 16'h00B6; #100;
A = 16'h00E; B = 16'h00B7; #100;
A = 16'h00E; B = 16'h00B8; #100;
A = 16'h00E; B = 16'h00B9; #100;
A = 16'h00E; B = 16'h00BA; #100;
A = 16'h00E; B = 16'h00BB; #100;
A = 16'h00E; B = 16'h00BC; #100;
A = 16'h00E; B = 16'h00BD; #100;
A = 16'h00E; B = 16'h00BE; #100;
A = 16'h00E; B = 16'h00BF; #100;
A = 16'h00E; B = 16'h00C0; #100;
A = 16'h00E; B = 16'h00C1; #100;
A = 16'h00E; B = 16'h00C2; #100;
A = 16'h00E; B = 16'h00C3; #100;
A = 16'h00E; B = 16'h00C4; #100;
A = 16'h00E; B = 16'h00C5; #100;
A = 16'h00E; B = 16'h00C6; #100;
A = 16'h00E; B = 16'h00C7; #100;
A = 16'h00E; B = 16'h00C8; #100;
A = 16'h00E; B = 16'h00C9; #100;
A = 16'h00E; B = 16'h00CA; #100;
A = 16'h00E; B = 16'h00CB; #100;
A = 16'h00E; B = 16'h00CC; #100;
A = 16'h00E; B = 16'h00CD; #100;
A = 16'h00E; B = 16'h00CE; #100;
A = 16'h00E; B = 16'h00CF; #100;
A = 16'h00E; B = 16'h00D0; #100;
A = 16'h00E; B = 16'h00D1; #100;
A = 16'h00E; B = 16'h00D2; #100;
A = 16'h00E; B = 16'h00D3; #100;
A = 16'h00E; B = 16'h00D4; #100;
A = 16'h00E; B = 16'h00D5; #100;
A = 16'h00E; B = 16'h00D6; #100;
A = 16'h00E; B = 16'h00D7; #100;
A = 16'h00E; B = 16'h00D8; #100;
A = 16'h00E; B = 16'h00D9; #100;
A = 16'h00E; B = 16'h00DA; #100;
A = 16'h00E; B = 16'h00DB; #100;
A = 16'h00E; B = 16'h00DC; #100;
A = 16'h00E; B = 16'h00DD; #100;
A = 16'h00E; B = 16'h00DE; #100;
A = 16'h00E; B = 16'h00DF; #100;
A = 16'h00E; B = 16'h00E0; #100;
A = 16'h00E; B = 16'h00E1; #100;
A = 16'h00E; B = 16'h00E2; #100;
A = 16'h00E; B = 16'h00E3; #100;
A = 16'h00E; B = 16'h00E4; #100;
A = 16'h00E; B = 16'h00E5; #100;
A = 16'h00E; B = 16'h00E6; #100;
A = 16'h00E; B = 16'h00E7; #100;
A = 16'h00E; B = 16'h00E8; #100;
A = 16'h00E; B = 16'h00E9; #100;
A = 16'h00E; B = 16'h00EA; #100;
A = 16'h00E; B = 16'h00EB; #100;
A = 16'h00E; B = 16'h00EC; #100;
A = 16'h00E; B = 16'h00ED; #100;
A = 16'h00E; B = 16'h00EE; #100;
A = 16'h00E; B = 16'h00EF; #100;
A = 16'h00E; B = 16'h00F0; #100;
A = 16'h00E; B = 16'h00F1; #100;
A = 16'h00E; B = 16'h00F2; #100;
A = 16'h00E; B = 16'h00F3; #100;
A = 16'h00E; B = 16'h00F4; #100;
A = 16'h00E; B = 16'h00F5; #100;
A = 16'h00E; B = 16'h00F6; #100;
A = 16'h00E; B = 16'h00F7; #100;
A = 16'h00E; B = 16'h00F8; #100;
A = 16'h00E; B = 16'h00F9; #100;
A = 16'h00E; B = 16'h00FA; #100;
A = 16'h00E; B = 16'h00FB; #100;
A = 16'h00E; B = 16'h00FC; #100;
A = 16'h00E; B = 16'h00FD; #100;
A = 16'h00E; B = 16'h00FE; #100;
A = 16'h00E; B = 16'h00FF; #100;
A = 16'h00F; B = 16'h000; #100;
A = 16'h00F; B = 16'h001; #100;
A = 16'h00F; B = 16'h002; #100;
A = 16'h00F; B = 16'h003; #100;
A = 16'h00F; B = 16'h004; #100;
A = 16'h00F; B = 16'h005; #100;
A = 16'h00F; B = 16'h006; #100;
A = 16'h00F; B = 16'h007; #100;
A = 16'h00F; B = 16'h008; #100;
A = 16'h00F; B = 16'h009; #100;
A = 16'h00F; B = 16'h00A; #100;
A = 16'h00F; B = 16'h00B; #100;
A = 16'h00F; B = 16'h00C; #100;
A = 16'h00F; B = 16'h00D; #100;
A = 16'h00F; B = 16'h00E; #100;
A = 16'h00F; B = 16'h00F; #100;
A = 16'h00F; B = 16'h0010; #100;
A = 16'h00F; B = 16'h0011; #100;
A = 16'h00F; B = 16'h0012; #100;
A = 16'h00F; B = 16'h0013; #100;
A = 16'h00F; B = 16'h0014; #100;
A = 16'h00F; B = 16'h0015; #100;
A = 16'h00F; B = 16'h0016; #100;
A = 16'h00F; B = 16'h0017; #100;
A = 16'h00F; B = 16'h0018; #100;
A = 16'h00F; B = 16'h0019; #100;
A = 16'h00F; B = 16'h001A; #100;
A = 16'h00F; B = 16'h001B; #100;
A = 16'h00F; B = 16'h001C; #100;
A = 16'h00F; B = 16'h001D; #100;
A = 16'h00F; B = 16'h001E; #100;
A = 16'h00F; B = 16'h001F; #100;
A = 16'h00F; B = 16'h0020; #100;
A = 16'h00F; B = 16'h0021; #100;
A = 16'h00F; B = 16'h0022; #100;
A = 16'h00F; B = 16'h0023; #100;
A = 16'h00F; B = 16'h0024; #100;
A = 16'h00F; B = 16'h0025; #100;
A = 16'h00F; B = 16'h0026; #100;
A = 16'h00F; B = 16'h0027; #100;
A = 16'h00F; B = 16'h0028; #100;
A = 16'h00F; B = 16'h0029; #100;
A = 16'h00F; B = 16'h002A; #100;
A = 16'h00F; B = 16'h002B; #100;
A = 16'h00F; B = 16'h002C; #100;
A = 16'h00F; B = 16'h002D; #100;
A = 16'h00F; B = 16'h002E; #100;
A = 16'h00F; B = 16'h002F; #100;
A = 16'h00F; B = 16'h0030; #100;
A = 16'h00F; B = 16'h0031; #100;
A = 16'h00F; B = 16'h0032; #100;
A = 16'h00F; B = 16'h0033; #100;
A = 16'h00F; B = 16'h0034; #100;
A = 16'h00F; B = 16'h0035; #100;
A = 16'h00F; B = 16'h0036; #100;
A = 16'h00F; B = 16'h0037; #100;
A = 16'h00F; B = 16'h0038; #100;
A = 16'h00F; B = 16'h0039; #100;
A = 16'h00F; B = 16'h003A; #100;
A = 16'h00F; B = 16'h003B; #100;
A = 16'h00F; B = 16'h003C; #100;
A = 16'h00F; B = 16'h003D; #100;
A = 16'h00F; B = 16'h003E; #100;
A = 16'h00F; B = 16'h003F; #100;
A = 16'h00F; B = 16'h0040; #100;
A = 16'h00F; B = 16'h0041; #100;
A = 16'h00F; B = 16'h0042; #100;
A = 16'h00F; B = 16'h0043; #100;
A = 16'h00F; B = 16'h0044; #100;
A = 16'h00F; B = 16'h0045; #100;
A = 16'h00F; B = 16'h0046; #100;
A = 16'h00F; B = 16'h0047; #100;
A = 16'h00F; B = 16'h0048; #100;
A = 16'h00F; B = 16'h0049; #100;
A = 16'h00F; B = 16'h004A; #100;
A = 16'h00F; B = 16'h004B; #100;
A = 16'h00F; B = 16'h004C; #100;
A = 16'h00F; B = 16'h004D; #100;
A = 16'h00F; B = 16'h004E; #100;
A = 16'h00F; B = 16'h004F; #100;
A = 16'h00F; B = 16'h0050; #100;
A = 16'h00F; B = 16'h0051; #100;
A = 16'h00F; B = 16'h0052; #100;
A = 16'h00F; B = 16'h0053; #100;
A = 16'h00F; B = 16'h0054; #100;
A = 16'h00F; B = 16'h0055; #100;
A = 16'h00F; B = 16'h0056; #100;
A = 16'h00F; B = 16'h0057; #100;
A = 16'h00F; B = 16'h0058; #100;
A = 16'h00F; B = 16'h0059; #100;
A = 16'h00F; B = 16'h005A; #100;
A = 16'h00F; B = 16'h005B; #100;
A = 16'h00F; B = 16'h005C; #100;
A = 16'h00F; B = 16'h005D; #100;
A = 16'h00F; B = 16'h005E; #100;
A = 16'h00F; B = 16'h005F; #100;
A = 16'h00F; B = 16'h0060; #100;
A = 16'h00F; B = 16'h0061; #100;
A = 16'h00F; B = 16'h0062; #100;
A = 16'h00F; B = 16'h0063; #100;
A = 16'h00F; B = 16'h0064; #100;
A = 16'h00F; B = 16'h0065; #100;
A = 16'h00F; B = 16'h0066; #100;
A = 16'h00F; B = 16'h0067; #100;
A = 16'h00F; B = 16'h0068; #100;
A = 16'h00F; B = 16'h0069; #100;
A = 16'h00F; B = 16'h006A; #100;
A = 16'h00F; B = 16'h006B; #100;
A = 16'h00F; B = 16'h006C; #100;
A = 16'h00F; B = 16'h006D; #100;
A = 16'h00F; B = 16'h006E; #100;
A = 16'h00F; B = 16'h006F; #100;
A = 16'h00F; B = 16'h0070; #100;
A = 16'h00F; B = 16'h0071; #100;
A = 16'h00F; B = 16'h0072; #100;
A = 16'h00F; B = 16'h0073; #100;
A = 16'h00F; B = 16'h0074; #100;
A = 16'h00F; B = 16'h0075; #100;
A = 16'h00F; B = 16'h0076; #100;
A = 16'h00F; B = 16'h0077; #100;
A = 16'h00F; B = 16'h0078; #100;
A = 16'h00F; B = 16'h0079; #100;
A = 16'h00F; B = 16'h007A; #100;
A = 16'h00F; B = 16'h007B; #100;
A = 16'h00F; B = 16'h007C; #100;
A = 16'h00F; B = 16'h007D; #100;
A = 16'h00F; B = 16'h007E; #100;
A = 16'h00F; B = 16'h007F; #100;
A = 16'h00F; B = 16'h0080; #100;
A = 16'h00F; B = 16'h0081; #100;
A = 16'h00F; B = 16'h0082; #100;
A = 16'h00F; B = 16'h0083; #100;
A = 16'h00F; B = 16'h0084; #100;
A = 16'h00F; B = 16'h0085; #100;
A = 16'h00F; B = 16'h0086; #100;
A = 16'h00F; B = 16'h0087; #100;
A = 16'h00F; B = 16'h0088; #100;
A = 16'h00F; B = 16'h0089; #100;
A = 16'h00F; B = 16'h008A; #100;
A = 16'h00F; B = 16'h008B; #100;
A = 16'h00F; B = 16'h008C; #100;
A = 16'h00F; B = 16'h008D; #100;
A = 16'h00F; B = 16'h008E; #100;
A = 16'h00F; B = 16'h008F; #100;
A = 16'h00F; B = 16'h0090; #100;
A = 16'h00F; B = 16'h0091; #100;
A = 16'h00F; B = 16'h0092; #100;
A = 16'h00F; B = 16'h0093; #100;
A = 16'h00F; B = 16'h0094; #100;
A = 16'h00F; B = 16'h0095; #100;
A = 16'h00F; B = 16'h0096; #100;
A = 16'h00F; B = 16'h0097; #100;
A = 16'h00F; B = 16'h0098; #100;
A = 16'h00F; B = 16'h0099; #100;
A = 16'h00F; B = 16'h009A; #100;
A = 16'h00F; B = 16'h009B; #100;
A = 16'h00F; B = 16'h009C; #100;
A = 16'h00F; B = 16'h009D; #100;
A = 16'h00F; B = 16'h009E; #100;
A = 16'h00F; B = 16'h009F; #100;
A = 16'h00F; B = 16'h00A0; #100;
A = 16'h00F; B = 16'h00A1; #100;
A = 16'h00F; B = 16'h00A2; #100;
A = 16'h00F; B = 16'h00A3; #100;
A = 16'h00F; B = 16'h00A4; #100;
A = 16'h00F; B = 16'h00A5; #100;
A = 16'h00F; B = 16'h00A6; #100;
A = 16'h00F; B = 16'h00A7; #100;
A = 16'h00F; B = 16'h00A8; #100;
A = 16'h00F; B = 16'h00A9; #100;
A = 16'h00F; B = 16'h00AA; #100;
A = 16'h00F; B = 16'h00AB; #100;
A = 16'h00F; B = 16'h00AC; #100;
A = 16'h00F; B = 16'h00AD; #100;
A = 16'h00F; B = 16'h00AE; #100;
A = 16'h00F; B = 16'h00AF; #100;
A = 16'h00F; B = 16'h00B0; #100;
A = 16'h00F; B = 16'h00B1; #100;
A = 16'h00F; B = 16'h00B2; #100;
A = 16'h00F; B = 16'h00B3; #100;
A = 16'h00F; B = 16'h00B4; #100;
A = 16'h00F; B = 16'h00B5; #100;
A = 16'h00F; B = 16'h00B6; #100;
A = 16'h00F; B = 16'h00B7; #100;
A = 16'h00F; B = 16'h00B8; #100;
A = 16'h00F; B = 16'h00B9; #100;
A = 16'h00F; B = 16'h00BA; #100;
A = 16'h00F; B = 16'h00BB; #100;
A = 16'h00F; B = 16'h00BC; #100;
A = 16'h00F; B = 16'h00BD; #100;
A = 16'h00F; B = 16'h00BE; #100;
A = 16'h00F; B = 16'h00BF; #100;
A = 16'h00F; B = 16'h00C0; #100;
A = 16'h00F; B = 16'h00C1; #100;
A = 16'h00F; B = 16'h00C2; #100;
A = 16'h00F; B = 16'h00C3; #100;
A = 16'h00F; B = 16'h00C4; #100;
A = 16'h00F; B = 16'h00C5; #100;
A = 16'h00F; B = 16'h00C6; #100;
A = 16'h00F; B = 16'h00C7; #100;
A = 16'h00F; B = 16'h00C8; #100;
A = 16'h00F; B = 16'h00C9; #100;
A = 16'h00F; B = 16'h00CA; #100;
A = 16'h00F; B = 16'h00CB; #100;
A = 16'h00F; B = 16'h00CC; #100;
A = 16'h00F; B = 16'h00CD; #100;
A = 16'h00F; B = 16'h00CE; #100;
A = 16'h00F; B = 16'h00CF; #100;
A = 16'h00F; B = 16'h00D0; #100;
A = 16'h00F; B = 16'h00D1; #100;
A = 16'h00F; B = 16'h00D2; #100;
A = 16'h00F; B = 16'h00D3; #100;
A = 16'h00F; B = 16'h00D4; #100;
A = 16'h00F; B = 16'h00D5; #100;
A = 16'h00F; B = 16'h00D6; #100;
A = 16'h00F; B = 16'h00D7; #100;
A = 16'h00F; B = 16'h00D8; #100;
A = 16'h00F; B = 16'h00D9; #100;
A = 16'h00F; B = 16'h00DA; #100;
A = 16'h00F; B = 16'h00DB; #100;
A = 16'h00F; B = 16'h00DC; #100;
A = 16'h00F; B = 16'h00DD; #100;
A = 16'h00F; B = 16'h00DE; #100;
A = 16'h00F; B = 16'h00DF; #100;
A = 16'h00F; B = 16'h00E0; #100;
A = 16'h00F; B = 16'h00E1; #100;
A = 16'h00F; B = 16'h00E2; #100;
A = 16'h00F; B = 16'h00E3; #100;
A = 16'h00F; B = 16'h00E4; #100;
A = 16'h00F; B = 16'h00E5; #100;
A = 16'h00F; B = 16'h00E6; #100;
A = 16'h00F; B = 16'h00E7; #100;
A = 16'h00F; B = 16'h00E8; #100;
A = 16'h00F; B = 16'h00E9; #100;
A = 16'h00F; B = 16'h00EA; #100;
A = 16'h00F; B = 16'h00EB; #100;
A = 16'h00F; B = 16'h00EC; #100;
A = 16'h00F; B = 16'h00ED; #100;
A = 16'h00F; B = 16'h00EE; #100;
A = 16'h00F; B = 16'h00EF; #100;
A = 16'h00F; B = 16'h00F0; #100;
A = 16'h00F; B = 16'h00F1; #100;
A = 16'h00F; B = 16'h00F2; #100;
A = 16'h00F; B = 16'h00F3; #100;
A = 16'h00F; B = 16'h00F4; #100;
A = 16'h00F; B = 16'h00F5; #100;
A = 16'h00F; B = 16'h00F6; #100;
A = 16'h00F; B = 16'h00F7; #100;
A = 16'h00F; B = 16'h00F8; #100;
A = 16'h00F; B = 16'h00F9; #100;
A = 16'h00F; B = 16'h00FA; #100;
A = 16'h00F; B = 16'h00FB; #100;
A = 16'h00F; B = 16'h00FC; #100;
A = 16'h00F; B = 16'h00FD; #100;
A = 16'h00F; B = 16'h00FE; #100;
A = 16'h00F; B = 16'h00FF; #100;
A = 16'h0010; B = 16'h000; #100;
A = 16'h0010; B = 16'h001; #100;
A = 16'h0010; B = 16'h002; #100;
A = 16'h0010; B = 16'h003; #100;
A = 16'h0010; B = 16'h004; #100;
A = 16'h0010; B = 16'h005; #100;
A = 16'h0010; B = 16'h006; #100;
A = 16'h0010; B = 16'h007; #100;
A = 16'h0010; B = 16'h008; #100;
A = 16'h0010; B = 16'h009; #100;
A = 16'h0010; B = 16'h00A; #100;
A = 16'h0010; B = 16'h00B; #100;
A = 16'h0010; B = 16'h00C; #100;
A = 16'h0010; B = 16'h00D; #100;
A = 16'h0010; B = 16'h00E; #100;
A = 16'h0010; B = 16'h00F; #100;
A = 16'h0010; B = 16'h0010; #100;
A = 16'h0010; B = 16'h0011; #100;
A = 16'h0010; B = 16'h0012; #100;
A = 16'h0010; B = 16'h0013; #100;
A = 16'h0010; B = 16'h0014; #100;
A = 16'h0010; B = 16'h0015; #100;
A = 16'h0010; B = 16'h0016; #100;
A = 16'h0010; B = 16'h0017; #100;
A = 16'h0010; B = 16'h0018; #100;
A = 16'h0010; B = 16'h0019; #100;
A = 16'h0010; B = 16'h001A; #100;
A = 16'h0010; B = 16'h001B; #100;
A = 16'h0010; B = 16'h001C; #100;
A = 16'h0010; B = 16'h001D; #100;
A = 16'h0010; B = 16'h001E; #100;
A = 16'h0010; B = 16'h001F; #100;
A = 16'h0010; B = 16'h0020; #100;
A = 16'h0010; B = 16'h0021; #100;
A = 16'h0010; B = 16'h0022; #100;
A = 16'h0010; B = 16'h0023; #100;
A = 16'h0010; B = 16'h0024; #100;
A = 16'h0010; B = 16'h0025; #100;
A = 16'h0010; B = 16'h0026; #100;
A = 16'h0010; B = 16'h0027; #100;
A = 16'h0010; B = 16'h0028; #100;
A = 16'h0010; B = 16'h0029; #100;
A = 16'h0010; B = 16'h002A; #100;
A = 16'h0010; B = 16'h002B; #100;
A = 16'h0010; B = 16'h002C; #100;
A = 16'h0010; B = 16'h002D; #100;
A = 16'h0010; B = 16'h002E; #100;
A = 16'h0010; B = 16'h002F; #100;
A = 16'h0010; B = 16'h0030; #100;
A = 16'h0010; B = 16'h0031; #100;
A = 16'h0010; B = 16'h0032; #100;
A = 16'h0010; B = 16'h0033; #100;
A = 16'h0010; B = 16'h0034; #100;
A = 16'h0010; B = 16'h0035; #100;
A = 16'h0010; B = 16'h0036; #100;
A = 16'h0010; B = 16'h0037; #100;
A = 16'h0010; B = 16'h0038; #100;
A = 16'h0010; B = 16'h0039; #100;
A = 16'h0010; B = 16'h003A; #100;
A = 16'h0010; B = 16'h003B; #100;
A = 16'h0010; B = 16'h003C; #100;
A = 16'h0010; B = 16'h003D; #100;
A = 16'h0010; B = 16'h003E; #100;
A = 16'h0010; B = 16'h003F; #100;
A = 16'h0010; B = 16'h0040; #100;
A = 16'h0010; B = 16'h0041; #100;
A = 16'h0010; B = 16'h0042; #100;
A = 16'h0010; B = 16'h0043; #100;
A = 16'h0010; B = 16'h0044; #100;
A = 16'h0010; B = 16'h0045; #100;
A = 16'h0010; B = 16'h0046; #100;
A = 16'h0010; B = 16'h0047; #100;
A = 16'h0010; B = 16'h0048; #100;
A = 16'h0010; B = 16'h0049; #100;
A = 16'h0010; B = 16'h004A; #100;
A = 16'h0010; B = 16'h004B; #100;
A = 16'h0010; B = 16'h004C; #100;
A = 16'h0010; B = 16'h004D; #100;
A = 16'h0010; B = 16'h004E; #100;
A = 16'h0010; B = 16'h004F; #100;
A = 16'h0010; B = 16'h0050; #100;
A = 16'h0010; B = 16'h0051; #100;
A = 16'h0010; B = 16'h0052; #100;
A = 16'h0010; B = 16'h0053; #100;
A = 16'h0010; B = 16'h0054; #100;
A = 16'h0010; B = 16'h0055; #100;
A = 16'h0010; B = 16'h0056; #100;
A = 16'h0010; B = 16'h0057; #100;
A = 16'h0010; B = 16'h0058; #100;
A = 16'h0010; B = 16'h0059; #100;
A = 16'h0010; B = 16'h005A; #100;
A = 16'h0010; B = 16'h005B; #100;
A = 16'h0010; B = 16'h005C; #100;
A = 16'h0010; B = 16'h005D; #100;
A = 16'h0010; B = 16'h005E; #100;
A = 16'h0010; B = 16'h005F; #100;
A = 16'h0010; B = 16'h0060; #100;
A = 16'h0010; B = 16'h0061; #100;
A = 16'h0010; B = 16'h0062; #100;
A = 16'h0010; B = 16'h0063; #100;
A = 16'h0010; B = 16'h0064; #100;
A = 16'h0010; B = 16'h0065; #100;
A = 16'h0010; B = 16'h0066; #100;
A = 16'h0010; B = 16'h0067; #100;
A = 16'h0010; B = 16'h0068; #100;
A = 16'h0010; B = 16'h0069; #100;
A = 16'h0010; B = 16'h006A; #100;
A = 16'h0010; B = 16'h006B; #100;
A = 16'h0010; B = 16'h006C; #100;
A = 16'h0010; B = 16'h006D; #100;
A = 16'h0010; B = 16'h006E; #100;
A = 16'h0010; B = 16'h006F; #100;
A = 16'h0010; B = 16'h0070; #100;
A = 16'h0010; B = 16'h0071; #100;
A = 16'h0010; B = 16'h0072; #100;
A = 16'h0010; B = 16'h0073; #100;
A = 16'h0010; B = 16'h0074; #100;
A = 16'h0010; B = 16'h0075; #100;
A = 16'h0010; B = 16'h0076; #100;
A = 16'h0010; B = 16'h0077; #100;
A = 16'h0010; B = 16'h0078; #100;
A = 16'h0010; B = 16'h0079; #100;
A = 16'h0010; B = 16'h007A; #100;
A = 16'h0010; B = 16'h007B; #100;
A = 16'h0010; B = 16'h007C; #100;
A = 16'h0010; B = 16'h007D; #100;
A = 16'h0010; B = 16'h007E; #100;
A = 16'h0010; B = 16'h007F; #100;
A = 16'h0010; B = 16'h0080; #100;
A = 16'h0010; B = 16'h0081; #100;
A = 16'h0010; B = 16'h0082; #100;
A = 16'h0010; B = 16'h0083; #100;
A = 16'h0010; B = 16'h0084; #100;
A = 16'h0010; B = 16'h0085; #100;
A = 16'h0010; B = 16'h0086; #100;
A = 16'h0010; B = 16'h0087; #100;
A = 16'h0010; B = 16'h0088; #100;
A = 16'h0010; B = 16'h0089; #100;
A = 16'h0010; B = 16'h008A; #100;
A = 16'h0010; B = 16'h008B; #100;
A = 16'h0010; B = 16'h008C; #100;
A = 16'h0010; B = 16'h008D; #100;
A = 16'h0010; B = 16'h008E; #100;
A = 16'h0010; B = 16'h008F; #100;
A = 16'h0010; B = 16'h0090; #100;
A = 16'h0010; B = 16'h0091; #100;
A = 16'h0010; B = 16'h0092; #100;
A = 16'h0010; B = 16'h0093; #100;
A = 16'h0010; B = 16'h0094; #100;
A = 16'h0010; B = 16'h0095; #100;
A = 16'h0010; B = 16'h0096; #100;
A = 16'h0010; B = 16'h0097; #100;
A = 16'h0010; B = 16'h0098; #100;
A = 16'h0010; B = 16'h0099; #100;
A = 16'h0010; B = 16'h009A; #100;
A = 16'h0010; B = 16'h009B; #100;
A = 16'h0010; B = 16'h009C; #100;
A = 16'h0010; B = 16'h009D; #100;
A = 16'h0010; B = 16'h009E; #100;
A = 16'h0010; B = 16'h009F; #100;
A = 16'h0010; B = 16'h00A0; #100;
A = 16'h0010; B = 16'h00A1; #100;
A = 16'h0010; B = 16'h00A2; #100;
A = 16'h0010; B = 16'h00A3; #100;
A = 16'h0010; B = 16'h00A4; #100;
A = 16'h0010; B = 16'h00A5; #100;
A = 16'h0010; B = 16'h00A6; #100;
A = 16'h0010; B = 16'h00A7; #100;
A = 16'h0010; B = 16'h00A8; #100;
A = 16'h0010; B = 16'h00A9; #100;
A = 16'h0010; B = 16'h00AA; #100;
A = 16'h0010; B = 16'h00AB; #100;
A = 16'h0010; B = 16'h00AC; #100;
A = 16'h0010; B = 16'h00AD; #100;
A = 16'h0010; B = 16'h00AE; #100;
A = 16'h0010; B = 16'h00AF; #100;
A = 16'h0010; B = 16'h00B0; #100;
A = 16'h0010; B = 16'h00B1; #100;
A = 16'h0010; B = 16'h00B2; #100;
A = 16'h0010; B = 16'h00B3; #100;
A = 16'h0010; B = 16'h00B4; #100;
A = 16'h0010; B = 16'h00B5; #100;
A = 16'h0010; B = 16'h00B6; #100;
A = 16'h0010; B = 16'h00B7; #100;
A = 16'h0010; B = 16'h00B8; #100;
A = 16'h0010; B = 16'h00B9; #100;
A = 16'h0010; B = 16'h00BA; #100;
A = 16'h0010; B = 16'h00BB; #100;
A = 16'h0010; B = 16'h00BC; #100;
A = 16'h0010; B = 16'h00BD; #100;
A = 16'h0010; B = 16'h00BE; #100;
A = 16'h0010; B = 16'h00BF; #100;
A = 16'h0010; B = 16'h00C0; #100;
A = 16'h0010; B = 16'h00C1; #100;
A = 16'h0010; B = 16'h00C2; #100;
A = 16'h0010; B = 16'h00C3; #100;
A = 16'h0010; B = 16'h00C4; #100;
A = 16'h0010; B = 16'h00C5; #100;
A = 16'h0010; B = 16'h00C6; #100;
A = 16'h0010; B = 16'h00C7; #100;
A = 16'h0010; B = 16'h00C8; #100;
A = 16'h0010; B = 16'h00C9; #100;
A = 16'h0010; B = 16'h00CA; #100;
A = 16'h0010; B = 16'h00CB; #100;
A = 16'h0010; B = 16'h00CC; #100;
A = 16'h0010; B = 16'h00CD; #100;
A = 16'h0010; B = 16'h00CE; #100;
A = 16'h0010; B = 16'h00CF; #100;
A = 16'h0010; B = 16'h00D0; #100;
A = 16'h0010; B = 16'h00D1; #100;
A = 16'h0010; B = 16'h00D2; #100;
A = 16'h0010; B = 16'h00D3; #100;
A = 16'h0010; B = 16'h00D4; #100;
A = 16'h0010; B = 16'h00D5; #100;
A = 16'h0010; B = 16'h00D6; #100;
A = 16'h0010; B = 16'h00D7; #100;
A = 16'h0010; B = 16'h00D8; #100;
A = 16'h0010; B = 16'h00D9; #100;
A = 16'h0010; B = 16'h00DA; #100;
A = 16'h0010; B = 16'h00DB; #100;
A = 16'h0010; B = 16'h00DC; #100;
A = 16'h0010; B = 16'h00DD; #100;
A = 16'h0010; B = 16'h00DE; #100;
A = 16'h0010; B = 16'h00DF; #100;
A = 16'h0010; B = 16'h00E0; #100;
A = 16'h0010; B = 16'h00E1; #100;
A = 16'h0010; B = 16'h00E2; #100;
A = 16'h0010; B = 16'h00E3; #100;
A = 16'h0010; B = 16'h00E4; #100;
A = 16'h0010; B = 16'h00E5; #100;
A = 16'h0010; B = 16'h00E6; #100;
A = 16'h0010; B = 16'h00E7; #100;
A = 16'h0010; B = 16'h00E8; #100;
A = 16'h0010; B = 16'h00E9; #100;
A = 16'h0010; B = 16'h00EA; #100;
A = 16'h0010; B = 16'h00EB; #100;
A = 16'h0010; B = 16'h00EC; #100;
A = 16'h0010; B = 16'h00ED; #100;
A = 16'h0010; B = 16'h00EE; #100;
A = 16'h0010; B = 16'h00EF; #100;
A = 16'h0010; B = 16'h00F0; #100;
A = 16'h0010; B = 16'h00F1; #100;
A = 16'h0010; B = 16'h00F2; #100;
A = 16'h0010; B = 16'h00F3; #100;
A = 16'h0010; B = 16'h00F4; #100;
A = 16'h0010; B = 16'h00F5; #100;
A = 16'h0010; B = 16'h00F6; #100;
A = 16'h0010; B = 16'h00F7; #100;
A = 16'h0010; B = 16'h00F8; #100;
A = 16'h0010; B = 16'h00F9; #100;
A = 16'h0010; B = 16'h00FA; #100;
A = 16'h0010; B = 16'h00FB; #100;
A = 16'h0010; B = 16'h00FC; #100;
A = 16'h0010; B = 16'h00FD; #100;
A = 16'h0010; B = 16'h00FE; #100;
A = 16'h0010; B = 16'h00FF; #100;
A = 16'h0011; B = 16'h000; #100;
A = 16'h0011; B = 16'h001; #100;
A = 16'h0011; B = 16'h002; #100;
A = 16'h0011; B = 16'h003; #100;
A = 16'h0011; B = 16'h004; #100;
A = 16'h0011; B = 16'h005; #100;
A = 16'h0011; B = 16'h006; #100;
A = 16'h0011; B = 16'h007; #100;
A = 16'h0011; B = 16'h008; #100;
A = 16'h0011; B = 16'h009; #100;
A = 16'h0011; B = 16'h00A; #100;
A = 16'h0011; B = 16'h00B; #100;
A = 16'h0011; B = 16'h00C; #100;
A = 16'h0011; B = 16'h00D; #100;
A = 16'h0011; B = 16'h00E; #100;
A = 16'h0011; B = 16'h00F; #100;
A = 16'h0011; B = 16'h0010; #100;
A = 16'h0011; B = 16'h0011; #100;
A = 16'h0011; B = 16'h0012; #100;
A = 16'h0011; B = 16'h0013; #100;
A = 16'h0011; B = 16'h0014; #100;
A = 16'h0011; B = 16'h0015; #100;
A = 16'h0011; B = 16'h0016; #100;
A = 16'h0011; B = 16'h0017; #100;
A = 16'h0011; B = 16'h0018; #100;
A = 16'h0011; B = 16'h0019; #100;
A = 16'h0011; B = 16'h001A; #100;
A = 16'h0011; B = 16'h001B; #100;
A = 16'h0011; B = 16'h001C; #100;
A = 16'h0011; B = 16'h001D; #100;
A = 16'h0011; B = 16'h001E; #100;
A = 16'h0011; B = 16'h001F; #100;
A = 16'h0011; B = 16'h0020; #100;
A = 16'h0011; B = 16'h0021; #100;
A = 16'h0011; B = 16'h0022; #100;
A = 16'h0011; B = 16'h0023; #100;
A = 16'h0011; B = 16'h0024; #100;
A = 16'h0011; B = 16'h0025; #100;
A = 16'h0011; B = 16'h0026; #100;
A = 16'h0011; B = 16'h0027; #100;
A = 16'h0011; B = 16'h0028; #100;
A = 16'h0011; B = 16'h0029; #100;
A = 16'h0011; B = 16'h002A; #100;
A = 16'h0011; B = 16'h002B; #100;
A = 16'h0011; B = 16'h002C; #100;
A = 16'h0011; B = 16'h002D; #100;
A = 16'h0011; B = 16'h002E; #100;
A = 16'h0011; B = 16'h002F; #100;
A = 16'h0011; B = 16'h0030; #100;
A = 16'h0011; B = 16'h0031; #100;
A = 16'h0011; B = 16'h0032; #100;
A = 16'h0011; B = 16'h0033; #100;
A = 16'h0011; B = 16'h0034; #100;
A = 16'h0011; B = 16'h0035; #100;
A = 16'h0011; B = 16'h0036; #100;
A = 16'h0011; B = 16'h0037; #100;
A = 16'h0011; B = 16'h0038; #100;
A = 16'h0011; B = 16'h0039; #100;
A = 16'h0011; B = 16'h003A; #100;
A = 16'h0011; B = 16'h003B; #100;
A = 16'h0011; B = 16'h003C; #100;
A = 16'h0011; B = 16'h003D; #100;
A = 16'h0011; B = 16'h003E; #100;
A = 16'h0011; B = 16'h003F; #100;
A = 16'h0011; B = 16'h0040; #100;
A = 16'h0011; B = 16'h0041; #100;
A = 16'h0011; B = 16'h0042; #100;
A = 16'h0011; B = 16'h0043; #100;
A = 16'h0011; B = 16'h0044; #100;
A = 16'h0011; B = 16'h0045; #100;
A = 16'h0011; B = 16'h0046; #100;
A = 16'h0011; B = 16'h0047; #100;
A = 16'h0011; B = 16'h0048; #100;
A = 16'h0011; B = 16'h0049; #100;
A = 16'h0011; B = 16'h004A; #100;
A = 16'h0011; B = 16'h004B; #100;
A = 16'h0011; B = 16'h004C; #100;
A = 16'h0011; B = 16'h004D; #100;
A = 16'h0011; B = 16'h004E; #100;
A = 16'h0011; B = 16'h004F; #100;
A = 16'h0011; B = 16'h0050; #100;
A = 16'h0011; B = 16'h0051; #100;
A = 16'h0011; B = 16'h0052; #100;
A = 16'h0011; B = 16'h0053; #100;
A = 16'h0011; B = 16'h0054; #100;
A = 16'h0011; B = 16'h0055; #100;
A = 16'h0011; B = 16'h0056; #100;
A = 16'h0011; B = 16'h0057; #100;
A = 16'h0011; B = 16'h0058; #100;
A = 16'h0011; B = 16'h0059; #100;
A = 16'h0011; B = 16'h005A; #100;
A = 16'h0011; B = 16'h005B; #100;
A = 16'h0011; B = 16'h005C; #100;
A = 16'h0011; B = 16'h005D; #100;
A = 16'h0011; B = 16'h005E; #100;
A = 16'h0011; B = 16'h005F; #100;
A = 16'h0011; B = 16'h0060; #100;
A = 16'h0011; B = 16'h0061; #100;
A = 16'h0011; B = 16'h0062; #100;
A = 16'h0011; B = 16'h0063; #100;
A = 16'h0011; B = 16'h0064; #100;
A = 16'h0011; B = 16'h0065; #100;
A = 16'h0011; B = 16'h0066; #100;
A = 16'h0011; B = 16'h0067; #100;
A = 16'h0011; B = 16'h0068; #100;
A = 16'h0011; B = 16'h0069; #100;
A = 16'h0011; B = 16'h006A; #100;
A = 16'h0011; B = 16'h006B; #100;
A = 16'h0011; B = 16'h006C; #100;
A = 16'h0011; B = 16'h006D; #100;
A = 16'h0011; B = 16'h006E; #100;
A = 16'h0011; B = 16'h006F; #100;
A = 16'h0011; B = 16'h0070; #100;
A = 16'h0011; B = 16'h0071; #100;
A = 16'h0011; B = 16'h0072; #100;
A = 16'h0011; B = 16'h0073; #100;
A = 16'h0011; B = 16'h0074; #100;
A = 16'h0011; B = 16'h0075; #100;
A = 16'h0011; B = 16'h0076; #100;
A = 16'h0011; B = 16'h0077; #100;
A = 16'h0011; B = 16'h0078; #100;
A = 16'h0011; B = 16'h0079; #100;
A = 16'h0011; B = 16'h007A; #100;
A = 16'h0011; B = 16'h007B; #100;
A = 16'h0011; B = 16'h007C; #100;
A = 16'h0011; B = 16'h007D; #100;
A = 16'h0011; B = 16'h007E; #100;
A = 16'h0011; B = 16'h007F; #100;
A = 16'h0011; B = 16'h0080; #100;
A = 16'h0011; B = 16'h0081; #100;
A = 16'h0011; B = 16'h0082; #100;
A = 16'h0011; B = 16'h0083; #100;
A = 16'h0011; B = 16'h0084; #100;
A = 16'h0011; B = 16'h0085; #100;
A = 16'h0011; B = 16'h0086; #100;
A = 16'h0011; B = 16'h0087; #100;
A = 16'h0011; B = 16'h0088; #100;
A = 16'h0011; B = 16'h0089; #100;
A = 16'h0011; B = 16'h008A; #100;
A = 16'h0011; B = 16'h008B; #100;
A = 16'h0011; B = 16'h008C; #100;
A = 16'h0011; B = 16'h008D; #100;
A = 16'h0011; B = 16'h008E; #100;
A = 16'h0011; B = 16'h008F; #100;
A = 16'h0011; B = 16'h0090; #100;
A = 16'h0011; B = 16'h0091; #100;
A = 16'h0011; B = 16'h0092; #100;
A = 16'h0011; B = 16'h0093; #100;
A = 16'h0011; B = 16'h0094; #100;
A = 16'h0011; B = 16'h0095; #100;
A = 16'h0011; B = 16'h0096; #100;
A = 16'h0011; B = 16'h0097; #100;
A = 16'h0011; B = 16'h0098; #100;
A = 16'h0011; B = 16'h0099; #100;
A = 16'h0011; B = 16'h009A; #100;
A = 16'h0011; B = 16'h009B; #100;
A = 16'h0011; B = 16'h009C; #100;
A = 16'h0011; B = 16'h009D; #100;
A = 16'h0011; B = 16'h009E; #100;
A = 16'h0011; B = 16'h009F; #100;
A = 16'h0011; B = 16'h00A0; #100;
A = 16'h0011; B = 16'h00A1; #100;
A = 16'h0011; B = 16'h00A2; #100;
A = 16'h0011; B = 16'h00A3; #100;
A = 16'h0011; B = 16'h00A4; #100;
A = 16'h0011; B = 16'h00A5; #100;
A = 16'h0011; B = 16'h00A6; #100;
A = 16'h0011; B = 16'h00A7; #100;
A = 16'h0011; B = 16'h00A8; #100;
A = 16'h0011; B = 16'h00A9; #100;
A = 16'h0011; B = 16'h00AA; #100;
A = 16'h0011; B = 16'h00AB; #100;
A = 16'h0011; B = 16'h00AC; #100;
A = 16'h0011; B = 16'h00AD; #100;
A = 16'h0011; B = 16'h00AE; #100;
A = 16'h0011; B = 16'h00AF; #100;
A = 16'h0011; B = 16'h00B0; #100;
A = 16'h0011; B = 16'h00B1; #100;
A = 16'h0011; B = 16'h00B2; #100;
A = 16'h0011; B = 16'h00B3; #100;
A = 16'h0011; B = 16'h00B4; #100;
A = 16'h0011; B = 16'h00B5; #100;
A = 16'h0011; B = 16'h00B6; #100;
A = 16'h0011; B = 16'h00B7; #100;
A = 16'h0011; B = 16'h00B8; #100;
A = 16'h0011; B = 16'h00B9; #100;
A = 16'h0011; B = 16'h00BA; #100;
A = 16'h0011; B = 16'h00BB; #100;
A = 16'h0011; B = 16'h00BC; #100;
A = 16'h0011; B = 16'h00BD; #100;
A = 16'h0011; B = 16'h00BE; #100;
A = 16'h0011; B = 16'h00BF; #100;
A = 16'h0011; B = 16'h00C0; #100;
A = 16'h0011; B = 16'h00C1; #100;
A = 16'h0011; B = 16'h00C2; #100;
A = 16'h0011; B = 16'h00C3; #100;
A = 16'h0011; B = 16'h00C4; #100;
A = 16'h0011; B = 16'h00C5; #100;
A = 16'h0011; B = 16'h00C6; #100;
A = 16'h0011; B = 16'h00C7; #100;
A = 16'h0011; B = 16'h00C8; #100;
A = 16'h0011; B = 16'h00C9; #100;
A = 16'h0011; B = 16'h00CA; #100;
A = 16'h0011; B = 16'h00CB; #100;
A = 16'h0011; B = 16'h00CC; #100;
A = 16'h0011; B = 16'h00CD; #100;
A = 16'h0011; B = 16'h00CE; #100;
A = 16'h0011; B = 16'h00CF; #100;
A = 16'h0011; B = 16'h00D0; #100;
A = 16'h0011; B = 16'h00D1; #100;
A = 16'h0011; B = 16'h00D2; #100;
A = 16'h0011; B = 16'h00D3; #100;
A = 16'h0011; B = 16'h00D4; #100;
A = 16'h0011; B = 16'h00D5; #100;
A = 16'h0011; B = 16'h00D6; #100;
A = 16'h0011; B = 16'h00D7; #100;
A = 16'h0011; B = 16'h00D8; #100;
A = 16'h0011; B = 16'h00D9; #100;
A = 16'h0011; B = 16'h00DA; #100;
A = 16'h0011; B = 16'h00DB; #100;
A = 16'h0011; B = 16'h00DC; #100;
A = 16'h0011; B = 16'h00DD; #100;
A = 16'h0011; B = 16'h00DE; #100;
A = 16'h0011; B = 16'h00DF; #100;
A = 16'h0011; B = 16'h00E0; #100;
A = 16'h0011; B = 16'h00E1; #100;
A = 16'h0011; B = 16'h00E2; #100;
A = 16'h0011; B = 16'h00E3; #100;
A = 16'h0011; B = 16'h00E4; #100;
A = 16'h0011; B = 16'h00E5; #100;
A = 16'h0011; B = 16'h00E6; #100;
A = 16'h0011; B = 16'h00E7; #100;
A = 16'h0011; B = 16'h00E8; #100;
A = 16'h0011; B = 16'h00E9; #100;
A = 16'h0011; B = 16'h00EA; #100;
A = 16'h0011; B = 16'h00EB; #100;
A = 16'h0011; B = 16'h00EC; #100;
A = 16'h0011; B = 16'h00ED; #100;
A = 16'h0011; B = 16'h00EE; #100;
A = 16'h0011; B = 16'h00EF; #100;
A = 16'h0011; B = 16'h00F0; #100;
A = 16'h0011; B = 16'h00F1; #100;
A = 16'h0011; B = 16'h00F2; #100;
A = 16'h0011; B = 16'h00F3; #100;
A = 16'h0011; B = 16'h00F4; #100;
A = 16'h0011; B = 16'h00F5; #100;
A = 16'h0011; B = 16'h00F6; #100;
A = 16'h0011; B = 16'h00F7; #100;
A = 16'h0011; B = 16'h00F8; #100;
A = 16'h0011; B = 16'h00F9; #100;
A = 16'h0011; B = 16'h00FA; #100;
A = 16'h0011; B = 16'h00FB; #100;
A = 16'h0011; B = 16'h00FC; #100;
A = 16'h0011; B = 16'h00FD; #100;
A = 16'h0011; B = 16'h00FE; #100;
A = 16'h0011; B = 16'h00FF; #100;
A = 16'h0012; B = 16'h000; #100;
A = 16'h0012; B = 16'h001; #100;
A = 16'h0012; B = 16'h002; #100;
A = 16'h0012; B = 16'h003; #100;
A = 16'h0012; B = 16'h004; #100;
A = 16'h0012; B = 16'h005; #100;
A = 16'h0012; B = 16'h006; #100;
A = 16'h0012; B = 16'h007; #100;
A = 16'h0012; B = 16'h008; #100;
A = 16'h0012; B = 16'h009; #100;
A = 16'h0012; B = 16'h00A; #100;
A = 16'h0012; B = 16'h00B; #100;
A = 16'h0012; B = 16'h00C; #100;
A = 16'h0012; B = 16'h00D; #100;
A = 16'h0012; B = 16'h00E; #100;
A = 16'h0012; B = 16'h00F; #100;
A = 16'h0012; B = 16'h0010; #100;
A = 16'h0012; B = 16'h0011; #100;
A = 16'h0012; B = 16'h0012; #100;
A = 16'h0012; B = 16'h0013; #100;
A = 16'h0012; B = 16'h0014; #100;
A = 16'h0012; B = 16'h0015; #100;
A = 16'h0012; B = 16'h0016; #100;
A = 16'h0012; B = 16'h0017; #100;
A = 16'h0012; B = 16'h0018; #100;
A = 16'h0012; B = 16'h0019; #100;
A = 16'h0012; B = 16'h001A; #100;
A = 16'h0012; B = 16'h001B; #100;
A = 16'h0012; B = 16'h001C; #100;
A = 16'h0012; B = 16'h001D; #100;
A = 16'h0012; B = 16'h001E; #100;
A = 16'h0012; B = 16'h001F; #100;
A = 16'h0012; B = 16'h0020; #100;
A = 16'h0012; B = 16'h0021; #100;
A = 16'h0012; B = 16'h0022; #100;
A = 16'h0012; B = 16'h0023; #100;
A = 16'h0012; B = 16'h0024; #100;
A = 16'h0012; B = 16'h0025; #100;
A = 16'h0012; B = 16'h0026; #100;
A = 16'h0012; B = 16'h0027; #100;
A = 16'h0012; B = 16'h0028; #100;
A = 16'h0012; B = 16'h0029; #100;
A = 16'h0012; B = 16'h002A; #100;
A = 16'h0012; B = 16'h002B; #100;
A = 16'h0012; B = 16'h002C; #100;
A = 16'h0012; B = 16'h002D; #100;
A = 16'h0012; B = 16'h002E; #100;
A = 16'h0012; B = 16'h002F; #100;
A = 16'h0012; B = 16'h0030; #100;
A = 16'h0012; B = 16'h0031; #100;
A = 16'h0012; B = 16'h0032; #100;
A = 16'h0012; B = 16'h0033; #100;
A = 16'h0012; B = 16'h0034; #100;
A = 16'h0012; B = 16'h0035; #100;
A = 16'h0012; B = 16'h0036; #100;
A = 16'h0012; B = 16'h0037; #100;
A = 16'h0012; B = 16'h0038; #100;
A = 16'h0012; B = 16'h0039; #100;
A = 16'h0012; B = 16'h003A; #100;
A = 16'h0012; B = 16'h003B; #100;
A = 16'h0012; B = 16'h003C; #100;
A = 16'h0012; B = 16'h003D; #100;
A = 16'h0012; B = 16'h003E; #100;
A = 16'h0012; B = 16'h003F; #100;
A = 16'h0012; B = 16'h0040; #100;
A = 16'h0012; B = 16'h0041; #100;
A = 16'h0012; B = 16'h0042; #100;
A = 16'h0012; B = 16'h0043; #100;
A = 16'h0012; B = 16'h0044; #100;
A = 16'h0012; B = 16'h0045; #100;
A = 16'h0012; B = 16'h0046; #100;
A = 16'h0012; B = 16'h0047; #100;
A = 16'h0012; B = 16'h0048; #100;
A = 16'h0012; B = 16'h0049; #100;
A = 16'h0012; B = 16'h004A; #100;
A = 16'h0012; B = 16'h004B; #100;
A = 16'h0012; B = 16'h004C; #100;
A = 16'h0012; B = 16'h004D; #100;
A = 16'h0012; B = 16'h004E; #100;
A = 16'h0012; B = 16'h004F; #100;
A = 16'h0012; B = 16'h0050; #100;
A = 16'h0012; B = 16'h0051; #100;
A = 16'h0012; B = 16'h0052; #100;
A = 16'h0012; B = 16'h0053; #100;
A = 16'h0012; B = 16'h0054; #100;
A = 16'h0012; B = 16'h0055; #100;
A = 16'h0012; B = 16'h0056; #100;
A = 16'h0012; B = 16'h0057; #100;
A = 16'h0012; B = 16'h0058; #100;
A = 16'h0012; B = 16'h0059; #100;
A = 16'h0012; B = 16'h005A; #100;
A = 16'h0012; B = 16'h005B; #100;
A = 16'h0012; B = 16'h005C; #100;
A = 16'h0012; B = 16'h005D; #100;
A = 16'h0012; B = 16'h005E; #100;
A = 16'h0012; B = 16'h005F; #100;
A = 16'h0012; B = 16'h0060; #100;
A = 16'h0012; B = 16'h0061; #100;
A = 16'h0012; B = 16'h0062; #100;
A = 16'h0012; B = 16'h0063; #100;
A = 16'h0012; B = 16'h0064; #100;
A = 16'h0012; B = 16'h0065; #100;
A = 16'h0012; B = 16'h0066; #100;
A = 16'h0012; B = 16'h0067; #100;
A = 16'h0012; B = 16'h0068; #100;
A = 16'h0012; B = 16'h0069; #100;
A = 16'h0012; B = 16'h006A; #100;
A = 16'h0012; B = 16'h006B; #100;
A = 16'h0012; B = 16'h006C; #100;
A = 16'h0012; B = 16'h006D; #100;
A = 16'h0012; B = 16'h006E; #100;
A = 16'h0012; B = 16'h006F; #100;
A = 16'h0012; B = 16'h0070; #100;
A = 16'h0012; B = 16'h0071; #100;
A = 16'h0012; B = 16'h0072; #100;
A = 16'h0012; B = 16'h0073; #100;
A = 16'h0012; B = 16'h0074; #100;
A = 16'h0012; B = 16'h0075; #100;
A = 16'h0012; B = 16'h0076; #100;
A = 16'h0012; B = 16'h0077; #100;
A = 16'h0012; B = 16'h0078; #100;
A = 16'h0012; B = 16'h0079; #100;
A = 16'h0012; B = 16'h007A; #100;
A = 16'h0012; B = 16'h007B; #100;
A = 16'h0012; B = 16'h007C; #100;
A = 16'h0012; B = 16'h007D; #100;
A = 16'h0012; B = 16'h007E; #100;
A = 16'h0012; B = 16'h007F; #100;
A = 16'h0012; B = 16'h0080; #100;
A = 16'h0012; B = 16'h0081; #100;
A = 16'h0012; B = 16'h0082; #100;
A = 16'h0012; B = 16'h0083; #100;
A = 16'h0012; B = 16'h0084; #100;
A = 16'h0012; B = 16'h0085; #100;
A = 16'h0012; B = 16'h0086; #100;
A = 16'h0012; B = 16'h0087; #100;
A = 16'h0012; B = 16'h0088; #100;
A = 16'h0012; B = 16'h0089; #100;
A = 16'h0012; B = 16'h008A; #100;
A = 16'h0012; B = 16'h008B; #100;
A = 16'h0012; B = 16'h008C; #100;
A = 16'h0012; B = 16'h008D; #100;
A = 16'h0012; B = 16'h008E; #100;
A = 16'h0012; B = 16'h008F; #100;
A = 16'h0012; B = 16'h0090; #100;
A = 16'h0012; B = 16'h0091; #100;
A = 16'h0012; B = 16'h0092; #100;
A = 16'h0012; B = 16'h0093; #100;
A = 16'h0012; B = 16'h0094; #100;
A = 16'h0012; B = 16'h0095; #100;
A = 16'h0012; B = 16'h0096; #100;
A = 16'h0012; B = 16'h0097; #100;
A = 16'h0012; B = 16'h0098; #100;
A = 16'h0012; B = 16'h0099; #100;
A = 16'h0012; B = 16'h009A; #100;
A = 16'h0012; B = 16'h009B; #100;
A = 16'h0012; B = 16'h009C; #100;
A = 16'h0012; B = 16'h009D; #100;
A = 16'h0012; B = 16'h009E; #100;
A = 16'h0012; B = 16'h009F; #100;
A = 16'h0012; B = 16'h00A0; #100;
A = 16'h0012; B = 16'h00A1; #100;
A = 16'h0012; B = 16'h00A2; #100;
A = 16'h0012; B = 16'h00A3; #100;
A = 16'h0012; B = 16'h00A4; #100;
A = 16'h0012; B = 16'h00A5; #100;
A = 16'h0012; B = 16'h00A6; #100;
A = 16'h0012; B = 16'h00A7; #100;
A = 16'h0012; B = 16'h00A8; #100;
A = 16'h0012; B = 16'h00A9; #100;
A = 16'h0012; B = 16'h00AA; #100;
A = 16'h0012; B = 16'h00AB; #100;
A = 16'h0012; B = 16'h00AC; #100;
A = 16'h0012; B = 16'h00AD; #100;
A = 16'h0012; B = 16'h00AE; #100;
A = 16'h0012; B = 16'h00AF; #100;
A = 16'h0012; B = 16'h00B0; #100;
A = 16'h0012; B = 16'h00B1; #100;
A = 16'h0012; B = 16'h00B2; #100;
A = 16'h0012; B = 16'h00B3; #100;
A = 16'h0012; B = 16'h00B4; #100;
A = 16'h0012; B = 16'h00B5; #100;
A = 16'h0012; B = 16'h00B6; #100;
A = 16'h0012; B = 16'h00B7; #100;
A = 16'h0012; B = 16'h00B8; #100;
A = 16'h0012; B = 16'h00B9; #100;
A = 16'h0012; B = 16'h00BA; #100;
A = 16'h0012; B = 16'h00BB; #100;
A = 16'h0012; B = 16'h00BC; #100;
A = 16'h0012; B = 16'h00BD; #100;
A = 16'h0012; B = 16'h00BE; #100;
A = 16'h0012; B = 16'h00BF; #100;
A = 16'h0012; B = 16'h00C0; #100;
A = 16'h0012; B = 16'h00C1; #100;
A = 16'h0012; B = 16'h00C2; #100;
A = 16'h0012; B = 16'h00C3; #100;
A = 16'h0012; B = 16'h00C4; #100;
A = 16'h0012; B = 16'h00C5; #100;
A = 16'h0012; B = 16'h00C6; #100;
A = 16'h0012; B = 16'h00C7; #100;
A = 16'h0012; B = 16'h00C8; #100;
A = 16'h0012; B = 16'h00C9; #100;
A = 16'h0012; B = 16'h00CA; #100;
A = 16'h0012; B = 16'h00CB; #100;
A = 16'h0012; B = 16'h00CC; #100;
A = 16'h0012; B = 16'h00CD; #100;
A = 16'h0012; B = 16'h00CE; #100;
A = 16'h0012; B = 16'h00CF; #100;
A = 16'h0012; B = 16'h00D0; #100;
A = 16'h0012; B = 16'h00D1; #100;
A = 16'h0012; B = 16'h00D2; #100;
A = 16'h0012; B = 16'h00D3; #100;
A = 16'h0012; B = 16'h00D4; #100;
A = 16'h0012; B = 16'h00D5; #100;
A = 16'h0012; B = 16'h00D6; #100;
A = 16'h0012; B = 16'h00D7; #100;
A = 16'h0012; B = 16'h00D8; #100;
A = 16'h0012; B = 16'h00D9; #100;
A = 16'h0012; B = 16'h00DA; #100;
A = 16'h0012; B = 16'h00DB; #100;
A = 16'h0012; B = 16'h00DC; #100;
A = 16'h0012; B = 16'h00DD; #100;
A = 16'h0012; B = 16'h00DE; #100;
A = 16'h0012; B = 16'h00DF; #100;
A = 16'h0012; B = 16'h00E0; #100;
A = 16'h0012; B = 16'h00E1; #100;
A = 16'h0012; B = 16'h00E2; #100;
A = 16'h0012; B = 16'h00E3; #100;
A = 16'h0012; B = 16'h00E4; #100;
A = 16'h0012; B = 16'h00E5; #100;
A = 16'h0012; B = 16'h00E6; #100;
A = 16'h0012; B = 16'h00E7; #100;
A = 16'h0012; B = 16'h00E8; #100;
A = 16'h0012; B = 16'h00E9; #100;
A = 16'h0012; B = 16'h00EA; #100;
A = 16'h0012; B = 16'h00EB; #100;
A = 16'h0012; B = 16'h00EC; #100;
A = 16'h0012; B = 16'h00ED; #100;
A = 16'h0012; B = 16'h00EE; #100;
A = 16'h0012; B = 16'h00EF; #100;
A = 16'h0012; B = 16'h00F0; #100;
A = 16'h0012; B = 16'h00F1; #100;
A = 16'h0012; B = 16'h00F2; #100;
A = 16'h0012; B = 16'h00F3; #100;
A = 16'h0012; B = 16'h00F4; #100;
A = 16'h0012; B = 16'h00F5; #100;
A = 16'h0012; B = 16'h00F6; #100;
A = 16'h0012; B = 16'h00F7; #100;
A = 16'h0012; B = 16'h00F8; #100;
A = 16'h0012; B = 16'h00F9; #100;
A = 16'h0012; B = 16'h00FA; #100;
A = 16'h0012; B = 16'h00FB; #100;
A = 16'h0012; B = 16'h00FC; #100;
A = 16'h0012; B = 16'h00FD; #100;
A = 16'h0012; B = 16'h00FE; #100;
A = 16'h0012; B = 16'h00FF; #100;
A = 16'h0013; B = 16'h000; #100;
A = 16'h0013; B = 16'h001; #100;
A = 16'h0013; B = 16'h002; #100;
A = 16'h0013; B = 16'h003; #100;
A = 16'h0013; B = 16'h004; #100;
A = 16'h0013; B = 16'h005; #100;
A = 16'h0013; B = 16'h006; #100;
A = 16'h0013; B = 16'h007; #100;
A = 16'h0013; B = 16'h008; #100;
A = 16'h0013; B = 16'h009; #100;
A = 16'h0013; B = 16'h00A; #100;
A = 16'h0013; B = 16'h00B; #100;
A = 16'h0013; B = 16'h00C; #100;
A = 16'h0013; B = 16'h00D; #100;
A = 16'h0013; B = 16'h00E; #100;
A = 16'h0013; B = 16'h00F; #100;
A = 16'h0013; B = 16'h0010; #100;
A = 16'h0013; B = 16'h0011; #100;
A = 16'h0013; B = 16'h0012; #100;
A = 16'h0013; B = 16'h0013; #100;
A = 16'h0013; B = 16'h0014; #100;
A = 16'h0013; B = 16'h0015; #100;
A = 16'h0013; B = 16'h0016; #100;
A = 16'h0013; B = 16'h0017; #100;
A = 16'h0013; B = 16'h0018; #100;
A = 16'h0013; B = 16'h0019; #100;
A = 16'h0013; B = 16'h001A; #100;
A = 16'h0013; B = 16'h001B; #100;
A = 16'h0013; B = 16'h001C; #100;
A = 16'h0013; B = 16'h001D; #100;
A = 16'h0013; B = 16'h001E; #100;
A = 16'h0013; B = 16'h001F; #100;
A = 16'h0013; B = 16'h0020; #100;
A = 16'h0013; B = 16'h0021; #100;
A = 16'h0013; B = 16'h0022; #100;
A = 16'h0013; B = 16'h0023; #100;
A = 16'h0013; B = 16'h0024; #100;
A = 16'h0013; B = 16'h0025; #100;
A = 16'h0013; B = 16'h0026; #100;
A = 16'h0013; B = 16'h0027; #100;
A = 16'h0013; B = 16'h0028; #100;
A = 16'h0013; B = 16'h0029; #100;
A = 16'h0013; B = 16'h002A; #100;
A = 16'h0013; B = 16'h002B; #100;
A = 16'h0013; B = 16'h002C; #100;
A = 16'h0013; B = 16'h002D; #100;
A = 16'h0013; B = 16'h002E; #100;
A = 16'h0013; B = 16'h002F; #100;
A = 16'h0013; B = 16'h0030; #100;
A = 16'h0013; B = 16'h0031; #100;
A = 16'h0013; B = 16'h0032; #100;
A = 16'h0013; B = 16'h0033; #100;
A = 16'h0013; B = 16'h0034; #100;
A = 16'h0013; B = 16'h0035; #100;
A = 16'h0013; B = 16'h0036; #100;
A = 16'h0013; B = 16'h0037; #100;
A = 16'h0013; B = 16'h0038; #100;
A = 16'h0013; B = 16'h0039; #100;
A = 16'h0013; B = 16'h003A; #100;
A = 16'h0013; B = 16'h003B; #100;
A = 16'h0013; B = 16'h003C; #100;
A = 16'h0013; B = 16'h003D; #100;
A = 16'h0013; B = 16'h003E; #100;
A = 16'h0013; B = 16'h003F; #100;
A = 16'h0013; B = 16'h0040; #100;
A = 16'h0013; B = 16'h0041; #100;
A = 16'h0013; B = 16'h0042; #100;
A = 16'h0013; B = 16'h0043; #100;
A = 16'h0013; B = 16'h0044; #100;
A = 16'h0013; B = 16'h0045; #100;
A = 16'h0013; B = 16'h0046; #100;
A = 16'h0013; B = 16'h0047; #100;
A = 16'h0013; B = 16'h0048; #100;
A = 16'h0013; B = 16'h0049; #100;
A = 16'h0013; B = 16'h004A; #100;
A = 16'h0013; B = 16'h004B; #100;
A = 16'h0013; B = 16'h004C; #100;
A = 16'h0013; B = 16'h004D; #100;
A = 16'h0013; B = 16'h004E; #100;
A = 16'h0013; B = 16'h004F; #100;
A = 16'h0013; B = 16'h0050; #100;
A = 16'h0013; B = 16'h0051; #100;
A = 16'h0013; B = 16'h0052; #100;
A = 16'h0013; B = 16'h0053; #100;
A = 16'h0013; B = 16'h0054; #100;
A = 16'h0013; B = 16'h0055; #100;
A = 16'h0013; B = 16'h0056; #100;
A = 16'h0013; B = 16'h0057; #100;
A = 16'h0013; B = 16'h0058; #100;
A = 16'h0013; B = 16'h0059; #100;
A = 16'h0013; B = 16'h005A; #100;
A = 16'h0013; B = 16'h005B; #100;
A = 16'h0013; B = 16'h005C; #100;
A = 16'h0013; B = 16'h005D; #100;
A = 16'h0013; B = 16'h005E; #100;
A = 16'h0013; B = 16'h005F; #100;
A = 16'h0013; B = 16'h0060; #100;
A = 16'h0013; B = 16'h0061; #100;
A = 16'h0013; B = 16'h0062; #100;
A = 16'h0013; B = 16'h0063; #100;
A = 16'h0013; B = 16'h0064; #100;
A = 16'h0013; B = 16'h0065; #100;
A = 16'h0013; B = 16'h0066; #100;
A = 16'h0013; B = 16'h0067; #100;
A = 16'h0013; B = 16'h0068; #100;
A = 16'h0013; B = 16'h0069; #100;
A = 16'h0013; B = 16'h006A; #100;
A = 16'h0013; B = 16'h006B; #100;
A = 16'h0013; B = 16'h006C; #100;
A = 16'h0013; B = 16'h006D; #100;
A = 16'h0013; B = 16'h006E; #100;
A = 16'h0013; B = 16'h006F; #100;
A = 16'h0013; B = 16'h0070; #100;
A = 16'h0013; B = 16'h0071; #100;
A = 16'h0013; B = 16'h0072; #100;
A = 16'h0013; B = 16'h0073; #100;
A = 16'h0013; B = 16'h0074; #100;
A = 16'h0013; B = 16'h0075; #100;
A = 16'h0013; B = 16'h0076; #100;
A = 16'h0013; B = 16'h0077; #100;
A = 16'h0013; B = 16'h0078; #100;
A = 16'h0013; B = 16'h0079; #100;
A = 16'h0013; B = 16'h007A; #100;
A = 16'h0013; B = 16'h007B; #100;
A = 16'h0013; B = 16'h007C; #100;
A = 16'h0013; B = 16'h007D; #100;
A = 16'h0013; B = 16'h007E; #100;
A = 16'h0013; B = 16'h007F; #100;
A = 16'h0013; B = 16'h0080; #100;
A = 16'h0013; B = 16'h0081; #100;
A = 16'h0013; B = 16'h0082; #100;
A = 16'h0013; B = 16'h0083; #100;
A = 16'h0013; B = 16'h0084; #100;
A = 16'h0013; B = 16'h0085; #100;
A = 16'h0013; B = 16'h0086; #100;
A = 16'h0013; B = 16'h0087; #100;
A = 16'h0013; B = 16'h0088; #100;
A = 16'h0013; B = 16'h0089; #100;
A = 16'h0013; B = 16'h008A; #100;
A = 16'h0013; B = 16'h008B; #100;
A = 16'h0013; B = 16'h008C; #100;
A = 16'h0013; B = 16'h008D; #100;
A = 16'h0013; B = 16'h008E; #100;
A = 16'h0013; B = 16'h008F; #100;
A = 16'h0013; B = 16'h0090; #100;
A = 16'h0013; B = 16'h0091; #100;
A = 16'h0013; B = 16'h0092; #100;
A = 16'h0013; B = 16'h0093; #100;
A = 16'h0013; B = 16'h0094; #100;
A = 16'h0013; B = 16'h0095; #100;
A = 16'h0013; B = 16'h0096; #100;
A = 16'h0013; B = 16'h0097; #100;
A = 16'h0013; B = 16'h0098; #100;
A = 16'h0013; B = 16'h0099; #100;
A = 16'h0013; B = 16'h009A; #100;
A = 16'h0013; B = 16'h009B; #100;
A = 16'h0013; B = 16'h009C; #100;
A = 16'h0013; B = 16'h009D; #100;
A = 16'h0013; B = 16'h009E; #100;
A = 16'h0013; B = 16'h009F; #100;
A = 16'h0013; B = 16'h00A0; #100;
A = 16'h0013; B = 16'h00A1; #100;
A = 16'h0013; B = 16'h00A2; #100;
A = 16'h0013; B = 16'h00A3; #100;
A = 16'h0013; B = 16'h00A4; #100;
A = 16'h0013; B = 16'h00A5; #100;
A = 16'h0013; B = 16'h00A6; #100;
A = 16'h0013; B = 16'h00A7; #100;
A = 16'h0013; B = 16'h00A8; #100;
A = 16'h0013; B = 16'h00A9; #100;
A = 16'h0013; B = 16'h00AA; #100;
A = 16'h0013; B = 16'h00AB; #100;
A = 16'h0013; B = 16'h00AC; #100;
A = 16'h0013; B = 16'h00AD; #100;
A = 16'h0013; B = 16'h00AE; #100;
A = 16'h0013; B = 16'h00AF; #100;
A = 16'h0013; B = 16'h00B0; #100;
A = 16'h0013; B = 16'h00B1; #100;
A = 16'h0013; B = 16'h00B2; #100;
A = 16'h0013; B = 16'h00B3; #100;
A = 16'h0013; B = 16'h00B4; #100;
A = 16'h0013; B = 16'h00B5; #100;
A = 16'h0013; B = 16'h00B6; #100;
A = 16'h0013; B = 16'h00B7; #100;
A = 16'h0013; B = 16'h00B8; #100;
A = 16'h0013; B = 16'h00B9; #100;
A = 16'h0013; B = 16'h00BA; #100;
A = 16'h0013; B = 16'h00BB; #100;
A = 16'h0013; B = 16'h00BC; #100;
A = 16'h0013; B = 16'h00BD; #100;
A = 16'h0013; B = 16'h00BE; #100;
A = 16'h0013; B = 16'h00BF; #100;
A = 16'h0013; B = 16'h00C0; #100;
A = 16'h0013; B = 16'h00C1; #100;
A = 16'h0013; B = 16'h00C2; #100;
A = 16'h0013; B = 16'h00C3; #100;
A = 16'h0013; B = 16'h00C4; #100;
A = 16'h0013; B = 16'h00C5; #100;
A = 16'h0013; B = 16'h00C6; #100;
A = 16'h0013; B = 16'h00C7; #100;
A = 16'h0013; B = 16'h00C8; #100;
A = 16'h0013; B = 16'h00C9; #100;
A = 16'h0013; B = 16'h00CA; #100;
A = 16'h0013; B = 16'h00CB; #100;
A = 16'h0013; B = 16'h00CC; #100;
A = 16'h0013; B = 16'h00CD; #100;
A = 16'h0013; B = 16'h00CE; #100;
A = 16'h0013; B = 16'h00CF; #100;
A = 16'h0013; B = 16'h00D0; #100;
A = 16'h0013; B = 16'h00D1; #100;
A = 16'h0013; B = 16'h00D2; #100;
A = 16'h0013; B = 16'h00D3; #100;
A = 16'h0013; B = 16'h00D4; #100;
A = 16'h0013; B = 16'h00D5; #100;
A = 16'h0013; B = 16'h00D6; #100;
A = 16'h0013; B = 16'h00D7; #100;
A = 16'h0013; B = 16'h00D8; #100;
A = 16'h0013; B = 16'h00D9; #100;
A = 16'h0013; B = 16'h00DA; #100;
A = 16'h0013; B = 16'h00DB; #100;
A = 16'h0013; B = 16'h00DC; #100;
A = 16'h0013; B = 16'h00DD; #100;
A = 16'h0013; B = 16'h00DE; #100;
A = 16'h0013; B = 16'h00DF; #100;
A = 16'h0013; B = 16'h00E0; #100;
A = 16'h0013; B = 16'h00E1; #100;
A = 16'h0013; B = 16'h00E2; #100;
A = 16'h0013; B = 16'h00E3; #100;
A = 16'h0013; B = 16'h00E4; #100;
A = 16'h0013; B = 16'h00E5; #100;
A = 16'h0013; B = 16'h00E6; #100;
A = 16'h0013; B = 16'h00E7; #100;
A = 16'h0013; B = 16'h00E8; #100;
A = 16'h0013; B = 16'h00E9; #100;
A = 16'h0013; B = 16'h00EA; #100;
A = 16'h0013; B = 16'h00EB; #100;
A = 16'h0013; B = 16'h00EC; #100;
A = 16'h0013; B = 16'h00ED; #100;
A = 16'h0013; B = 16'h00EE; #100;
A = 16'h0013; B = 16'h00EF; #100;
A = 16'h0013; B = 16'h00F0; #100;
A = 16'h0013; B = 16'h00F1; #100;
A = 16'h0013; B = 16'h00F2; #100;
A = 16'h0013; B = 16'h00F3; #100;
A = 16'h0013; B = 16'h00F4; #100;
A = 16'h0013; B = 16'h00F5; #100;
A = 16'h0013; B = 16'h00F6; #100;
A = 16'h0013; B = 16'h00F7; #100;
A = 16'h0013; B = 16'h00F8; #100;
A = 16'h0013; B = 16'h00F9; #100;
A = 16'h0013; B = 16'h00FA; #100;
A = 16'h0013; B = 16'h00FB; #100;
A = 16'h0013; B = 16'h00FC; #100;
A = 16'h0013; B = 16'h00FD; #100;
A = 16'h0013; B = 16'h00FE; #100;
A = 16'h0013; B = 16'h00FF; #100;
A = 16'h0014; B = 16'h000; #100;
A = 16'h0014; B = 16'h001; #100;
A = 16'h0014; B = 16'h002; #100;
A = 16'h0014; B = 16'h003; #100;
A = 16'h0014; B = 16'h004; #100;
A = 16'h0014; B = 16'h005; #100;
A = 16'h0014; B = 16'h006; #100;
A = 16'h0014; B = 16'h007; #100;
A = 16'h0014; B = 16'h008; #100;
A = 16'h0014; B = 16'h009; #100;
A = 16'h0014; B = 16'h00A; #100;
A = 16'h0014; B = 16'h00B; #100;
A = 16'h0014; B = 16'h00C; #100;
A = 16'h0014; B = 16'h00D; #100;
A = 16'h0014; B = 16'h00E; #100;
A = 16'h0014; B = 16'h00F; #100;
A = 16'h0014; B = 16'h0010; #100;
A = 16'h0014; B = 16'h0011; #100;
A = 16'h0014; B = 16'h0012; #100;
A = 16'h0014; B = 16'h0013; #100;
A = 16'h0014; B = 16'h0014; #100;
A = 16'h0014; B = 16'h0015; #100;
A = 16'h0014; B = 16'h0016; #100;
A = 16'h0014; B = 16'h0017; #100;
A = 16'h0014; B = 16'h0018; #100;
A = 16'h0014; B = 16'h0019; #100;
A = 16'h0014; B = 16'h001A; #100;
A = 16'h0014; B = 16'h001B; #100;
A = 16'h0014; B = 16'h001C; #100;
A = 16'h0014; B = 16'h001D; #100;
A = 16'h0014; B = 16'h001E; #100;
A = 16'h0014; B = 16'h001F; #100;
A = 16'h0014; B = 16'h0020; #100;
A = 16'h0014; B = 16'h0021; #100;
A = 16'h0014; B = 16'h0022; #100;
A = 16'h0014; B = 16'h0023; #100;
A = 16'h0014; B = 16'h0024; #100;
A = 16'h0014; B = 16'h0025; #100;
A = 16'h0014; B = 16'h0026; #100;
A = 16'h0014; B = 16'h0027; #100;
A = 16'h0014; B = 16'h0028; #100;
A = 16'h0014; B = 16'h0029; #100;
A = 16'h0014; B = 16'h002A; #100;
A = 16'h0014; B = 16'h002B; #100;
A = 16'h0014; B = 16'h002C; #100;
A = 16'h0014; B = 16'h002D; #100;
A = 16'h0014; B = 16'h002E; #100;
A = 16'h0014; B = 16'h002F; #100;
A = 16'h0014; B = 16'h0030; #100;
A = 16'h0014; B = 16'h0031; #100;
A = 16'h0014; B = 16'h0032; #100;
A = 16'h0014; B = 16'h0033; #100;
A = 16'h0014; B = 16'h0034; #100;
A = 16'h0014; B = 16'h0035; #100;
A = 16'h0014; B = 16'h0036; #100;
A = 16'h0014; B = 16'h0037; #100;
A = 16'h0014; B = 16'h0038; #100;
A = 16'h0014; B = 16'h0039; #100;
A = 16'h0014; B = 16'h003A; #100;
A = 16'h0014; B = 16'h003B; #100;
A = 16'h0014; B = 16'h003C; #100;
A = 16'h0014; B = 16'h003D; #100;
A = 16'h0014; B = 16'h003E; #100;
A = 16'h0014; B = 16'h003F; #100;
A = 16'h0014; B = 16'h0040; #100;
A = 16'h0014; B = 16'h0041; #100;
A = 16'h0014; B = 16'h0042; #100;
A = 16'h0014; B = 16'h0043; #100;
A = 16'h0014; B = 16'h0044; #100;
A = 16'h0014; B = 16'h0045; #100;
A = 16'h0014; B = 16'h0046; #100;
A = 16'h0014; B = 16'h0047; #100;
A = 16'h0014; B = 16'h0048; #100;
A = 16'h0014; B = 16'h0049; #100;
A = 16'h0014; B = 16'h004A; #100;
A = 16'h0014; B = 16'h004B; #100;
A = 16'h0014; B = 16'h004C; #100;
A = 16'h0014; B = 16'h004D; #100;
A = 16'h0014; B = 16'h004E; #100;
A = 16'h0014; B = 16'h004F; #100;
A = 16'h0014; B = 16'h0050; #100;
A = 16'h0014; B = 16'h0051; #100;
A = 16'h0014; B = 16'h0052; #100;
A = 16'h0014; B = 16'h0053; #100;
A = 16'h0014; B = 16'h0054; #100;
A = 16'h0014; B = 16'h0055; #100;
A = 16'h0014; B = 16'h0056; #100;
A = 16'h0014; B = 16'h0057; #100;
A = 16'h0014; B = 16'h0058; #100;
A = 16'h0014; B = 16'h0059; #100;
A = 16'h0014; B = 16'h005A; #100;
A = 16'h0014; B = 16'h005B; #100;
A = 16'h0014; B = 16'h005C; #100;
A = 16'h0014; B = 16'h005D; #100;
A = 16'h0014; B = 16'h005E; #100;
A = 16'h0014; B = 16'h005F; #100;
A = 16'h0014; B = 16'h0060; #100;
A = 16'h0014; B = 16'h0061; #100;
A = 16'h0014; B = 16'h0062; #100;
A = 16'h0014; B = 16'h0063; #100;
A = 16'h0014; B = 16'h0064; #100;
A = 16'h0014; B = 16'h0065; #100;
A = 16'h0014; B = 16'h0066; #100;
A = 16'h0014; B = 16'h0067; #100;
A = 16'h0014; B = 16'h0068; #100;
A = 16'h0014; B = 16'h0069; #100;
A = 16'h0014; B = 16'h006A; #100;
A = 16'h0014; B = 16'h006B; #100;
A = 16'h0014; B = 16'h006C; #100;
A = 16'h0014; B = 16'h006D; #100;
A = 16'h0014; B = 16'h006E; #100;
A = 16'h0014; B = 16'h006F; #100;
A = 16'h0014; B = 16'h0070; #100;
A = 16'h0014; B = 16'h0071; #100;
A = 16'h0014; B = 16'h0072; #100;
A = 16'h0014; B = 16'h0073; #100;
A = 16'h0014; B = 16'h0074; #100;
A = 16'h0014; B = 16'h0075; #100;
A = 16'h0014; B = 16'h0076; #100;
A = 16'h0014; B = 16'h0077; #100;
A = 16'h0014; B = 16'h0078; #100;
A = 16'h0014; B = 16'h0079; #100;
A = 16'h0014; B = 16'h007A; #100;
A = 16'h0014; B = 16'h007B; #100;
A = 16'h0014; B = 16'h007C; #100;
A = 16'h0014; B = 16'h007D; #100;
A = 16'h0014; B = 16'h007E; #100;
A = 16'h0014; B = 16'h007F; #100;
A = 16'h0014; B = 16'h0080; #100;
A = 16'h0014; B = 16'h0081; #100;
A = 16'h0014; B = 16'h0082; #100;
A = 16'h0014; B = 16'h0083; #100;
A = 16'h0014; B = 16'h0084; #100;
A = 16'h0014; B = 16'h0085; #100;
A = 16'h0014; B = 16'h0086; #100;
A = 16'h0014; B = 16'h0087; #100;
A = 16'h0014; B = 16'h0088; #100;
A = 16'h0014; B = 16'h0089; #100;
A = 16'h0014; B = 16'h008A; #100;
A = 16'h0014; B = 16'h008B; #100;
A = 16'h0014; B = 16'h008C; #100;
A = 16'h0014; B = 16'h008D; #100;
A = 16'h0014; B = 16'h008E; #100;
A = 16'h0014; B = 16'h008F; #100;
A = 16'h0014; B = 16'h0090; #100;
A = 16'h0014; B = 16'h0091; #100;
A = 16'h0014; B = 16'h0092; #100;
A = 16'h0014; B = 16'h0093; #100;
A = 16'h0014; B = 16'h0094; #100;
A = 16'h0014; B = 16'h0095; #100;
A = 16'h0014; B = 16'h0096; #100;
A = 16'h0014; B = 16'h0097; #100;
A = 16'h0014; B = 16'h0098; #100;
A = 16'h0014; B = 16'h0099; #100;
A = 16'h0014; B = 16'h009A; #100;
A = 16'h0014; B = 16'h009B; #100;
A = 16'h0014; B = 16'h009C; #100;
A = 16'h0014; B = 16'h009D; #100;
A = 16'h0014; B = 16'h009E; #100;
A = 16'h0014; B = 16'h009F; #100;
A = 16'h0014; B = 16'h00A0; #100;
A = 16'h0014; B = 16'h00A1; #100;
A = 16'h0014; B = 16'h00A2; #100;
A = 16'h0014; B = 16'h00A3; #100;
A = 16'h0014; B = 16'h00A4; #100;
A = 16'h0014; B = 16'h00A5; #100;
A = 16'h0014; B = 16'h00A6; #100;
A = 16'h0014; B = 16'h00A7; #100;
A = 16'h0014; B = 16'h00A8; #100;
A = 16'h0014; B = 16'h00A9; #100;
A = 16'h0014; B = 16'h00AA; #100;
A = 16'h0014; B = 16'h00AB; #100;
A = 16'h0014; B = 16'h00AC; #100;
A = 16'h0014; B = 16'h00AD; #100;
A = 16'h0014; B = 16'h00AE; #100;
A = 16'h0014; B = 16'h00AF; #100;
A = 16'h0014; B = 16'h00B0; #100;
A = 16'h0014; B = 16'h00B1; #100;
A = 16'h0014; B = 16'h00B2; #100;
A = 16'h0014; B = 16'h00B3; #100;
A = 16'h0014; B = 16'h00B4; #100;
A = 16'h0014; B = 16'h00B5; #100;
A = 16'h0014; B = 16'h00B6; #100;
A = 16'h0014; B = 16'h00B7; #100;
A = 16'h0014; B = 16'h00B8; #100;
A = 16'h0014; B = 16'h00B9; #100;
A = 16'h0014; B = 16'h00BA; #100;
A = 16'h0014; B = 16'h00BB; #100;
A = 16'h0014; B = 16'h00BC; #100;
A = 16'h0014; B = 16'h00BD; #100;
A = 16'h0014; B = 16'h00BE; #100;
A = 16'h0014; B = 16'h00BF; #100;
A = 16'h0014; B = 16'h00C0; #100;
A = 16'h0014; B = 16'h00C1; #100;
A = 16'h0014; B = 16'h00C2; #100;
A = 16'h0014; B = 16'h00C3; #100;
A = 16'h0014; B = 16'h00C4; #100;
A = 16'h0014; B = 16'h00C5; #100;
A = 16'h0014; B = 16'h00C6; #100;
A = 16'h0014; B = 16'h00C7; #100;
A = 16'h0014; B = 16'h00C8; #100;
A = 16'h0014; B = 16'h00C9; #100;
A = 16'h0014; B = 16'h00CA; #100;
A = 16'h0014; B = 16'h00CB; #100;
A = 16'h0014; B = 16'h00CC; #100;
A = 16'h0014; B = 16'h00CD; #100;
A = 16'h0014; B = 16'h00CE; #100;
A = 16'h0014; B = 16'h00CF; #100;
A = 16'h0014; B = 16'h00D0; #100;
A = 16'h0014; B = 16'h00D1; #100;
A = 16'h0014; B = 16'h00D2; #100;
A = 16'h0014; B = 16'h00D3; #100;
A = 16'h0014; B = 16'h00D4; #100;
A = 16'h0014; B = 16'h00D5; #100;
A = 16'h0014; B = 16'h00D6; #100;
A = 16'h0014; B = 16'h00D7; #100;
A = 16'h0014; B = 16'h00D8; #100;
A = 16'h0014; B = 16'h00D9; #100;
A = 16'h0014; B = 16'h00DA; #100;
A = 16'h0014; B = 16'h00DB; #100;
A = 16'h0014; B = 16'h00DC; #100;
A = 16'h0014; B = 16'h00DD; #100;
A = 16'h0014; B = 16'h00DE; #100;
A = 16'h0014; B = 16'h00DF; #100;
A = 16'h0014; B = 16'h00E0; #100;
A = 16'h0014; B = 16'h00E1; #100;
A = 16'h0014; B = 16'h00E2; #100;
A = 16'h0014; B = 16'h00E3; #100;
A = 16'h0014; B = 16'h00E4; #100;
A = 16'h0014; B = 16'h00E5; #100;
A = 16'h0014; B = 16'h00E6; #100;
A = 16'h0014; B = 16'h00E7; #100;
A = 16'h0014; B = 16'h00E8; #100;
A = 16'h0014; B = 16'h00E9; #100;
A = 16'h0014; B = 16'h00EA; #100;
A = 16'h0014; B = 16'h00EB; #100;
A = 16'h0014; B = 16'h00EC; #100;
A = 16'h0014; B = 16'h00ED; #100;
A = 16'h0014; B = 16'h00EE; #100;
A = 16'h0014; B = 16'h00EF; #100;
A = 16'h0014; B = 16'h00F0; #100;
A = 16'h0014; B = 16'h00F1; #100;
A = 16'h0014; B = 16'h00F2; #100;
A = 16'h0014; B = 16'h00F3; #100;
A = 16'h0014; B = 16'h00F4; #100;
A = 16'h0014; B = 16'h00F5; #100;
A = 16'h0014; B = 16'h00F6; #100;
A = 16'h0014; B = 16'h00F7; #100;
A = 16'h0014; B = 16'h00F8; #100;
A = 16'h0014; B = 16'h00F9; #100;
A = 16'h0014; B = 16'h00FA; #100;
A = 16'h0014; B = 16'h00FB; #100;
A = 16'h0014; B = 16'h00FC; #100;
A = 16'h0014; B = 16'h00FD; #100;
A = 16'h0014; B = 16'h00FE; #100;
A = 16'h0014; B = 16'h00FF; #100;
A = 16'h0015; B = 16'h000; #100;
A = 16'h0015; B = 16'h001; #100;
A = 16'h0015; B = 16'h002; #100;
A = 16'h0015; B = 16'h003; #100;
A = 16'h0015; B = 16'h004; #100;
A = 16'h0015; B = 16'h005; #100;
A = 16'h0015; B = 16'h006; #100;
A = 16'h0015; B = 16'h007; #100;
A = 16'h0015; B = 16'h008; #100;
A = 16'h0015; B = 16'h009; #100;
A = 16'h0015; B = 16'h00A; #100;
A = 16'h0015; B = 16'h00B; #100;
A = 16'h0015; B = 16'h00C; #100;
A = 16'h0015; B = 16'h00D; #100;
A = 16'h0015; B = 16'h00E; #100;
A = 16'h0015; B = 16'h00F; #100;
A = 16'h0015; B = 16'h0010; #100;
A = 16'h0015; B = 16'h0011; #100;
A = 16'h0015; B = 16'h0012; #100;
A = 16'h0015; B = 16'h0013; #100;
A = 16'h0015; B = 16'h0014; #100;
A = 16'h0015; B = 16'h0015; #100;
A = 16'h0015; B = 16'h0016; #100;
A = 16'h0015; B = 16'h0017; #100;
A = 16'h0015; B = 16'h0018; #100;
A = 16'h0015; B = 16'h0019; #100;
A = 16'h0015; B = 16'h001A; #100;
A = 16'h0015; B = 16'h001B; #100;
A = 16'h0015; B = 16'h001C; #100;
A = 16'h0015; B = 16'h001D; #100;
A = 16'h0015; B = 16'h001E; #100;
A = 16'h0015; B = 16'h001F; #100;
A = 16'h0015; B = 16'h0020; #100;
A = 16'h0015; B = 16'h0021; #100;
A = 16'h0015; B = 16'h0022; #100;
A = 16'h0015; B = 16'h0023; #100;
A = 16'h0015; B = 16'h0024; #100;
A = 16'h0015; B = 16'h0025; #100;
A = 16'h0015; B = 16'h0026; #100;
A = 16'h0015; B = 16'h0027; #100;
A = 16'h0015; B = 16'h0028; #100;
A = 16'h0015; B = 16'h0029; #100;
A = 16'h0015; B = 16'h002A; #100;
A = 16'h0015; B = 16'h002B; #100;
A = 16'h0015; B = 16'h002C; #100;
A = 16'h0015; B = 16'h002D; #100;
A = 16'h0015; B = 16'h002E; #100;
A = 16'h0015; B = 16'h002F; #100;
A = 16'h0015; B = 16'h0030; #100;
A = 16'h0015; B = 16'h0031; #100;
A = 16'h0015; B = 16'h0032; #100;
A = 16'h0015; B = 16'h0033; #100;
A = 16'h0015; B = 16'h0034; #100;
A = 16'h0015; B = 16'h0035; #100;
A = 16'h0015; B = 16'h0036; #100;
A = 16'h0015; B = 16'h0037; #100;
A = 16'h0015; B = 16'h0038; #100;
A = 16'h0015; B = 16'h0039; #100;
A = 16'h0015; B = 16'h003A; #100;
A = 16'h0015; B = 16'h003B; #100;
A = 16'h0015; B = 16'h003C; #100;
A = 16'h0015; B = 16'h003D; #100;
A = 16'h0015; B = 16'h003E; #100;
A = 16'h0015; B = 16'h003F; #100;
A = 16'h0015; B = 16'h0040; #100;
A = 16'h0015; B = 16'h0041; #100;
A = 16'h0015; B = 16'h0042; #100;
A = 16'h0015; B = 16'h0043; #100;
A = 16'h0015; B = 16'h0044; #100;
A = 16'h0015; B = 16'h0045; #100;
A = 16'h0015; B = 16'h0046; #100;
A = 16'h0015; B = 16'h0047; #100;
A = 16'h0015; B = 16'h0048; #100;
A = 16'h0015; B = 16'h0049; #100;
A = 16'h0015; B = 16'h004A; #100;
A = 16'h0015; B = 16'h004B; #100;
A = 16'h0015; B = 16'h004C; #100;
A = 16'h0015; B = 16'h004D; #100;
A = 16'h0015; B = 16'h004E; #100;
A = 16'h0015; B = 16'h004F; #100;
A = 16'h0015; B = 16'h0050; #100;
A = 16'h0015; B = 16'h0051; #100;
A = 16'h0015; B = 16'h0052; #100;
A = 16'h0015; B = 16'h0053; #100;
A = 16'h0015; B = 16'h0054; #100;
A = 16'h0015; B = 16'h0055; #100;
A = 16'h0015; B = 16'h0056; #100;
A = 16'h0015; B = 16'h0057; #100;
A = 16'h0015; B = 16'h0058; #100;
A = 16'h0015; B = 16'h0059; #100;
A = 16'h0015; B = 16'h005A; #100;
A = 16'h0015; B = 16'h005B; #100;
A = 16'h0015; B = 16'h005C; #100;
A = 16'h0015; B = 16'h005D; #100;
A = 16'h0015; B = 16'h005E; #100;
A = 16'h0015; B = 16'h005F; #100;
A = 16'h0015; B = 16'h0060; #100;
A = 16'h0015; B = 16'h0061; #100;
A = 16'h0015; B = 16'h0062; #100;
A = 16'h0015; B = 16'h0063; #100;
A = 16'h0015; B = 16'h0064; #100;
A = 16'h0015; B = 16'h0065; #100;
A = 16'h0015; B = 16'h0066; #100;
A = 16'h0015; B = 16'h0067; #100;
A = 16'h0015; B = 16'h0068; #100;
A = 16'h0015; B = 16'h0069; #100;
A = 16'h0015; B = 16'h006A; #100;
A = 16'h0015; B = 16'h006B; #100;
A = 16'h0015; B = 16'h006C; #100;
A = 16'h0015; B = 16'h006D; #100;
A = 16'h0015; B = 16'h006E; #100;
A = 16'h0015; B = 16'h006F; #100;
A = 16'h0015; B = 16'h0070; #100;
A = 16'h0015; B = 16'h0071; #100;
A = 16'h0015; B = 16'h0072; #100;
A = 16'h0015; B = 16'h0073; #100;
A = 16'h0015; B = 16'h0074; #100;
A = 16'h0015; B = 16'h0075; #100;
A = 16'h0015; B = 16'h0076; #100;
A = 16'h0015; B = 16'h0077; #100;
A = 16'h0015; B = 16'h0078; #100;
A = 16'h0015; B = 16'h0079; #100;
A = 16'h0015; B = 16'h007A; #100;
A = 16'h0015; B = 16'h007B; #100;
A = 16'h0015; B = 16'h007C; #100;
A = 16'h0015; B = 16'h007D; #100;
A = 16'h0015; B = 16'h007E; #100;
A = 16'h0015; B = 16'h007F; #100;
A = 16'h0015; B = 16'h0080; #100;
A = 16'h0015; B = 16'h0081; #100;
A = 16'h0015; B = 16'h0082; #100;
A = 16'h0015; B = 16'h0083; #100;
A = 16'h0015; B = 16'h0084; #100;
A = 16'h0015; B = 16'h0085; #100;
A = 16'h0015; B = 16'h0086; #100;
A = 16'h0015; B = 16'h0087; #100;
A = 16'h0015; B = 16'h0088; #100;
A = 16'h0015; B = 16'h0089; #100;
A = 16'h0015; B = 16'h008A; #100;
A = 16'h0015; B = 16'h008B; #100;
A = 16'h0015; B = 16'h008C; #100;
A = 16'h0015; B = 16'h008D; #100;
A = 16'h0015; B = 16'h008E; #100;
A = 16'h0015; B = 16'h008F; #100;
A = 16'h0015; B = 16'h0090; #100;
A = 16'h0015; B = 16'h0091; #100;
A = 16'h0015; B = 16'h0092; #100;
A = 16'h0015; B = 16'h0093; #100;
A = 16'h0015; B = 16'h0094; #100;
A = 16'h0015; B = 16'h0095; #100;
A = 16'h0015; B = 16'h0096; #100;
A = 16'h0015; B = 16'h0097; #100;
A = 16'h0015; B = 16'h0098; #100;
A = 16'h0015; B = 16'h0099; #100;
A = 16'h0015; B = 16'h009A; #100;
A = 16'h0015; B = 16'h009B; #100;
A = 16'h0015; B = 16'h009C; #100;
A = 16'h0015; B = 16'h009D; #100;
A = 16'h0015; B = 16'h009E; #100;
A = 16'h0015; B = 16'h009F; #100;
A = 16'h0015; B = 16'h00A0; #100;
A = 16'h0015; B = 16'h00A1; #100;
A = 16'h0015; B = 16'h00A2; #100;
A = 16'h0015; B = 16'h00A3; #100;
A = 16'h0015; B = 16'h00A4; #100;
A = 16'h0015; B = 16'h00A5; #100;
A = 16'h0015; B = 16'h00A6; #100;
A = 16'h0015; B = 16'h00A7; #100;
A = 16'h0015; B = 16'h00A8; #100;
A = 16'h0015; B = 16'h00A9; #100;
A = 16'h0015; B = 16'h00AA; #100;
A = 16'h0015; B = 16'h00AB; #100;
A = 16'h0015; B = 16'h00AC; #100;
A = 16'h0015; B = 16'h00AD; #100;
A = 16'h0015; B = 16'h00AE; #100;
A = 16'h0015; B = 16'h00AF; #100;
A = 16'h0015; B = 16'h00B0; #100;
A = 16'h0015; B = 16'h00B1; #100;
A = 16'h0015; B = 16'h00B2; #100;
A = 16'h0015; B = 16'h00B3; #100;
A = 16'h0015; B = 16'h00B4; #100;
A = 16'h0015; B = 16'h00B5; #100;
A = 16'h0015; B = 16'h00B6; #100;
A = 16'h0015; B = 16'h00B7; #100;
A = 16'h0015; B = 16'h00B8; #100;
A = 16'h0015; B = 16'h00B9; #100;
A = 16'h0015; B = 16'h00BA; #100;
A = 16'h0015; B = 16'h00BB; #100;
A = 16'h0015; B = 16'h00BC; #100;
A = 16'h0015; B = 16'h00BD; #100;
A = 16'h0015; B = 16'h00BE; #100;
A = 16'h0015; B = 16'h00BF; #100;
A = 16'h0015; B = 16'h00C0; #100;
A = 16'h0015; B = 16'h00C1; #100;
A = 16'h0015; B = 16'h00C2; #100;
A = 16'h0015; B = 16'h00C3; #100;
A = 16'h0015; B = 16'h00C4; #100;
A = 16'h0015; B = 16'h00C5; #100;
A = 16'h0015; B = 16'h00C6; #100;
A = 16'h0015; B = 16'h00C7; #100;
A = 16'h0015; B = 16'h00C8; #100;
A = 16'h0015; B = 16'h00C9; #100;
A = 16'h0015; B = 16'h00CA; #100;
A = 16'h0015; B = 16'h00CB; #100;
A = 16'h0015; B = 16'h00CC; #100;
A = 16'h0015; B = 16'h00CD; #100;
A = 16'h0015; B = 16'h00CE; #100;
A = 16'h0015; B = 16'h00CF; #100;
A = 16'h0015; B = 16'h00D0; #100;
A = 16'h0015; B = 16'h00D1; #100;
A = 16'h0015; B = 16'h00D2; #100;
A = 16'h0015; B = 16'h00D3; #100;
A = 16'h0015; B = 16'h00D4; #100;
A = 16'h0015; B = 16'h00D5; #100;
A = 16'h0015; B = 16'h00D6; #100;
A = 16'h0015; B = 16'h00D7; #100;
A = 16'h0015; B = 16'h00D8; #100;
A = 16'h0015; B = 16'h00D9; #100;
A = 16'h0015; B = 16'h00DA; #100;
A = 16'h0015; B = 16'h00DB; #100;
A = 16'h0015; B = 16'h00DC; #100;
A = 16'h0015; B = 16'h00DD; #100;
A = 16'h0015; B = 16'h00DE; #100;
A = 16'h0015; B = 16'h00DF; #100;
A = 16'h0015; B = 16'h00E0; #100;
A = 16'h0015; B = 16'h00E1; #100;
A = 16'h0015; B = 16'h00E2; #100;
A = 16'h0015; B = 16'h00E3; #100;
A = 16'h0015; B = 16'h00E4; #100;
A = 16'h0015; B = 16'h00E5; #100;
A = 16'h0015; B = 16'h00E6; #100;
A = 16'h0015; B = 16'h00E7; #100;
A = 16'h0015; B = 16'h00E8; #100;
A = 16'h0015; B = 16'h00E9; #100;
A = 16'h0015; B = 16'h00EA; #100;
A = 16'h0015; B = 16'h00EB; #100;
A = 16'h0015; B = 16'h00EC; #100;
A = 16'h0015; B = 16'h00ED; #100;
A = 16'h0015; B = 16'h00EE; #100;
A = 16'h0015; B = 16'h00EF; #100;
A = 16'h0015; B = 16'h00F0; #100;
A = 16'h0015; B = 16'h00F1; #100;
A = 16'h0015; B = 16'h00F2; #100;
A = 16'h0015; B = 16'h00F3; #100;
A = 16'h0015; B = 16'h00F4; #100;
A = 16'h0015; B = 16'h00F5; #100;
A = 16'h0015; B = 16'h00F6; #100;
A = 16'h0015; B = 16'h00F7; #100;
A = 16'h0015; B = 16'h00F8; #100;
A = 16'h0015; B = 16'h00F9; #100;
A = 16'h0015; B = 16'h00FA; #100;
A = 16'h0015; B = 16'h00FB; #100;
A = 16'h0015; B = 16'h00FC; #100;
A = 16'h0015; B = 16'h00FD; #100;
A = 16'h0015; B = 16'h00FE; #100;
A = 16'h0015; B = 16'h00FF; #100;
A = 16'h0016; B = 16'h000; #100;
A = 16'h0016; B = 16'h001; #100;
A = 16'h0016; B = 16'h002; #100;
A = 16'h0016; B = 16'h003; #100;
A = 16'h0016; B = 16'h004; #100;
A = 16'h0016; B = 16'h005; #100;
A = 16'h0016; B = 16'h006; #100;
A = 16'h0016; B = 16'h007; #100;
A = 16'h0016; B = 16'h008; #100;
A = 16'h0016; B = 16'h009; #100;
A = 16'h0016; B = 16'h00A; #100;
A = 16'h0016; B = 16'h00B; #100;
A = 16'h0016; B = 16'h00C; #100;
A = 16'h0016; B = 16'h00D; #100;
A = 16'h0016; B = 16'h00E; #100;
A = 16'h0016; B = 16'h00F; #100;
A = 16'h0016; B = 16'h0010; #100;
A = 16'h0016; B = 16'h0011; #100;
A = 16'h0016; B = 16'h0012; #100;
A = 16'h0016; B = 16'h0013; #100;
A = 16'h0016; B = 16'h0014; #100;
A = 16'h0016; B = 16'h0015; #100;
A = 16'h0016; B = 16'h0016; #100;
A = 16'h0016; B = 16'h0017; #100;
A = 16'h0016; B = 16'h0018; #100;
A = 16'h0016; B = 16'h0019; #100;
A = 16'h0016; B = 16'h001A; #100;
A = 16'h0016; B = 16'h001B; #100;
A = 16'h0016; B = 16'h001C; #100;
A = 16'h0016; B = 16'h001D; #100;
A = 16'h0016; B = 16'h001E; #100;
A = 16'h0016; B = 16'h001F; #100;
A = 16'h0016; B = 16'h0020; #100;
A = 16'h0016; B = 16'h0021; #100;
A = 16'h0016; B = 16'h0022; #100;
A = 16'h0016; B = 16'h0023; #100;
A = 16'h0016; B = 16'h0024; #100;
A = 16'h0016; B = 16'h0025; #100;
A = 16'h0016; B = 16'h0026; #100;
A = 16'h0016; B = 16'h0027; #100;
A = 16'h0016; B = 16'h0028; #100;
A = 16'h0016; B = 16'h0029; #100;
A = 16'h0016; B = 16'h002A; #100;
A = 16'h0016; B = 16'h002B; #100;
A = 16'h0016; B = 16'h002C; #100;
A = 16'h0016; B = 16'h002D; #100;
A = 16'h0016; B = 16'h002E; #100;
A = 16'h0016; B = 16'h002F; #100;
A = 16'h0016; B = 16'h0030; #100;
A = 16'h0016; B = 16'h0031; #100;
A = 16'h0016; B = 16'h0032; #100;
A = 16'h0016; B = 16'h0033; #100;
A = 16'h0016; B = 16'h0034; #100;
A = 16'h0016; B = 16'h0035; #100;
A = 16'h0016; B = 16'h0036; #100;
A = 16'h0016; B = 16'h0037; #100;
A = 16'h0016; B = 16'h0038; #100;
A = 16'h0016; B = 16'h0039; #100;
A = 16'h0016; B = 16'h003A; #100;
A = 16'h0016; B = 16'h003B; #100;
A = 16'h0016; B = 16'h003C; #100;
A = 16'h0016; B = 16'h003D; #100;
A = 16'h0016; B = 16'h003E; #100;
A = 16'h0016; B = 16'h003F; #100;
A = 16'h0016; B = 16'h0040; #100;
A = 16'h0016; B = 16'h0041; #100;
A = 16'h0016; B = 16'h0042; #100;
A = 16'h0016; B = 16'h0043; #100;
A = 16'h0016; B = 16'h0044; #100;
A = 16'h0016; B = 16'h0045; #100;
A = 16'h0016; B = 16'h0046; #100;
A = 16'h0016; B = 16'h0047; #100;
A = 16'h0016; B = 16'h0048; #100;
A = 16'h0016; B = 16'h0049; #100;
A = 16'h0016; B = 16'h004A; #100;
A = 16'h0016; B = 16'h004B; #100;
A = 16'h0016; B = 16'h004C; #100;
A = 16'h0016; B = 16'h004D; #100;
A = 16'h0016; B = 16'h004E; #100;
A = 16'h0016; B = 16'h004F; #100;
A = 16'h0016; B = 16'h0050; #100;
A = 16'h0016; B = 16'h0051; #100;
A = 16'h0016; B = 16'h0052; #100;
A = 16'h0016; B = 16'h0053; #100;
A = 16'h0016; B = 16'h0054; #100;
A = 16'h0016; B = 16'h0055; #100;
A = 16'h0016; B = 16'h0056; #100;
A = 16'h0016; B = 16'h0057; #100;
A = 16'h0016; B = 16'h0058; #100;
A = 16'h0016; B = 16'h0059; #100;
A = 16'h0016; B = 16'h005A; #100;
A = 16'h0016; B = 16'h005B; #100;
A = 16'h0016; B = 16'h005C; #100;
A = 16'h0016; B = 16'h005D; #100;
A = 16'h0016; B = 16'h005E; #100;
A = 16'h0016; B = 16'h005F; #100;
A = 16'h0016; B = 16'h0060; #100;
A = 16'h0016; B = 16'h0061; #100;
A = 16'h0016; B = 16'h0062; #100;
A = 16'h0016; B = 16'h0063; #100;
A = 16'h0016; B = 16'h0064; #100;
A = 16'h0016; B = 16'h0065; #100;
A = 16'h0016; B = 16'h0066; #100;
A = 16'h0016; B = 16'h0067; #100;
A = 16'h0016; B = 16'h0068; #100;
A = 16'h0016; B = 16'h0069; #100;
A = 16'h0016; B = 16'h006A; #100;
A = 16'h0016; B = 16'h006B; #100;
A = 16'h0016; B = 16'h006C; #100;
A = 16'h0016; B = 16'h006D; #100;
A = 16'h0016; B = 16'h006E; #100;
A = 16'h0016; B = 16'h006F; #100;
A = 16'h0016; B = 16'h0070; #100;
A = 16'h0016; B = 16'h0071; #100;
A = 16'h0016; B = 16'h0072; #100;
A = 16'h0016; B = 16'h0073; #100;
A = 16'h0016; B = 16'h0074; #100;
A = 16'h0016; B = 16'h0075; #100;
A = 16'h0016; B = 16'h0076; #100;
A = 16'h0016; B = 16'h0077; #100;
A = 16'h0016; B = 16'h0078; #100;
A = 16'h0016; B = 16'h0079; #100;
A = 16'h0016; B = 16'h007A; #100;
A = 16'h0016; B = 16'h007B; #100;
A = 16'h0016; B = 16'h007C; #100;
A = 16'h0016; B = 16'h007D; #100;
A = 16'h0016; B = 16'h007E; #100;
A = 16'h0016; B = 16'h007F; #100;
A = 16'h0016; B = 16'h0080; #100;
A = 16'h0016; B = 16'h0081; #100;
A = 16'h0016; B = 16'h0082; #100;
A = 16'h0016; B = 16'h0083; #100;
A = 16'h0016; B = 16'h0084; #100;
A = 16'h0016; B = 16'h0085; #100;
A = 16'h0016; B = 16'h0086; #100;
A = 16'h0016; B = 16'h0087; #100;
A = 16'h0016; B = 16'h0088; #100;
A = 16'h0016; B = 16'h0089; #100;
A = 16'h0016; B = 16'h008A; #100;
A = 16'h0016; B = 16'h008B; #100;
A = 16'h0016; B = 16'h008C; #100;
A = 16'h0016; B = 16'h008D; #100;
A = 16'h0016; B = 16'h008E; #100;
A = 16'h0016; B = 16'h008F; #100;
A = 16'h0016; B = 16'h0090; #100;
A = 16'h0016; B = 16'h0091; #100;
A = 16'h0016; B = 16'h0092; #100;
A = 16'h0016; B = 16'h0093; #100;
A = 16'h0016; B = 16'h0094; #100;
A = 16'h0016; B = 16'h0095; #100;
A = 16'h0016; B = 16'h0096; #100;
A = 16'h0016; B = 16'h0097; #100;
A = 16'h0016; B = 16'h0098; #100;
A = 16'h0016; B = 16'h0099; #100;
A = 16'h0016; B = 16'h009A; #100;
A = 16'h0016; B = 16'h009B; #100;
A = 16'h0016; B = 16'h009C; #100;
A = 16'h0016; B = 16'h009D; #100;
A = 16'h0016; B = 16'h009E; #100;
A = 16'h0016; B = 16'h009F; #100;
A = 16'h0016; B = 16'h00A0; #100;
A = 16'h0016; B = 16'h00A1; #100;
A = 16'h0016; B = 16'h00A2; #100;
A = 16'h0016; B = 16'h00A3; #100;
A = 16'h0016; B = 16'h00A4; #100;
A = 16'h0016; B = 16'h00A5; #100;
A = 16'h0016; B = 16'h00A6; #100;
A = 16'h0016; B = 16'h00A7; #100;
A = 16'h0016; B = 16'h00A8; #100;
A = 16'h0016; B = 16'h00A9; #100;
A = 16'h0016; B = 16'h00AA; #100;
A = 16'h0016; B = 16'h00AB; #100;
A = 16'h0016; B = 16'h00AC; #100;
A = 16'h0016; B = 16'h00AD; #100;
A = 16'h0016; B = 16'h00AE; #100;
A = 16'h0016; B = 16'h00AF; #100;
A = 16'h0016; B = 16'h00B0; #100;
A = 16'h0016; B = 16'h00B1; #100;
A = 16'h0016; B = 16'h00B2; #100;
A = 16'h0016; B = 16'h00B3; #100;
A = 16'h0016; B = 16'h00B4; #100;
A = 16'h0016; B = 16'h00B5; #100;
A = 16'h0016; B = 16'h00B6; #100;
A = 16'h0016; B = 16'h00B7; #100;
A = 16'h0016; B = 16'h00B8; #100;
A = 16'h0016; B = 16'h00B9; #100;
A = 16'h0016; B = 16'h00BA; #100;
A = 16'h0016; B = 16'h00BB; #100;
A = 16'h0016; B = 16'h00BC; #100;
A = 16'h0016; B = 16'h00BD; #100;
A = 16'h0016; B = 16'h00BE; #100;
A = 16'h0016; B = 16'h00BF; #100;
A = 16'h0016; B = 16'h00C0; #100;
A = 16'h0016; B = 16'h00C1; #100;
A = 16'h0016; B = 16'h00C2; #100;
A = 16'h0016; B = 16'h00C3; #100;
A = 16'h0016; B = 16'h00C4; #100;
A = 16'h0016; B = 16'h00C5; #100;
A = 16'h0016; B = 16'h00C6; #100;
A = 16'h0016; B = 16'h00C7; #100;
A = 16'h0016; B = 16'h00C8; #100;
A = 16'h0016; B = 16'h00C9; #100;
A = 16'h0016; B = 16'h00CA; #100;
A = 16'h0016; B = 16'h00CB; #100;
A = 16'h0016; B = 16'h00CC; #100;
A = 16'h0016; B = 16'h00CD; #100;
A = 16'h0016; B = 16'h00CE; #100;
A = 16'h0016; B = 16'h00CF; #100;
A = 16'h0016; B = 16'h00D0; #100;
A = 16'h0016; B = 16'h00D1; #100;
A = 16'h0016; B = 16'h00D2; #100;
A = 16'h0016; B = 16'h00D3; #100;
A = 16'h0016; B = 16'h00D4; #100;
A = 16'h0016; B = 16'h00D5; #100;
A = 16'h0016; B = 16'h00D6; #100;
A = 16'h0016; B = 16'h00D7; #100;
A = 16'h0016; B = 16'h00D8; #100;
A = 16'h0016; B = 16'h00D9; #100;
A = 16'h0016; B = 16'h00DA; #100;
A = 16'h0016; B = 16'h00DB; #100;
A = 16'h0016; B = 16'h00DC; #100;
A = 16'h0016; B = 16'h00DD; #100;
A = 16'h0016; B = 16'h00DE; #100;
A = 16'h0016; B = 16'h00DF; #100;
A = 16'h0016; B = 16'h00E0; #100;
A = 16'h0016; B = 16'h00E1; #100;
A = 16'h0016; B = 16'h00E2; #100;
A = 16'h0016; B = 16'h00E3; #100;
A = 16'h0016; B = 16'h00E4; #100;
A = 16'h0016; B = 16'h00E5; #100;
A = 16'h0016; B = 16'h00E6; #100;
A = 16'h0016; B = 16'h00E7; #100;
A = 16'h0016; B = 16'h00E8; #100;
A = 16'h0016; B = 16'h00E9; #100;
A = 16'h0016; B = 16'h00EA; #100;
A = 16'h0016; B = 16'h00EB; #100;
A = 16'h0016; B = 16'h00EC; #100;
A = 16'h0016; B = 16'h00ED; #100;
A = 16'h0016; B = 16'h00EE; #100;
A = 16'h0016; B = 16'h00EF; #100;
A = 16'h0016; B = 16'h00F0; #100;
A = 16'h0016; B = 16'h00F1; #100;
A = 16'h0016; B = 16'h00F2; #100;
A = 16'h0016; B = 16'h00F3; #100;
A = 16'h0016; B = 16'h00F4; #100;
A = 16'h0016; B = 16'h00F5; #100;
A = 16'h0016; B = 16'h00F6; #100;
A = 16'h0016; B = 16'h00F7; #100;
A = 16'h0016; B = 16'h00F8; #100;
A = 16'h0016; B = 16'h00F9; #100;
A = 16'h0016; B = 16'h00FA; #100;
A = 16'h0016; B = 16'h00FB; #100;
A = 16'h0016; B = 16'h00FC; #100;
A = 16'h0016; B = 16'h00FD; #100;
A = 16'h0016; B = 16'h00FE; #100;
A = 16'h0016; B = 16'h00FF; #100;
A = 16'h0017; B = 16'h000; #100;
A = 16'h0017; B = 16'h001; #100;
A = 16'h0017; B = 16'h002; #100;
A = 16'h0017; B = 16'h003; #100;
A = 16'h0017; B = 16'h004; #100;
A = 16'h0017; B = 16'h005; #100;
A = 16'h0017; B = 16'h006; #100;
A = 16'h0017; B = 16'h007; #100;
A = 16'h0017; B = 16'h008; #100;
A = 16'h0017; B = 16'h009; #100;
A = 16'h0017; B = 16'h00A; #100;
A = 16'h0017; B = 16'h00B; #100;
A = 16'h0017; B = 16'h00C; #100;
A = 16'h0017; B = 16'h00D; #100;
A = 16'h0017; B = 16'h00E; #100;
A = 16'h0017; B = 16'h00F; #100;
A = 16'h0017; B = 16'h0010; #100;
A = 16'h0017; B = 16'h0011; #100;
A = 16'h0017; B = 16'h0012; #100;
A = 16'h0017; B = 16'h0013; #100;
A = 16'h0017; B = 16'h0014; #100;
A = 16'h0017; B = 16'h0015; #100;
A = 16'h0017; B = 16'h0016; #100;
A = 16'h0017; B = 16'h0017; #100;
A = 16'h0017; B = 16'h0018; #100;
A = 16'h0017; B = 16'h0019; #100;
A = 16'h0017; B = 16'h001A; #100;
A = 16'h0017; B = 16'h001B; #100;
A = 16'h0017; B = 16'h001C; #100;
A = 16'h0017; B = 16'h001D; #100;
A = 16'h0017; B = 16'h001E; #100;
A = 16'h0017; B = 16'h001F; #100;
A = 16'h0017; B = 16'h0020; #100;
A = 16'h0017; B = 16'h0021; #100;
A = 16'h0017; B = 16'h0022; #100;
A = 16'h0017; B = 16'h0023; #100;
A = 16'h0017; B = 16'h0024; #100;
A = 16'h0017; B = 16'h0025; #100;
A = 16'h0017; B = 16'h0026; #100;
A = 16'h0017; B = 16'h0027; #100;
A = 16'h0017; B = 16'h0028; #100;
A = 16'h0017; B = 16'h0029; #100;
A = 16'h0017; B = 16'h002A; #100;
A = 16'h0017; B = 16'h002B; #100;
A = 16'h0017; B = 16'h002C; #100;
A = 16'h0017; B = 16'h002D; #100;
A = 16'h0017; B = 16'h002E; #100;
A = 16'h0017; B = 16'h002F; #100;
A = 16'h0017; B = 16'h0030; #100;
A = 16'h0017; B = 16'h0031; #100;
A = 16'h0017; B = 16'h0032; #100;
A = 16'h0017; B = 16'h0033; #100;
A = 16'h0017; B = 16'h0034; #100;
A = 16'h0017; B = 16'h0035; #100;
A = 16'h0017; B = 16'h0036; #100;
A = 16'h0017; B = 16'h0037; #100;
A = 16'h0017; B = 16'h0038; #100;
A = 16'h0017; B = 16'h0039; #100;
A = 16'h0017; B = 16'h003A; #100;
A = 16'h0017; B = 16'h003B; #100;
A = 16'h0017; B = 16'h003C; #100;
A = 16'h0017; B = 16'h003D; #100;
A = 16'h0017; B = 16'h003E; #100;
A = 16'h0017; B = 16'h003F; #100;
A = 16'h0017; B = 16'h0040; #100;
A = 16'h0017; B = 16'h0041; #100;
A = 16'h0017; B = 16'h0042; #100;
A = 16'h0017; B = 16'h0043; #100;
A = 16'h0017; B = 16'h0044; #100;
A = 16'h0017; B = 16'h0045; #100;
A = 16'h0017; B = 16'h0046; #100;
A = 16'h0017; B = 16'h0047; #100;
A = 16'h0017; B = 16'h0048; #100;
A = 16'h0017; B = 16'h0049; #100;
A = 16'h0017; B = 16'h004A; #100;
A = 16'h0017; B = 16'h004B; #100;
A = 16'h0017; B = 16'h004C; #100;
A = 16'h0017; B = 16'h004D; #100;
A = 16'h0017; B = 16'h004E; #100;
A = 16'h0017; B = 16'h004F; #100;
A = 16'h0017; B = 16'h0050; #100;
A = 16'h0017; B = 16'h0051; #100;
A = 16'h0017; B = 16'h0052; #100;
A = 16'h0017; B = 16'h0053; #100;
A = 16'h0017; B = 16'h0054; #100;
A = 16'h0017; B = 16'h0055; #100;
A = 16'h0017; B = 16'h0056; #100;
A = 16'h0017; B = 16'h0057; #100;
A = 16'h0017; B = 16'h0058; #100;
A = 16'h0017; B = 16'h0059; #100;
A = 16'h0017; B = 16'h005A; #100;
A = 16'h0017; B = 16'h005B; #100;
A = 16'h0017; B = 16'h005C; #100;
A = 16'h0017; B = 16'h005D; #100;
A = 16'h0017; B = 16'h005E; #100;
A = 16'h0017; B = 16'h005F; #100;
A = 16'h0017; B = 16'h0060; #100;
A = 16'h0017; B = 16'h0061; #100;
A = 16'h0017; B = 16'h0062; #100;
A = 16'h0017; B = 16'h0063; #100;
A = 16'h0017; B = 16'h0064; #100;
A = 16'h0017; B = 16'h0065; #100;
A = 16'h0017; B = 16'h0066; #100;
A = 16'h0017; B = 16'h0067; #100;
A = 16'h0017; B = 16'h0068; #100;
A = 16'h0017; B = 16'h0069; #100;
A = 16'h0017; B = 16'h006A; #100;
A = 16'h0017; B = 16'h006B; #100;
A = 16'h0017; B = 16'h006C; #100;
A = 16'h0017; B = 16'h006D; #100;
A = 16'h0017; B = 16'h006E; #100;
A = 16'h0017; B = 16'h006F; #100;
A = 16'h0017; B = 16'h0070; #100;
A = 16'h0017; B = 16'h0071; #100;
A = 16'h0017; B = 16'h0072; #100;
A = 16'h0017; B = 16'h0073; #100;
A = 16'h0017; B = 16'h0074; #100;
A = 16'h0017; B = 16'h0075; #100;
A = 16'h0017; B = 16'h0076; #100;
A = 16'h0017; B = 16'h0077; #100;
A = 16'h0017; B = 16'h0078; #100;
A = 16'h0017; B = 16'h0079; #100;
A = 16'h0017; B = 16'h007A; #100;
A = 16'h0017; B = 16'h007B; #100;
A = 16'h0017; B = 16'h007C; #100;
A = 16'h0017; B = 16'h007D; #100;
A = 16'h0017; B = 16'h007E; #100;
A = 16'h0017; B = 16'h007F; #100;
A = 16'h0017; B = 16'h0080; #100;
A = 16'h0017; B = 16'h0081; #100;
A = 16'h0017; B = 16'h0082; #100;
A = 16'h0017; B = 16'h0083; #100;
A = 16'h0017; B = 16'h0084; #100;
A = 16'h0017; B = 16'h0085; #100;
A = 16'h0017; B = 16'h0086; #100;
A = 16'h0017; B = 16'h0087; #100;
A = 16'h0017; B = 16'h0088; #100;
A = 16'h0017; B = 16'h0089; #100;
A = 16'h0017; B = 16'h008A; #100;
A = 16'h0017; B = 16'h008B; #100;
A = 16'h0017; B = 16'h008C; #100;
A = 16'h0017; B = 16'h008D; #100;
A = 16'h0017; B = 16'h008E; #100;
A = 16'h0017; B = 16'h008F; #100;
A = 16'h0017; B = 16'h0090; #100;
A = 16'h0017; B = 16'h0091; #100;
A = 16'h0017; B = 16'h0092; #100;
A = 16'h0017; B = 16'h0093; #100;
A = 16'h0017; B = 16'h0094; #100;
A = 16'h0017; B = 16'h0095; #100;
A = 16'h0017; B = 16'h0096; #100;
A = 16'h0017; B = 16'h0097; #100;
A = 16'h0017; B = 16'h0098; #100;
A = 16'h0017; B = 16'h0099; #100;
A = 16'h0017; B = 16'h009A; #100;
A = 16'h0017; B = 16'h009B; #100;
A = 16'h0017; B = 16'h009C; #100;
A = 16'h0017; B = 16'h009D; #100;
A = 16'h0017; B = 16'h009E; #100;
A = 16'h0017; B = 16'h009F; #100;
A = 16'h0017; B = 16'h00A0; #100;
A = 16'h0017; B = 16'h00A1; #100;
A = 16'h0017; B = 16'h00A2; #100;
A = 16'h0017; B = 16'h00A3; #100;
A = 16'h0017; B = 16'h00A4; #100;
A = 16'h0017; B = 16'h00A5; #100;
A = 16'h0017; B = 16'h00A6; #100;
A = 16'h0017; B = 16'h00A7; #100;
A = 16'h0017; B = 16'h00A8; #100;
A = 16'h0017; B = 16'h00A9; #100;
A = 16'h0017; B = 16'h00AA; #100;
A = 16'h0017; B = 16'h00AB; #100;
A = 16'h0017; B = 16'h00AC; #100;
A = 16'h0017; B = 16'h00AD; #100;
A = 16'h0017; B = 16'h00AE; #100;
A = 16'h0017; B = 16'h00AF; #100;
A = 16'h0017; B = 16'h00B0; #100;
A = 16'h0017; B = 16'h00B1; #100;
A = 16'h0017; B = 16'h00B2; #100;
A = 16'h0017; B = 16'h00B3; #100;
A = 16'h0017; B = 16'h00B4; #100;
A = 16'h0017; B = 16'h00B5; #100;
A = 16'h0017; B = 16'h00B6; #100;
A = 16'h0017; B = 16'h00B7; #100;
A = 16'h0017; B = 16'h00B8; #100;
A = 16'h0017; B = 16'h00B9; #100;
A = 16'h0017; B = 16'h00BA; #100;
A = 16'h0017; B = 16'h00BB; #100;
A = 16'h0017; B = 16'h00BC; #100;
A = 16'h0017; B = 16'h00BD; #100;
A = 16'h0017; B = 16'h00BE; #100;
A = 16'h0017; B = 16'h00BF; #100;
A = 16'h0017; B = 16'h00C0; #100;
A = 16'h0017; B = 16'h00C1; #100;
A = 16'h0017; B = 16'h00C2; #100;
A = 16'h0017; B = 16'h00C3; #100;
A = 16'h0017; B = 16'h00C4; #100;
A = 16'h0017; B = 16'h00C5; #100;
A = 16'h0017; B = 16'h00C6; #100;
A = 16'h0017; B = 16'h00C7; #100;
A = 16'h0017; B = 16'h00C8; #100;
A = 16'h0017; B = 16'h00C9; #100;
A = 16'h0017; B = 16'h00CA; #100;
A = 16'h0017; B = 16'h00CB; #100;
A = 16'h0017; B = 16'h00CC; #100;
A = 16'h0017; B = 16'h00CD; #100;
A = 16'h0017; B = 16'h00CE; #100;
A = 16'h0017; B = 16'h00CF; #100;
A = 16'h0017; B = 16'h00D0; #100;
A = 16'h0017; B = 16'h00D1; #100;
A = 16'h0017; B = 16'h00D2; #100;
A = 16'h0017; B = 16'h00D3; #100;
A = 16'h0017; B = 16'h00D4; #100;
A = 16'h0017; B = 16'h00D5; #100;
A = 16'h0017; B = 16'h00D6; #100;
A = 16'h0017; B = 16'h00D7; #100;
A = 16'h0017; B = 16'h00D8; #100;
A = 16'h0017; B = 16'h00D9; #100;
A = 16'h0017; B = 16'h00DA; #100;
A = 16'h0017; B = 16'h00DB; #100;
A = 16'h0017; B = 16'h00DC; #100;
A = 16'h0017; B = 16'h00DD; #100;
A = 16'h0017; B = 16'h00DE; #100;
A = 16'h0017; B = 16'h00DF; #100;
A = 16'h0017; B = 16'h00E0; #100;
A = 16'h0017; B = 16'h00E1; #100;
A = 16'h0017; B = 16'h00E2; #100;
A = 16'h0017; B = 16'h00E3; #100;
A = 16'h0017; B = 16'h00E4; #100;
A = 16'h0017; B = 16'h00E5; #100;
A = 16'h0017; B = 16'h00E6; #100;
A = 16'h0017; B = 16'h00E7; #100;
A = 16'h0017; B = 16'h00E8; #100;
A = 16'h0017; B = 16'h00E9; #100;
A = 16'h0017; B = 16'h00EA; #100;
A = 16'h0017; B = 16'h00EB; #100;
A = 16'h0017; B = 16'h00EC; #100;
A = 16'h0017; B = 16'h00ED; #100;
A = 16'h0017; B = 16'h00EE; #100;
A = 16'h0017; B = 16'h00EF; #100;
A = 16'h0017; B = 16'h00F0; #100;
A = 16'h0017; B = 16'h00F1; #100;
A = 16'h0017; B = 16'h00F2; #100;
A = 16'h0017; B = 16'h00F3; #100;
A = 16'h0017; B = 16'h00F4; #100;
A = 16'h0017; B = 16'h00F5; #100;
A = 16'h0017; B = 16'h00F6; #100;
A = 16'h0017; B = 16'h00F7; #100;
A = 16'h0017; B = 16'h00F8; #100;
A = 16'h0017; B = 16'h00F9; #100;
A = 16'h0017; B = 16'h00FA; #100;
A = 16'h0017; B = 16'h00FB; #100;
A = 16'h0017; B = 16'h00FC; #100;
A = 16'h0017; B = 16'h00FD; #100;
A = 16'h0017; B = 16'h00FE; #100;
A = 16'h0017; B = 16'h00FF; #100;
A = 16'h0018; B = 16'h000; #100;
A = 16'h0018; B = 16'h001; #100;
A = 16'h0018; B = 16'h002; #100;
A = 16'h0018; B = 16'h003; #100;
A = 16'h0018; B = 16'h004; #100;
A = 16'h0018; B = 16'h005; #100;
A = 16'h0018; B = 16'h006; #100;
A = 16'h0018; B = 16'h007; #100;
A = 16'h0018; B = 16'h008; #100;
A = 16'h0018; B = 16'h009; #100;
A = 16'h0018; B = 16'h00A; #100;
A = 16'h0018; B = 16'h00B; #100;
A = 16'h0018; B = 16'h00C; #100;
A = 16'h0018; B = 16'h00D; #100;
A = 16'h0018; B = 16'h00E; #100;
A = 16'h0018; B = 16'h00F; #100;
A = 16'h0018; B = 16'h0010; #100;
A = 16'h0018; B = 16'h0011; #100;
A = 16'h0018; B = 16'h0012; #100;
A = 16'h0018; B = 16'h0013; #100;
A = 16'h0018; B = 16'h0014; #100;
A = 16'h0018; B = 16'h0015; #100;
A = 16'h0018; B = 16'h0016; #100;
A = 16'h0018; B = 16'h0017; #100;
A = 16'h0018; B = 16'h0018; #100;
A = 16'h0018; B = 16'h0019; #100;
A = 16'h0018; B = 16'h001A; #100;
A = 16'h0018; B = 16'h001B; #100;
A = 16'h0018; B = 16'h001C; #100;
A = 16'h0018; B = 16'h001D; #100;
A = 16'h0018; B = 16'h001E; #100;
A = 16'h0018; B = 16'h001F; #100;
A = 16'h0018; B = 16'h0020; #100;
A = 16'h0018; B = 16'h0021; #100;
A = 16'h0018; B = 16'h0022; #100;
A = 16'h0018; B = 16'h0023; #100;
A = 16'h0018; B = 16'h0024; #100;
A = 16'h0018; B = 16'h0025; #100;
A = 16'h0018; B = 16'h0026; #100;
A = 16'h0018; B = 16'h0027; #100;
A = 16'h0018; B = 16'h0028; #100;
A = 16'h0018; B = 16'h0029; #100;
A = 16'h0018; B = 16'h002A; #100;
A = 16'h0018; B = 16'h002B; #100;
A = 16'h0018; B = 16'h002C; #100;
A = 16'h0018; B = 16'h002D; #100;
A = 16'h0018; B = 16'h002E; #100;
A = 16'h0018; B = 16'h002F; #100;
A = 16'h0018; B = 16'h0030; #100;
A = 16'h0018; B = 16'h0031; #100;
A = 16'h0018; B = 16'h0032; #100;
A = 16'h0018; B = 16'h0033; #100;
A = 16'h0018; B = 16'h0034; #100;
A = 16'h0018; B = 16'h0035; #100;
A = 16'h0018; B = 16'h0036; #100;
A = 16'h0018; B = 16'h0037; #100;
A = 16'h0018; B = 16'h0038; #100;
A = 16'h0018; B = 16'h0039; #100;
A = 16'h0018; B = 16'h003A; #100;
A = 16'h0018; B = 16'h003B; #100;
A = 16'h0018; B = 16'h003C; #100;
A = 16'h0018; B = 16'h003D; #100;
A = 16'h0018; B = 16'h003E; #100;
A = 16'h0018; B = 16'h003F; #100;
A = 16'h0018; B = 16'h0040; #100;
A = 16'h0018; B = 16'h0041; #100;
A = 16'h0018; B = 16'h0042; #100;
A = 16'h0018; B = 16'h0043; #100;
A = 16'h0018; B = 16'h0044; #100;
A = 16'h0018; B = 16'h0045; #100;
A = 16'h0018; B = 16'h0046; #100;
A = 16'h0018; B = 16'h0047; #100;
A = 16'h0018; B = 16'h0048; #100;
A = 16'h0018; B = 16'h0049; #100;
A = 16'h0018; B = 16'h004A; #100;
A = 16'h0018; B = 16'h004B; #100;
A = 16'h0018; B = 16'h004C; #100;
A = 16'h0018; B = 16'h004D; #100;
A = 16'h0018; B = 16'h004E; #100;
A = 16'h0018; B = 16'h004F; #100;
A = 16'h0018; B = 16'h0050; #100;
A = 16'h0018; B = 16'h0051; #100;
A = 16'h0018; B = 16'h0052; #100;
A = 16'h0018; B = 16'h0053; #100;
A = 16'h0018; B = 16'h0054; #100;
A = 16'h0018; B = 16'h0055; #100;
A = 16'h0018; B = 16'h0056; #100;
A = 16'h0018; B = 16'h0057; #100;
A = 16'h0018; B = 16'h0058; #100;
A = 16'h0018; B = 16'h0059; #100;
A = 16'h0018; B = 16'h005A; #100;
A = 16'h0018; B = 16'h005B; #100;
A = 16'h0018; B = 16'h005C; #100;
A = 16'h0018; B = 16'h005D; #100;
A = 16'h0018; B = 16'h005E; #100;
A = 16'h0018; B = 16'h005F; #100;
A = 16'h0018; B = 16'h0060; #100;
A = 16'h0018; B = 16'h0061; #100;
A = 16'h0018; B = 16'h0062; #100;
A = 16'h0018; B = 16'h0063; #100;
A = 16'h0018; B = 16'h0064; #100;
A = 16'h0018; B = 16'h0065; #100;
A = 16'h0018; B = 16'h0066; #100;
A = 16'h0018; B = 16'h0067; #100;
A = 16'h0018; B = 16'h0068; #100;
A = 16'h0018; B = 16'h0069; #100;
A = 16'h0018; B = 16'h006A; #100;
A = 16'h0018; B = 16'h006B; #100;
A = 16'h0018; B = 16'h006C; #100;
A = 16'h0018; B = 16'h006D; #100;
A = 16'h0018; B = 16'h006E; #100;
A = 16'h0018; B = 16'h006F; #100;
A = 16'h0018; B = 16'h0070; #100;
A = 16'h0018; B = 16'h0071; #100;
A = 16'h0018; B = 16'h0072; #100;
A = 16'h0018; B = 16'h0073; #100;
A = 16'h0018; B = 16'h0074; #100;
A = 16'h0018; B = 16'h0075; #100;
A = 16'h0018; B = 16'h0076; #100;
A = 16'h0018; B = 16'h0077; #100;
A = 16'h0018; B = 16'h0078; #100;
A = 16'h0018; B = 16'h0079; #100;
A = 16'h0018; B = 16'h007A; #100;
A = 16'h0018; B = 16'h007B; #100;
A = 16'h0018; B = 16'h007C; #100;
A = 16'h0018; B = 16'h007D; #100;
A = 16'h0018; B = 16'h007E; #100;
A = 16'h0018; B = 16'h007F; #100;
A = 16'h0018; B = 16'h0080; #100;
A = 16'h0018; B = 16'h0081; #100;
A = 16'h0018; B = 16'h0082; #100;
A = 16'h0018; B = 16'h0083; #100;
A = 16'h0018; B = 16'h0084; #100;
A = 16'h0018; B = 16'h0085; #100;
A = 16'h0018; B = 16'h0086; #100;
A = 16'h0018; B = 16'h0087; #100;
A = 16'h0018; B = 16'h0088; #100;
A = 16'h0018; B = 16'h0089; #100;
A = 16'h0018; B = 16'h008A; #100;
A = 16'h0018; B = 16'h008B; #100;
A = 16'h0018; B = 16'h008C; #100;
A = 16'h0018; B = 16'h008D; #100;
A = 16'h0018; B = 16'h008E; #100;
A = 16'h0018; B = 16'h008F; #100;
A = 16'h0018; B = 16'h0090; #100;
A = 16'h0018; B = 16'h0091; #100;
A = 16'h0018; B = 16'h0092; #100;
A = 16'h0018; B = 16'h0093; #100;
A = 16'h0018; B = 16'h0094; #100;
A = 16'h0018; B = 16'h0095; #100;
A = 16'h0018; B = 16'h0096; #100;
A = 16'h0018; B = 16'h0097; #100;
A = 16'h0018; B = 16'h0098; #100;
A = 16'h0018; B = 16'h0099; #100;
A = 16'h0018; B = 16'h009A; #100;
A = 16'h0018; B = 16'h009B; #100;
A = 16'h0018; B = 16'h009C; #100;
A = 16'h0018; B = 16'h009D; #100;
A = 16'h0018; B = 16'h009E; #100;
A = 16'h0018; B = 16'h009F; #100;
A = 16'h0018; B = 16'h00A0; #100;
A = 16'h0018; B = 16'h00A1; #100;
A = 16'h0018; B = 16'h00A2; #100;
A = 16'h0018; B = 16'h00A3; #100;
A = 16'h0018; B = 16'h00A4; #100;
A = 16'h0018; B = 16'h00A5; #100;
A = 16'h0018; B = 16'h00A6; #100;
A = 16'h0018; B = 16'h00A7; #100;
A = 16'h0018; B = 16'h00A8; #100;
A = 16'h0018; B = 16'h00A9; #100;
A = 16'h0018; B = 16'h00AA; #100;
A = 16'h0018; B = 16'h00AB; #100;
A = 16'h0018; B = 16'h00AC; #100;
A = 16'h0018; B = 16'h00AD; #100;
A = 16'h0018; B = 16'h00AE; #100;
A = 16'h0018; B = 16'h00AF; #100;
A = 16'h0018; B = 16'h00B0; #100;
A = 16'h0018; B = 16'h00B1; #100;
A = 16'h0018; B = 16'h00B2; #100;
A = 16'h0018; B = 16'h00B3; #100;
A = 16'h0018; B = 16'h00B4; #100;
A = 16'h0018; B = 16'h00B5; #100;
A = 16'h0018; B = 16'h00B6; #100;
A = 16'h0018; B = 16'h00B7; #100;
A = 16'h0018; B = 16'h00B8; #100;
A = 16'h0018; B = 16'h00B9; #100;
A = 16'h0018; B = 16'h00BA; #100;
A = 16'h0018; B = 16'h00BB; #100;
A = 16'h0018; B = 16'h00BC; #100;
A = 16'h0018; B = 16'h00BD; #100;
A = 16'h0018; B = 16'h00BE; #100;
A = 16'h0018; B = 16'h00BF; #100;
A = 16'h0018; B = 16'h00C0; #100;
A = 16'h0018; B = 16'h00C1; #100;
A = 16'h0018; B = 16'h00C2; #100;
A = 16'h0018; B = 16'h00C3; #100;
A = 16'h0018; B = 16'h00C4; #100;
A = 16'h0018; B = 16'h00C5; #100;
A = 16'h0018; B = 16'h00C6; #100;
A = 16'h0018; B = 16'h00C7; #100;
A = 16'h0018; B = 16'h00C8; #100;
A = 16'h0018; B = 16'h00C9; #100;
A = 16'h0018; B = 16'h00CA; #100;
A = 16'h0018; B = 16'h00CB; #100;
A = 16'h0018; B = 16'h00CC; #100;
A = 16'h0018; B = 16'h00CD; #100;
A = 16'h0018; B = 16'h00CE; #100;
A = 16'h0018; B = 16'h00CF; #100;
A = 16'h0018; B = 16'h00D0; #100;
A = 16'h0018; B = 16'h00D1; #100;
A = 16'h0018; B = 16'h00D2; #100;
A = 16'h0018; B = 16'h00D3; #100;
A = 16'h0018; B = 16'h00D4; #100;
A = 16'h0018; B = 16'h00D5; #100;
A = 16'h0018; B = 16'h00D6; #100;
A = 16'h0018; B = 16'h00D7; #100;
A = 16'h0018; B = 16'h00D8; #100;
A = 16'h0018; B = 16'h00D9; #100;
A = 16'h0018; B = 16'h00DA; #100;
A = 16'h0018; B = 16'h00DB; #100;
A = 16'h0018; B = 16'h00DC; #100;
A = 16'h0018; B = 16'h00DD; #100;
A = 16'h0018; B = 16'h00DE; #100;
A = 16'h0018; B = 16'h00DF; #100;
A = 16'h0018; B = 16'h00E0; #100;
A = 16'h0018; B = 16'h00E1; #100;
A = 16'h0018; B = 16'h00E2; #100;
A = 16'h0018; B = 16'h00E3; #100;
A = 16'h0018; B = 16'h00E4; #100;
A = 16'h0018; B = 16'h00E5; #100;
A = 16'h0018; B = 16'h00E6; #100;
A = 16'h0018; B = 16'h00E7; #100;
A = 16'h0018; B = 16'h00E8; #100;
A = 16'h0018; B = 16'h00E9; #100;
A = 16'h0018; B = 16'h00EA; #100;
A = 16'h0018; B = 16'h00EB; #100;
A = 16'h0018; B = 16'h00EC; #100;
A = 16'h0018; B = 16'h00ED; #100;
A = 16'h0018; B = 16'h00EE; #100;
A = 16'h0018; B = 16'h00EF; #100;
A = 16'h0018; B = 16'h00F0; #100;
A = 16'h0018; B = 16'h00F1; #100;
A = 16'h0018; B = 16'h00F2; #100;
A = 16'h0018; B = 16'h00F3; #100;
A = 16'h0018; B = 16'h00F4; #100;
A = 16'h0018; B = 16'h00F5; #100;
A = 16'h0018; B = 16'h00F6; #100;
A = 16'h0018; B = 16'h00F7; #100;
A = 16'h0018; B = 16'h00F8; #100;
A = 16'h0018; B = 16'h00F9; #100;
A = 16'h0018; B = 16'h00FA; #100;
A = 16'h0018; B = 16'h00FB; #100;
A = 16'h0018; B = 16'h00FC; #100;
A = 16'h0018; B = 16'h00FD; #100;
A = 16'h0018; B = 16'h00FE; #100;
A = 16'h0018; B = 16'h00FF; #100;
A = 16'h0019; B = 16'h000; #100;
A = 16'h0019; B = 16'h001; #100;
A = 16'h0019; B = 16'h002; #100;
A = 16'h0019; B = 16'h003; #100;
A = 16'h0019; B = 16'h004; #100;
A = 16'h0019; B = 16'h005; #100;
A = 16'h0019; B = 16'h006; #100;
A = 16'h0019; B = 16'h007; #100;
A = 16'h0019; B = 16'h008; #100;
A = 16'h0019; B = 16'h009; #100;
A = 16'h0019; B = 16'h00A; #100;
A = 16'h0019; B = 16'h00B; #100;
A = 16'h0019; B = 16'h00C; #100;
A = 16'h0019; B = 16'h00D; #100;
A = 16'h0019; B = 16'h00E; #100;
A = 16'h0019; B = 16'h00F; #100;
A = 16'h0019; B = 16'h0010; #100;
A = 16'h0019; B = 16'h0011; #100;
A = 16'h0019; B = 16'h0012; #100;
A = 16'h0019; B = 16'h0013; #100;
A = 16'h0019; B = 16'h0014; #100;
A = 16'h0019; B = 16'h0015; #100;
A = 16'h0019; B = 16'h0016; #100;
A = 16'h0019; B = 16'h0017; #100;
A = 16'h0019; B = 16'h0018; #100;
A = 16'h0019; B = 16'h0019; #100;
A = 16'h0019; B = 16'h001A; #100;
A = 16'h0019; B = 16'h001B; #100;
A = 16'h0019; B = 16'h001C; #100;
A = 16'h0019; B = 16'h001D; #100;
A = 16'h0019; B = 16'h001E; #100;
A = 16'h0019; B = 16'h001F; #100;
A = 16'h0019; B = 16'h0020; #100;
A = 16'h0019; B = 16'h0021; #100;
A = 16'h0019; B = 16'h0022; #100;
A = 16'h0019; B = 16'h0023; #100;
A = 16'h0019; B = 16'h0024; #100;
A = 16'h0019; B = 16'h0025; #100;
A = 16'h0019; B = 16'h0026; #100;
A = 16'h0019; B = 16'h0027; #100;
A = 16'h0019; B = 16'h0028; #100;
A = 16'h0019; B = 16'h0029; #100;
A = 16'h0019; B = 16'h002A; #100;
A = 16'h0019; B = 16'h002B; #100;
A = 16'h0019; B = 16'h002C; #100;
A = 16'h0019; B = 16'h002D; #100;
A = 16'h0019; B = 16'h002E; #100;
A = 16'h0019; B = 16'h002F; #100;
A = 16'h0019; B = 16'h0030; #100;
A = 16'h0019; B = 16'h0031; #100;
A = 16'h0019; B = 16'h0032; #100;
A = 16'h0019; B = 16'h0033; #100;
A = 16'h0019; B = 16'h0034; #100;
A = 16'h0019; B = 16'h0035; #100;
A = 16'h0019; B = 16'h0036; #100;
A = 16'h0019; B = 16'h0037; #100;
A = 16'h0019; B = 16'h0038; #100;
A = 16'h0019; B = 16'h0039; #100;
A = 16'h0019; B = 16'h003A; #100;
A = 16'h0019; B = 16'h003B; #100;
A = 16'h0019; B = 16'h003C; #100;
A = 16'h0019; B = 16'h003D; #100;
A = 16'h0019; B = 16'h003E; #100;
A = 16'h0019; B = 16'h003F; #100;
A = 16'h0019; B = 16'h0040; #100;
A = 16'h0019; B = 16'h0041; #100;
A = 16'h0019; B = 16'h0042; #100;
A = 16'h0019; B = 16'h0043; #100;
A = 16'h0019; B = 16'h0044; #100;
A = 16'h0019; B = 16'h0045; #100;
A = 16'h0019; B = 16'h0046; #100;
A = 16'h0019; B = 16'h0047; #100;
A = 16'h0019; B = 16'h0048; #100;
A = 16'h0019; B = 16'h0049; #100;
A = 16'h0019; B = 16'h004A; #100;
A = 16'h0019; B = 16'h004B; #100;
A = 16'h0019; B = 16'h004C; #100;
A = 16'h0019; B = 16'h004D; #100;
A = 16'h0019; B = 16'h004E; #100;
A = 16'h0019; B = 16'h004F; #100;
A = 16'h0019; B = 16'h0050; #100;
A = 16'h0019; B = 16'h0051; #100;
A = 16'h0019; B = 16'h0052; #100;
A = 16'h0019; B = 16'h0053; #100;
A = 16'h0019; B = 16'h0054; #100;
A = 16'h0019; B = 16'h0055; #100;
A = 16'h0019; B = 16'h0056; #100;
A = 16'h0019; B = 16'h0057; #100;
A = 16'h0019; B = 16'h0058; #100;
A = 16'h0019; B = 16'h0059; #100;
A = 16'h0019; B = 16'h005A; #100;
A = 16'h0019; B = 16'h005B; #100;
A = 16'h0019; B = 16'h005C; #100;
A = 16'h0019; B = 16'h005D; #100;
A = 16'h0019; B = 16'h005E; #100;
A = 16'h0019; B = 16'h005F; #100;
A = 16'h0019; B = 16'h0060; #100;
A = 16'h0019; B = 16'h0061; #100;
A = 16'h0019; B = 16'h0062; #100;
A = 16'h0019; B = 16'h0063; #100;
A = 16'h0019; B = 16'h0064; #100;
A = 16'h0019; B = 16'h0065; #100;
A = 16'h0019; B = 16'h0066; #100;
A = 16'h0019; B = 16'h0067; #100;
A = 16'h0019; B = 16'h0068; #100;
A = 16'h0019; B = 16'h0069; #100;
A = 16'h0019; B = 16'h006A; #100;
A = 16'h0019; B = 16'h006B; #100;
A = 16'h0019; B = 16'h006C; #100;
A = 16'h0019; B = 16'h006D; #100;
A = 16'h0019; B = 16'h006E; #100;
A = 16'h0019; B = 16'h006F; #100;
A = 16'h0019; B = 16'h0070; #100;
A = 16'h0019; B = 16'h0071; #100;
A = 16'h0019; B = 16'h0072; #100;
A = 16'h0019; B = 16'h0073; #100;
A = 16'h0019; B = 16'h0074; #100;
A = 16'h0019; B = 16'h0075; #100;
A = 16'h0019; B = 16'h0076; #100;
A = 16'h0019; B = 16'h0077; #100;
A = 16'h0019; B = 16'h0078; #100;
A = 16'h0019; B = 16'h0079; #100;
A = 16'h0019; B = 16'h007A; #100;
A = 16'h0019; B = 16'h007B; #100;
A = 16'h0019; B = 16'h007C; #100;
A = 16'h0019; B = 16'h007D; #100;
A = 16'h0019; B = 16'h007E; #100;
A = 16'h0019; B = 16'h007F; #100;
A = 16'h0019; B = 16'h0080; #100;
A = 16'h0019; B = 16'h0081; #100;
A = 16'h0019; B = 16'h0082; #100;
A = 16'h0019; B = 16'h0083; #100;
A = 16'h0019; B = 16'h0084; #100;
A = 16'h0019; B = 16'h0085; #100;
A = 16'h0019; B = 16'h0086; #100;
A = 16'h0019; B = 16'h0087; #100;
A = 16'h0019; B = 16'h0088; #100;
A = 16'h0019; B = 16'h0089; #100;
A = 16'h0019; B = 16'h008A; #100;
A = 16'h0019; B = 16'h008B; #100;
A = 16'h0019; B = 16'h008C; #100;
A = 16'h0019; B = 16'h008D; #100;
A = 16'h0019; B = 16'h008E; #100;
A = 16'h0019; B = 16'h008F; #100;
A = 16'h0019; B = 16'h0090; #100;
A = 16'h0019; B = 16'h0091; #100;
A = 16'h0019; B = 16'h0092; #100;
A = 16'h0019; B = 16'h0093; #100;
A = 16'h0019; B = 16'h0094; #100;
A = 16'h0019; B = 16'h0095; #100;
A = 16'h0019; B = 16'h0096; #100;
A = 16'h0019; B = 16'h0097; #100;
A = 16'h0019; B = 16'h0098; #100;
A = 16'h0019; B = 16'h0099; #100;
A = 16'h0019; B = 16'h009A; #100;
A = 16'h0019; B = 16'h009B; #100;
A = 16'h0019; B = 16'h009C; #100;
A = 16'h0019; B = 16'h009D; #100;
A = 16'h0019; B = 16'h009E; #100;
A = 16'h0019; B = 16'h009F; #100;
A = 16'h0019; B = 16'h00A0; #100;
A = 16'h0019; B = 16'h00A1; #100;
A = 16'h0019; B = 16'h00A2; #100;
A = 16'h0019; B = 16'h00A3; #100;
A = 16'h0019; B = 16'h00A4; #100;
A = 16'h0019; B = 16'h00A5; #100;
A = 16'h0019; B = 16'h00A6; #100;
A = 16'h0019; B = 16'h00A7; #100;
A = 16'h0019; B = 16'h00A8; #100;
A = 16'h0019; B = 16'h00A9; #100;
A = 16'h0019; B = 16'h00AA; #100;
A = 16'h0019; B = 16'h00AB; #100;
A = 16'h0019; B = 16'h00AC; #100;
A = 16'h0019; B = 16'h00AD; #100;
A = 16'h0019; B = 16'h00AE; #100;
A = 16'h0019; B = 16'h00AF; #100;
A = 16'h0019; B = 16'h00B0; #100;
A = 16'h0019; B = 16'h00B1; #100;
A = 16'h0019; B = 16'h00B2; #100;
A = 16'h0019; B = 16'h00B3; #100;
A = 16'h0019; B = 16'h00B4; #100;
A = 16'h0019; B = 16'h00B5; #100;
A = 16'h0019; B = 16'h00B6; #100;
A = 16'h0019; B = 16'h00B7; #100;
A = 16'h0019; B = 16'h00B8; #100;
A = 16'h0019; B = 16'h00B9; #100;
A = 16'h0019; B = 16'h00BA; #100;
A = 16'h0019; B = 16'h00BB; #100;
A = 16'h0019; B = 16'h00BC; #100;
A = 16'h0019; B = 16'h00BD; #100;
A = 16'h0019; B = 16'h00BE; #100;
A = 16'h0019; B = 16'h00BF; #100;
A = 16'h0019; B = 16'h00C0; #100;
A = 16'h0019; B = 16'h00C1; #100;
A = 16'h0019; B = 16'h00C2; #100;
A = 16'h0019; B = 16'h00C3; #100;
A = 16'h0019; B = 16'h00C4; #100;
A = 16'h0019; B = 16'h00C5; #100;
A = 16'h0019; B = 16'h00C6; #100;
A = 16'h0019; B = 16'h00C7; #100;
A = 16'h0019; B = 16'h00C8; #100;
A = 16'h0019; B = 16'h00C9; #100;
A = 16'h0019; B = 16'h00CA; #100;
A = 16'h0019; B = 16'h00CB; #100;
A = 16'h0019; B = 16'h00CC; #100;
A = 16'h0019; B = 16'h00CD; #100;
A = 16'h0019; B = 16'h00CE; #100;
A = 16'h0019; B = 16'h00CF; #100;
A = 16'h0019; B = 16'h00D0; #100;
A = 16'h0019; B = 16'h00D1; #100;
A = 16'h0019; B = 16'h00D2; #100;
A = 16'h0019; B = 16'h00D3; #100;
A = 16'h0019; B = 16'h00D4; #100;
A = 16'h0019; B = 16'h00D5; #100;
A = 16'h0019; B = 16'h00D6; #100;
A = 16'h0019; B = 16'h00D7; #100;
A = 16'h0019; B = 16'h00D8; #100;
A = 16'h0019; B = 16'h00D9; #100;
A = 16'h0019; B = 16'h00DA; #100;
A = 16'h0019; B = 16'h00DB; #100;
A = 16'h0019; B = 16'h00DC; #100;
A = 16'h0019; B = 16'h00DD; #100;
A = 16'h0019; B = 16'h00DE; #100;
A = 16'h0019; B = 16'h00DF; #100;
A = 16'h0019; B = 16'h00E0; #100;
A = 16'h0019; B = 16'h00E1; #100;
A = 16'h0019; B = 16'h00E2; #100;
A = 16'h0019; B = 16'h00E3; #100;
A = 16'h0019; B = 16'h00E4; #100;
A = 16'h0019; B = 16'h00E5; #100;
A = 16'h0019; B = 16'h00E6; #100;
A = 16'h0019; B = 16'h00E7; #100;
A = 16'h0019; B = 16'h00E8; #100;
A = 16'h0019; B = 16'h00E9; #100;
A = 16'h0019; B = 16'h00EA; #100;
A = 16'h0019; B = 16'h00EB; #100;
A = 16'h0019; B = 16'h00EC; #100;
A = 16'h0019; B = 16'h00ED; #100;
A = 16'h0019; B = 16'h00EE; #100;
A = 16'h0019; B = 16'h00EF; #100;
A = 16'h0019; B = 16'h00F0; #100;
A = 16'h0019; B = 16'h00F1; #100;
A = 16'h0019; B = 16'h00F2; #100;
A = 16'h0019; B = 16'h00F3; #100;
A = 16'h0019; B = 16'h00F4; #100;
A = 16'h0019; B = 16'h00F5; #100;
A = 16'h0019; B = 16'h00F6; #100;
A = 16'h0019; B = 16'h00F7; #100;
A = 16'h0019; B = 16'h00F8; #100;
A = 16'h0019; B = 16'h00F9; #100;
A = 16'h0019; B = 16'h00FA; #100;
A = 16'h0019; B = 16'h00FB; #100;
A = 16'h0019; B = 16'h00FC; #100;
A = 16'h0019; B = 16'h00FD; #100;
A = 16'h0019; B = 16'h00FE; #100;
A = 16'h0019; B = 16'h00FF; #100;
A = 16'h001A; B = 16'h000; #100;
A = 16'h001A; B = 16'h001; #100;
A = 16'h001A; B = 16'h002; #100;
A = 16'h001A; B = 16'h003; #100;
A = 16'h001A; B = 16'h004; #100;
A = 16'h001A; B = 16'h005; #100;
A = 16'h001A; B = 16'h006; #100;
A = 16'h001A; B = 16'h007; #100;
A = 16'h001A; B = 16'h008; #100;
A = 16'h001A; B = 16'h009; #100;
A = 16'h001A; B = 16'h00A; #100;
A = 16'h001A; B = 16'h00B; #100;
A = 16'h001A; B = 16'h00C; #100;
A = 16'h001A; B = 16'h00D; #100;
A = 16'h001A; B = 16'h00E; #100;
A = 16'h001A; B = 16'h00F; #100;
A = 16'h001A; B = 16'h0010; #100;
A = 16'h001A; B = 16'h0011; #100;
A = 16'h001A; B = 16'h0012; #100;
A = 16'h001A; B = 16'h0013; #100;
A = 16'h001A; B = 16'h0014; #100;
A = 16'h001A; B = 16'h0015; #100;
A = 16'h001A; B = 16'h0016; #100;
A = 16'h001A; B = 16'h0017; #100;
A = 16'h001A; B = 16'h0018; #100;
A = 16'h001A; B = 16'h0019; #100;
A = 16'h001A; B = 16'h001A; #100;
A = 16'h001A; B = 16'h001B; #100;
A = 16'h001A; B = 16'h001C; #100;
A = 16'h001A; B = 16'h001D; #100;
A = 16'h001A; B = 16'h001E; #100;
A = 16'h001A; B = 16'h001F; #100;
A = 16'h001A; B = 16'h0020; #100;
A = 16'h001A; B = 16'h0021; #100;
A = 16'h001A; B = 16'h0022; #100;
A = 16'h001A; B = 16'h0023; #100;
A = 16'h001A; B = 16'h0024; #100;
A = 16'h001A; B = 16'h0025; #100;
A = 16'h001A; B = 16'h0026; #100;
A = 16'h001A; B = 16'h0027; #100;
A = 16'h001A; B = 16'h0028; #100;
A = 16'h001A; B = 16'h0029; #100;
A = 16'h001A; B = 16'h002A; #100;
A = 16'h001A; B = 16'h002B; #100;
A = 16'h001A; B = 16'h002C; #100;
A = 16'h001A; B = 16'h002D; #100;
A = 16'h001A; B = 16'h002E; #100;
A = 16'h001A; B = 16'h002F; #100;
A = 16'h001A; B = 16'h0030; #100;
A = 16'h001A; B = 16'h0031; #100;
A = 16'h001A; B = 16'h0032; #100;
A = 16'h001A; B = 16'h0033; #100;
A = 16'h001A; B = 16'h0034; #100;
A = 16'h001A; B = 16'h0035; #100;
A = 16'h001A; B = 16'h0036; #100;
A = 16'h001A; B = 16'h0037; #100;
A = 16'h001A; B = 16'h0038; #100;
A = 16'h001A; B = 16'h0039; #100;
A = 16'h001A; B = 16'h003A; #100;
A = 16'h001A; B = 16'h003B; #100;
A = 16'h001A; B = 16'h003C; #100;
A = 16'h001A; B = 16'h003D; #100;
A = 16'h001A; B = 16'h003E; #100;
A = 16'h001A; B = 16'h003F; #100;
A = 16'h001A; B = 16'h0040; #100;
A = 16'h001A; B = 16'h0041; #100;
A = 16'h001A; B = 16'h0042; #100;
A = 16'h001A; B = 16'h0043; #100;
A = 16'h001A; B = 16'h0044; #100;
A = 16'h001A; B = 16'h0045; #100;
A = 16'h001A; B = 16'h0046; #100;
A = 16'h001A; B = 16'h0047; #100;
A = 16'h001A; B = 16'h0048; #100;
A = 16'h001A; B = 16'h0049; #100;
A = 16'h001A; B = 16'h004A; #100;
A = 16'h001A; B = 16'h004B; #100;
A = 16'h001A; B = 16'h004C; #100;
A = 16'h001A; B = 16'h004D; #100;
A = 16'h001A; B = 16'h004E; #100;
A = 16'h001A; B = 16'h004F; #100;
A = 16'h001A; B = 16'h0050; #100;
A = 16'h001A; B = 16'h0051; #100;
A = 16'h001A; B = 16'h0052; #100;
A = 16'h001A; B = 16'h0053; #100;
A = 16'h001A; B = 16'h0054; #100;
A = 16'h001A; B = 16'h0055; #100;
A = 16'h001A; B = 16'h0056; #100;
A = 16'h001A; B = 16'h0057; #100;
A = 16'h001A; B = 16'h0058; #100;
A = 16'h001A; B = 16'h0059; #100;
A = 16'h001A; B = 16'h005A; #100;
A = 16'h001A; B = 16'h005B; #100;
A = 16'h001A; B = 16'h005C; #100;
A = 16'h001A; B = 16'h005D; #100;
A = 16'h001A; B = 16'h005E; #100;
A = 16'h001A; B = 16'h005F; #100;
A = 16'h001A; B = 16'h0060; #100;
A = 16'h001A; B = 16'h0061; #100;
A = 16'h001A; B = 16'h0062; #100;
A = 16'h001A; B = 16'h0063; #100;
A = 16'h001A; B = 16'h0064; #100;
A = 16'h001A; B = 16'h0065; #100;
A = 16'h001A; B = 16'h0066; #100;
A = 16'h001A; B = 16'h0067; #100;
A = 16'h001A; B = 16'h0068; #100;
A = 16'h001A; B = 16'h0069; #100;
A = 16'h001A; B = 16'h006A; #100;
A = 16'h001A; B = 16'h006B; #100;
A = 16'h001A; B = 16'h006C; #100;
A = 16'h001A; B = 16'h006D; #100;
A = 16'h001A; B = 16'h006E; #100;
A = 16'h001A; B = 16'h006F; #100;
A = 16'h001A; B = 16'h0070; #100;
A = 16'h001A; B = 16'h0071; #100;
A = 16'h001A; B = 16'h0072; #100;
A = 16'h001A; B = 16'h0073; #100;
A = 16'h001A; B = 16'h0074; #100;
A = 16'h001A; B = 16'h0075; #100;
A = 16'h001A; B = 16'h0076; #100;
A = 16'h001A; B = 16'h0077; #100;
A = 16'h001A; B = 16'h0078; #100;
A = 16'h001A; B = 16'h0079; #100;
A = 16'h001A; B = 16'h007A; #100;
A = 16'h001A; B = 16'h007B; #100;
A = 16'h001A; B = 16'h007C; #100;
A = 16'h001A; B = 16'h007D; #100;
A = 16'h001A; B = 16'h007E; #100;
A = 16'h001A; B = 16'h007F; #100;
A = 16'h001A; B = 16'h0080; #100;
A = 16'h001A; B = 16'h0081; #100;
A = 16'h001A; B = 16'h0082; #100;
A = 16'h001A; B = 16'h0083; #100;
A = 16'h001A; B = 16'h0084; #100;
A = 16'h001A; B = 16'h0085; #100;
A = 16'h001A; B = 16'h0086; #100;
A = 16'h001A; B = 16'h0087; #100;
A = 16'h001A; B = 16'h0088; #100;
A = 16'h001A; B = 16'h0089; #100;
A = 16'h001A; B = 16'h008A; #100;
A = 16'h001A; B = 16'h008B; #100;
A = 16'h001A; B = 16'h008C; #100;
A = 16'h001A; B = 16'h008D; #100;
A = 16'h001A; B = 16'h008E; #100;
A = 16'h001A; B = 16'h008F; #100;
A = 16'h001A; B = 16'h0090; #100;
A = 16'h001A; B = 16'h0091; #100;
A = 16'h001A; B = 16'h0092; #100;
A = 16'h001A; B = 16'h0093; #100;
A = 16'h001A; B = 16'h0094; #100;
A = 16'h001A; B = 16'h0095; #100;
A = 16'h001A; B = 16'h0096; #100;
A = 16'h001A; B = 16'h0097; #100;
A = 16'h001A; B = 16'h0098; #100;
A = 16'h001A; B = 16'h0099; #100;
A = 16'h001A; B = 16'h009A; #100;
A = 16'h001A; B = 16'h009B; #100;
A = 16'h001A; B = 16'h009C; #100;
A = 16'h001A; B = 16'h009D; #100;
A = 16'h001A; B = 16'h009E; #100;
A = 16'h001A; B = 16'h009F; #100;
A = 16'h001A; B = 16'h00A0; #100;
A = 16'h001A; B = 16'h00A1; #100;
A = 16'h001A; B = 16'h00A2; #100;
A = 16'h001A; B = 16'h00A3; #100;
A = 16'h001A; B = 16'h00A4; #100;
A = 16'h001A; B = 16'h00A5; #100;
A = 16'h001A; B = 16'h00A6; #100;
A = 16'h001A; B = 16'h00A7; #100;
A = 16'h001A; B = 16'h00A8; #100;
A = 16'h001A; B = 16'h00A9; #100;
A = 16'h001A; B = 16'h00AA; #100;
A = 16'h001A; B = 16'h00AB; #100;
A = 16'h001A; B = 16'h00AC; #100;
A = 16'h001A; B = 16'h00AD; #100;
A = 16'h001A; B = 16'h00AE; #100;
A = 16'h001A; B = 16'h00AF; #100;
A = 16'h001A; B = 16'h00B0; #100;
A = 16'h001A; B = 16'h00B1; #100;
A = 16'h001A; B = 16'h00B2; #100;
A = 16'h001A; B = 16'h00B3; #100;
A = 16'h001A; B = 16'h00B4; #100;
A = 16'h001A; B = 16'h00B5; #100;
A = 16'h001A; B = 16'h00B6; #100;
A = 16'h001A; B = 16'h00B7; #100;
A = 16'h001A; B = 16'h00B8; #100;
A = 16'h001A; B = 16'h00B9; #100;
A = 16'h001A; B = 16'h00BA; #100;
A = 16'h001A; B = 16'h00BB; #100;
A = 16'h001A; B = 16'h00BC; #100;
A = 16'h001A; B = 16'h00BD; #100;
A = 16'h001A; B = 16'h00BE; #100;
A = 16'h001A; B = 16'h00BF; #100;
A = 16'h001A; B = 16'h00C0; #100;
A = 16'h001A; B = 16'h00C1; #100;
A = 16'h001A; B = 16'h00C2; #100;
A = 16'h001A; B = 16'h00C3; #100;
A = 16'h001A; B = 16'h00C4; #100;
A = 16'h001A; B = 16'h00C5; #100;
A = 16'h001A; B = 16'h00C6; #100;
A = 16'h001A; B = 16'h00C7; #100;
A = 16'h001A; B = 16'h00C8; #100;
A = 16'h001A; B = 16'h00C9; #100;
A = 16'h001A; B = 16'h00CA; #100;
A = 16'h001A; B = 16'h00CB; #100;
A = 16'h001A; B = 16'h00CC; #100;
A = 16'h001A; B = 16'h00CD; #100;
A = 16'h001A; B = 16'h00CE; #100;
A = 16'h001A; B = 16'h00CF; #100;
A = 16'h001A; B = 16'h00D0; #100;
A = 16'h001A; B = 16'h00D1; #100;
A = 16'h001A; B = 16'h00D2; #100;
A = 16'h001A; B = 16'h00D3; #100;
A = 16'h001A; B = 16'h00D4; #100;
A = 16'h001A; B = 16'h00D5; #100;
A = 16'h001A; B = 16'h00D6; #100;
A = 16'h001A; B = 16'h00D7; #100;
A = 16'h001A; B = 16'h00D8; #100;
A = 16'h001A; B = 16'h00D9; #100;
A = 16'h001A; B = 16'h00DA; #100;
A = 16'h001A; B = 16'h00DB; #100;
A = 16'h001A; B = 16'h00DC; #100;
A = 16'h001A; B = 16'h00DD; #100;
A = 16'h001A; B = 16'h00DE; #100;
A = 16'h001A; B = 16'h00DF; #100;
A = 16'h001A; B = 16'h00E0; #100;
A = 16'h001A; B = 16'h00E1; #100;
A = 16'h001A; B = 16'h00E2; #100;
A = 16'h001A; B = 16'h00E3; #100;
A = 16'h001A; B = 16'h00E4; #100;
A = 16'h001A; B = 16'h00E5; #100;
A = 16'h001A; B = 16'h00E6; #100;
A = 16'h001A; B = 16'h00E7; #100;
A = 16'h001A; B = 16'h00E8; #100;
A = 16'h001A; B = 16'h00E9; #100;
A = 16'h001A; B = 16'h00EA; #100;
A = 16'h001A; B = 16'h00EB; #100;
A = 16'h001A; B = 16'h00EC; #100;
A = 16'h001A; B = 16'h00ED; #100;
A = 16'h001A; B = 16'h00EE; #100;
A = 16'h001A; B = 16'h00EF; #100;
A = 16'h001A; B = 16'h00F0; #100;
A = 16'h001A; B = 16'h00F1; #100;
A = 16'h001A; B = 16'h00F2; #100;
A = 16'h001A; B = 16'h00F3; #100;
A = 16'h001A; B = 16'h00F4; #100;
A = 16'h001A; B = 16'h00F5; #100;
A = 16'h001A; B = 16'h00F6; #100;
A = 16'h001A; B = 16'h00F7; #100;
A = 16'h001A; B = 16'h00F8; #100;
A = 16'h001A; B = 16'h00F9; #100;
A = 16'h001A; B = 16'h00FA; #100;
A = 16'h001A; B = 16'h00FB; #100;
A = 16'h001A; B = 16'h00FC; #100;
A = 16'h001A; B = 16'h00FD; #100;
A = 16'h001A; B = 16'h00FE; #100;
A = 16'h001A; B = 16'h00FF; #100;
A = 16'h001B; B = 16'h000; #100;
A = 16'h001B; B = 16'h001; #100;
A = 16'h001B; B = 16'h002; #100;
A = 16'h001B; B = 16'h003; #100;
A = 16'h001B; B = 16'h004; #100;
A = 16'h001B; B = 16'h005; #100;
A = 16'h001B; B = 16'h006; #100;
A = 16'h001B; B = 16'h007; #100;
A = 16'h001B; B = 16'h008; #100;
A = 16'h001B; B = 16'h009; #100;
A = 16'h001B; B = 16'h00A; #100;
A = 16'h001B; B = 16'h00B; #100;
A = 16'h001B; B = 16'h00C; #100;
A = 16'h001B; B = 16'h00D; #100;
A = 16'h001B; B = 16'h00E; #100;
A = 16'h001B; B = 16'h00F; #100;
A = 16'h001B; B = 16'h0010; #100;
A = 16'h001B; B = 16'h0011; #100;
A = 16'h001B; B = 16'h0012; #100;
A = 16'h001B; B = 16'h0013; #100;
A = 16'h001B; B = 16'h0014; #100;
A = 16'h001B; B = 16'h0015; #100;
A = 16'h001B; B = 16'h0016; #100;
A = 16'h001B; B = 16'h0017; #100;
A = 16'h001B; B = 16'h0018; #100;
A = 16'h001B; B = 16'h0019; #100;
A = 16'h001B; B = 16'h001A; #100;
A = 16'h001B; B = 16'h001B; #100;
A = 16'h001B; B = 16'h001C; #100;
A = 16'h001B; B = 16'h001D; #100;
A = 16'h001B; B = 16'h001E; #100;
A = 16'h001B; B = 16'h001F; #100;
A = 16'h001B; B = 16'h0020; #100;
A = 16'h001B; B = 16'h0021; #100;
A = 16'h001B; B = 16'h0022; #100;
A = 16'h001B; B = 16'h0023; #100;
A = 16'h001B; B = 16'h0024; #100;
A = 16'h001B; B = 16'h0025; #100;
A = 16'h001B; B = 16'h0026; #100;
A = 16'h001B; B = 16'h0027; #100;
A = 16'h001B; B = 16'h0028; #100;
A = 16'h001B; B = 16'h0029; #100;
A = 16'h001B; B = 16'h002A; #100;
A = 16'h001B; B = 16'h002B; #100;
A = 16'h001B; B = 16'h002C; #100;
A = 16'h001B; B = 16'h002D; #100;
A = 16'h001B; B = 16'h002E; #100;
A = 16'h001B; B = 16'h002F; #100;
A = 16'h001B; B = 16'h0030; #100;
A = 16'h001B; B = 16'h0031; #100;
A = 16'h001B; B = 16'h0032; #100;
A = 16'h001B; B = 16'h0033; #100;
A = 16'h001B; B = 16'h0034; #100;
A = 16'h001B; B = 16'h0035; #100;
A = 16'h001B; B = 16'h0036; #100;
A = 16'h001B; B = 16'h0037; #100;
A = 16'h001B; B = 16'h0038; #100;
A = 16'h001B; B = 16'h0039; #100;
A = 16'h001B; B = 16'h003A; #100;
A = 16'h001B; B = 16'h003B; #100;
A = 16'h001B; B = 16'h003C; #100;
A = 16'h001B; B = 16'h003D; #100;
A = 16'h001B; B = 16'h003E; #100;
A = 16'h001B; B = 16'h003F; #100;
A = 16'h001B; B = 16'h0040; #100;
A = 16'h001B; B = 16'h0041; #100;
A = 16'h001B; B = 16'h0042; #100;
A = 16'h001B; B = 16'h0043; #100;
A = 16'h001B; B = 16'h0044; #100;
A = 16'h001B; B = 16'h0045; #100;
A = 16'h001B; B = 16'h0046; #100;
A = 16'h001B; B = 16'h0047; #100;
A = 16'h001B; B = 16'h0048; #100;
A = 16'h001B; B = 16'h0049; #100;
A = 16'h001B; B = 16'h004A; #100;
A = 16'h001B; B = 16'h004B; #100;
A = 16'h001B; B = 16'h004C; #100;
A = 16'h001B; B = 16'h004D; #100;
A = 16'h001B; B = 16'h004E; #100;
A = 16'h001B; B = 16'h004F; #100;
A = 16'h001B; B = 16'h0050; #100;
A = 16'h001B; B = 16'h0051; #100;
A = 16'h001B; B = 16'h0052; #100;
A = 16'h001B; B = 16'h0053; #100;
A = 16'h001B; B = 16'h0054; #100;
A = 16'h001B; B = 16'h0055; #100;
A = 16'h001B; B = 16'h0056; #100;
A = 16'h001B; B = 16'h0057; #100;
A = 16'h001B; B = 16'h0058; #100;
A = 16'h001B; B = 16'h0059; #100;
A = 16'h001B; B = 16'h005A; #100;
A = 16'h001B; B = 16'h005B; #100;
A = 16'h001B; B = 16'h005C; #100;
A = 16'h001B; B = 16'h005D; #100;
A = 16'h001B; B = 16'h005E; #100;
A = 16'h001B; B = 16'h005F; #100;
A = 16'h001B; B = 16'h0060; #100;
A = 16'h001B; B = 16'h0061; #100;
A = 16'h001B; B = 16'h0062; #100;
A = 16'h001B; B = 16'h0063; #100;
A = 16'h001B; B = 16'h0064; #100;
A = 16'h001B; B = 16'h0065; #100;
A = 16'h001B; B = 16'h0066; #100;
A = 16'h001B; B = 16'h0067; #100;
A = 16'h001B; B = 16'h0068; #100;
A = 16'h001B; B = 16'h0069; #100;
A = 16'h001B; B = 16'h006A; #100;
A = 16'h001B; B = 16'h006B; #100;
A = 16'h001B; B = 16'h006C; #100;
A = 16'h001B; B = 16'h006D; #100;
A = 16'h001B; B = 16'h006E; #100;
A = 16'h001B; B = 16'h006F; #100;
A = 16'h001B; B = 16'h0070; #100;
A = 16'h001B; B = 16'h0071; #100;
A = 16'h001B; B = 16'h0072; #100;
A = 16'h001B; B = 16'h0073; #100;
A = 16'h001B; B = 16'h0074; #100;
A = 16'h001B; B = 16'h0075; #100;
A = 16'h001B; B = 16'h0076; #100;
A = 16'h001B; B = 16'h0077; #100;
A = 16'h001B; B = 16'h0078; #100;
A = 16'h001B; B = 16'h0079; #100;
A = 16'h001B; B = 16'h007A; #100;
A = 16'h001B; B = 16'h007B; #100;
A = 16'h001B; B = 16'h007C; #100;
A = 16'h001B; B = 16'h007D; #100;
A = 16'h001B; B = 16'h007E; #100;
A = 16'h001B; B = 16'h007F; #100;
A = 16'h001B; B = 16'h0080; #100;
A = 16'h001B; B = 16'h0081; #100;
A = 16'h001B; B = 16'h0082; #100;
A = 16'h001B; B = 16'h0083; #100;
A = 16'h001B; B = 16'h0084; #100;
A = 16'h001B; B = 16'h0085; #100;
A = 16'h001B; B = 16'h0086; #100;
A = 16'h001B; B = 16'h0087; #100;
A = 16'h001B; B = 16'h0088; #100;
A = 16'h001B; B = 16'h0089; #100;
A = 16'h001B; B = 16'h008A; #100;
A = 16'h001B; B = 16'h008B; #100;
A = 16'h001B; B = 16'h008C; #100;
A = 16'h001B; B = 16'h008D; #100;
A = 16'h001B; B = 16'h008E; #100;
A = 16'h001B; B = 16'h008F; #100;
A = 16'h001B; B = 16'h0090; #100;
A = 16'h001B; B = 16'h0091; #100;
A = 16'h001B; B = 16'h0092; #100;
A = 16'h001B; B = 16'h0093; #100;
A = 16'h001B; B = 16'h0094; #100;
A = 16'h001B; B = 16'h0095; #100;
A = 16'h001B; B = 16'h0096; #100;
A = 16'h001B; B = 16'h0097; #100;
A = 16'h001B; B = 16'h0098; #100;
A = 16'h001B; B = 16'h0099; #100;
A = 16'h001B; B = 16'h009A; #100;
A = 16'h001B; B = 16'h009B; #100;
A = 16'h001B; B = 16'h009C; #100;
A = 16'h001B; B = 16'h009D; #100;
A = 16'h001B; B = 16'h009E; #100;
A = 16'h001B; B = 16'h009F; #100;
A = 16'h001B; B = 16'h00A0; #100;
A = 16'h001B; B = 16'h00A1; #100;
A = 16'h001B; B = 16'h00A2; #100;
A = 16'h001B; B = 16'h00A3; #100;
A = 16'h001B; B = 16'h00A4; #100;
A = 16'h001B; B = 16'h00A5; #100;
A = 16'h001B; B = 16'h00A6; #100;
A = 16'h001B; B = 16'h00A7; #100;
A = 16'h001B; B = 16'h00A8; #100;
A = 16'h001B; B = 16'h00A9; #100;
A = 16'h001B; B = 16'h00AA; #100;
A = 16'h001B; B = 16'h00AB; #100;
A = 16'h001B; B = 16'h00AC; #100;
A = 16'h001B; B = 16'h00AD; #100;
A = 16'h001B; B = 16'h00AE; #100;
A = 16'h001B; B = 16'h00AF; #100;
A = 16'h001B; B = 16'h00B0; #100;
A = 16'h001B; B = 16'h00B1; #100;
A = 16'h001B; B = 16'h00B2; #100;
A = 16'h001B; B = 16'h00B3; #100;
A = 16'h001B; B = 16'h00B4; #100;
A = 16'h001B; B = 16'h00B5; #100;
A = 16'h001B; B = 16'h00B6; #100;
A = 16'h001B; B = 16'h00B7; #100;
A = 16'h001B; B = 16'h00B8; #100;
A = 16'h001B; B = 16'h00B9; #100;
A = 16'h001B; B = 16'h00BA; #100;
A = 16'h001B; B = 16'h00BB; #100;
A = 16'h001B; B = 16'h00BC; #100;
A = 16'h001B; B = 16'h00BD; #100;
A = 16'h001B; B = 16'h00BE; #100;
A = 16'h001B; B = 16'h00BF; #100;
A = 16'h001B; B = 16'h00C0; #100;
A = 16'h001B; B = 16'h00C1; #100;
A = 16'h001B; B = 16'h00C2; #100;
A = 16'h001B; B = 16'h00C3; #100;
A = 16'h001B; B = 16'h00C4; #100;
A = 16'h001B; B = 16'h00C5; #100;
A = 16'h001B; B = 16'h00C6; #100;
A = 16'h001B; B = 16'h00C7; #100;
A = 16'h001B; B = 16'h00C8; #100;
A = 16'h001B; B = 16'h00C9; #100;
A = 16'h001B; B = 16'h00CA; #100;
A = 16'h001B; B = 16'h00CB; #100;
A = 16'h001B; B = 16'h00CC; #100;
A = 16'h001B; B = 16'h00CD; #100;
A = 16'h001B; B = 16'h00CE; #100;
A = 16'h001B; B = 16'h00CF; #100;
A = 16'h001B; B = 16'h00D0; #100;
A = 16'h001B; B = 16'h00D1; #100;
A = 16'h001B; B = 16'h00D2; #100;
A = 16'h001B; B = 16'h00D3; #100;
A = 16'h001B; B = 16'h00D4; #100;
A = 16'h001B; B = 16'h00D5; #100;
A = 16'h001B; B = 16'h00D6; #100;
A = 16'h001B; B = 16'h00D7; #100;
A = 16'h001B; B = 16'h00D8; #100;
A = 16'h001B; B = 16'h00D9; #100;
A = 16'h001B; B = 16'h00DA; #100;
A = 16'h001B; B = 16'h00DB; #100;
A = 16'h001B; B = 16'h00DC; #100;
A = 16'h001B; B = 16'h00DD; #100;
A = 16'h001B; B = 16'h00DE; #100;
A = 16'h001B; B = 16'h00DF; #100;
A = 16'h001B; B = 16'h00E0; #100;
A = 16'h001B; B = 16'h00E1; #100;
A = 16'h001B; B = 16'h00E2; #100;
A = 16'h001B; B = 16'h00E3; #100;
A = 16'h001B; B = 16'h00E4; #100;
A = 16'h001B; B = 16'h00E5; #100;
A = 16'h001B; B = 16'h00E6; #100;
A = 16'h001B; B = 16'h00E7; #100;
A = 16'h001B; B = 16'h00E8; #100;
A = 16'h001B; B = 16'h00E9; #100;
A = 16'h001B; B = 16'h00EA; #100;
A = 16'h001B; B = 16'h00EB; #100;
A = 16'h001B; B = 16'h00EC; #100;
A = 16'h001B; B = 16'h00ED; #100;
A = 16'h001B; B = 16'h00EE; #100;
A = 16'h001B; B = 16'h00EF; #100;
A = 16'h001B; B = 16'h00F0; #100;
A = 16'h001B; B = 16'h00F1; #100;
A = 16'h001B; B = 16'h00F2; #100;
A = 16'h001B; B = 16'h00F3; #100;
A = 16'h001B; B = 16'h00F4; #100;
A = 16'h001B; B = 16'h00F5; #100;
A = 16'h001B; B = 16'h00F6; #100;
A = 16'h001B; B = 16'h00F7; #100;
A = 16'h001B; B = 16'h00F8; #100;
A = 16'h001B; B = 16'h00F9; #100;
A = 16'h001B; B = 16'h00FA; #100;
A = 16'h001B; B = 16'h00FB; #100;
A = 16'h001B; B = 16'h00FC; #100;
A = 16'h001B; B = 16'h00FD; #100;
A = 16'h001B; B = 16'h00FE; #100;
A = 16'h001B; B = 16'h00FF; #100;
A = 16'h001C; B = 16'h000; #100;
A = 16'h001C; B = 16'h001; #100;
A = 16'h001C; B = 16'h002; #100;
A = 16'h001C; B = 16'h003; #100;
A = 16'h001C; B = 16'h004; #100;
A = 16'h001C; B = 16'h005; #100;
A = 16'h001C; B = 16'h006; #100;
A = 16'h001C; B = 16'h007; #100;
A = 16'h001C; B = 16'h008; #100;
A = 16'h001C; B = 16'h009; #100;
A = 16'h001C; B = 16'h00A; #100;
A = 16'h001C; B = 16'h00B; #100;
A = 16'h001C; B = 16'h00C; #100;
A = 16'h001C; B = 16'h00D; #100;
A = 16'h001C; B = 16'h00E; #100;
A = 16'h001C; B = 16'h00F; #100;
A = 16'h001C; B = 16'h0010; #100;
A = 16'h001C; B = 16'h0011; #100;
A = 16'h001C; B = 16'h0012; #100;
A = 16'h001C; B = 16'h0013; #100;
A = 16'h001C; B = 16'h0014; #100;
A = 16'h001C; B = 16'h0015; #100;
A = 16'h001C; B = 16'h0016; #100;
A = 16'h001C; B = 16'h0017; #100;
A = 16'h001C; B = 16'h0018; #100;
A = 16'h001C; B = 16'h0019; #100;
A = 16'h001C; B = 16'h001A; #100;
A = 16'h001C; B = 16'h001B; #100;
A = 16'h001C; B = 16'h001C; #100;
A = 16'h001C; B = 16'h001D; #100;
A = 16'h001C; B = 16'h001E; #100;
A = 16'h001C; B = 16'h001F; #100;
A = 16'h001C; B = 16'h0020; #100;
A = 16'h001C; B = 16'h0021; #100;
A = 16'h001C; B = 16'h0022; #100;
A = 16'h001C; B = 16'h0023; #100;
A = 16'h001C; B = 16'h0024; #100;
A = 16'h001C; B = 16'h0025; #100;
A = 16'h001C; B = 16'h0026; #100;
A = 16'h001C; B = 16'h0027; #100;
A = 16'h001C; B = 16'h0028; #100;
A = 16'h001C; B = 16'h0029; #100;
A = 16'h001C; B = 16'h002A; #100;
A = 16'h001C; B = 16'h002B; #100;
A = 16'h001C; B = 16'h002C; #100;
A = 16'h001C; B = 16'h002D; #100;
A = 16'h001C; B = 16'h002E; #100;
A = 16'h001C; B = 16'h002F; #100;
A = 16'h001C; B = 16'h0030; #100;
A = 16'h001C; B = 16'h0031; #100;
A = 16'h001C; B = 16'h0032; #100;
A = 16'h001C; B = 16'h0033; #100;
A = 16'h001C; B = 16'h0034; #100;
A = 16'h001C; B = 16'h0035; #100;
A = 16'h001C; B = 16'h0036; #100;
A = 16'h001C; B = 16'h0037; #100;
A = 16'h001C; B = 16'h0038; #100;
A = 16'h001C; B = 16'h0039; #100;
A = 16'h001C; B = 16'h003A; #100;
A = 16'h001C; B = 16'h003B; #100;
A = 16'h001C; B = 16'h003C; #100;
A = 16'h001C; B = 16'h003D; #100;
A = 16'h001C; B = 16'h003E; #100;
A = 16'h001C; B = 16'h003F; #100;
A = 16'h001C; B = 16'h0040; #100;
A = 16'h001C; B = 16'h0041; #100;
A = 16'h001C; B = 16'h0042; #100;
A = 16'h001C; B = 16'h0043; #100;
A = 16'h001C; B = 16'h0044; #100;
A = 16'h001C; B = 16'h0045; #100;
A = 16'h001C; B = 16'h0046; #100;
A = 16'h001C; B = 16'h0047; #100;
A = 16'h001C; B = 16'h0048; #100;
A = 16'h001C; B = 16'h0049; #100;
A = 16'h001C; B = 16'h004A; #100;
A = 16'h001C; B = 16'h004B; #100;
A = 16'h001C; B = 16'h004C; #100;
A = 16'h001C; B = 16'h004D; #100;
A = 16'h001C; B = 16'h004E; #100;
A = 16'h001C; B = 16'h004F; #100;
A = 16'h001C; B = 16'h0050; #100;
A = 16'h001C; B = 16'h0051; #100;
A = 16'h001C; B = 16'h0052; #100;
A = 16'h001C; B = 16'h0053; #100;
A = 16'h001C; B = 16'h0054; #100;
A = 16'h001C; B = 16'h0055; #100;
A = 16'h001C; B = 16'h0056; #100;
A = 16'h001C; B = 16'h0057; #100;
A = 16'h001C; B = 16'h0058; #100;
A = 16'h001C; B = 16'h0059; #100;
A = 16'h001C; B = 16'h005A; #100;
A = 16'h001C; B = 16'h005B; #100;
A = 16'h001C; B = 16'h005C; #100;
A = 16'h001C; B = 16'h005D; #100;
A = 16'h001C; B = 16'h005E; #100;
A = 16'h001C; B = 16'h005F; #100;
A = 16'h001C; B = 16'h0060; #100;
A = 16'h001C; B = 16'h0061; #100;
A = 16'h001C; B = 16'h0062; #100;
A = 16'h001C; B = 16'h0063; #100;
A = 16'h001C; B = 16'h0064; #100;
A = 16'h001C; B = 16'h0065; #100;
A = 16'h001C; B = 16'h0066; #100;
A = 16'h001C; B = 16'h0067; #100;
A = 16'h001C; B = 16'h0068; #100;
A = 16'h001C; B = 16'h0069; #100;
A = 16'h001C; B = 16'h006A; #100;
A = 16'h001C; B = 16'h006B; #100;
A = 16'h001C; B = 16'h006C; #100;
A = 16'h001C; B = 16'h006D; #100;
A = 16'h001C; B = 16'h006E; #100;
A = 16'h001C; B = 16'h006F; #100;
A = 16'h001C; B = 16'h0070; #100;
A = 16'h001C; B = 16'h0071; #100;
A = 16'h001C; B = 16'h0072; #100;
A = 16'h001C; B = 16'h0073; #100;
A = 16'h001C; B = 16'h0074; #100;
A = 16'h001C; B = 16'h0075; #100;
A = 16'h001C; B = 16'h0076; #100;
A = 16'h001C; B = 16'h0077; #100;
A = 16'h001C; B = 16'h0078; #100;
A = 16'h001C; B = 16'h0079; #100;
A = 16'h001C; B = 16'h007A; #100;
A = 16'h001C; B = 16'h007B; #100;
A = 16'h001C; B = 16'h007C; #100;
A = 16'h001C; B = 16'h007D; #100;
A = 16'h001C; B = 16'h007E; #100;
A = 16'h001C; B = 16'h007F; #100;
A = 16'h001C; B = 16'h0080; #100;
A = 16'h001C; B = 16'h0081; #100;
A = 16'h001C; B = 16'h0082; #100;
A = 16'h001C; B = 16'h0083; #100;
A = 16'h001C; B = 16'h0084; #100;
A = 16'h001C; B = 16'h0085; #100;
A = 16'h001C; B = 16'h0086; #100;
A = 16'h001C; B = 16'h0087; #100;
A = 16'h001C; B = 16'h0088; #100;
A = 16'h001C; B = 16'h0089; #100;
A = 16'h001C; B = 16'h008A; #100;
A = 16'h001C; B = 16'h008B; #100;
A = 16'h001C; B = 16'h008C; #100;
A = 16'h001C; B = 16'h008D; #100;
A = 16'h001C; B = 16'h008E; #100;
A = 16'h001C; B = 16'h008F; #100;
A = 16'h001C; B = 16'h0090; #100;
A = 16'h001C; B = 16'h0091; #100;
A = 16'h001C; B = 16'h0092; #100;
A = 16'h001C; B = 16'h0093; #100;
A = 16'h001C; B = 16'h0094; #100;
A = 16'h001C; B = 16'h0095; #100;
A = 16'h001C; B = 16'h0096; #100;
A = 16'h001C; B = 16'h0097; #100;
A = 16'h001C; B = 16'h0098; #100;
A = 16'h001C; B = 16'h0099; #100;
A = 16'h001C; B = 16'h009A; #100;
A = 16'h001C; B = 16'h009B; #100;
A = 16'h001C; B = 16'h009C; #100;
A = 16'h001C; B = 16'h009D; #100;
A = 16'h001C; B = 16'h009E; #100;
A = 16'h001C; B = 16'h009F; #100;
A = 16'h001C; B = 16'h00A0; #100;
A = 16'h001C; B = 16'h00A1; #100;
A = 16'h001C; B = 16'h00A2; #100;
A = 16'h001C; B = 16'h00A3; #100;
A = 16'h001C; B = 16'h00A4; #100;
A = 16'h001C; B = 16'h00A5; #100;
A = 16'h001C; B = 16'h00A6; #100;
A = 16'h001C; B = 16'h00A7; #100;
A = 16'h001C; B = 16'h00A8; #100;
A = 16'h001C; B = 16'h00A9; #100;
A = 16'h001C; B = 16'h00AA; #100;
A = 16'h001C; B = 16'h00AB; #100;
A = 16'h001C; B = 16'h00AC; #100;
A = 16'h001C; B = 16'h00AD; #100;
A = 16'h001C; B = 16'h00AE; #100;
A = 16'h001C; B = 16'h00AF; #100;
A = 16'h001C; B = 16'h00B0; #100;
A = 16'h001C; B = 16'h00B1; #100;
A = 16'h001C; B = 16'h00B2; #100;
A = 16'h001C; B = 16'h00B3; #100;
A = 16'h001C; B = 16'h00B4; #100;
A = 16'h001C; B = 16'h00B5; #100;
A = 16'h001C; B = 16'h00B6; #100;
A = 16'h001C; B = 16'h00B7; #100;
A = 16'h001C; B = 16'h00B8; #100;
A = 16'h001C; B = 16'h00B9; #100;
A = 16'h001C; B = 16'h00BA; #100;
A = 16'h001C; B = 16'h00BB; #100;
A = 16'h001C; B = 16'h00BC; #100;
A = 16'h001C; B = 16'h00BD; #100;
A = 16'h001C; B = 16'h00BE; #100;
A = 16'h001C; B = 16'h00BF; #100;
A = 16'h001C; B = 16'h00C0; #100;
A = 16'h001C; B = 16'h00C1; #100;
A = 16'h001C; B = 16'h00C2; #100;
A = 16'h001C; B = 16'h00C3; #100;
A = 16'h001C; B = 16'h00C4; #100;
A = 16'h001C; B = 16'h00C5; #100;
A = 16'h001C; B = 16'h00C6; #100;
A = 16'h001C; B = 16'h00C7; #100;
A = 16'h001C; B = 16'h00C8; #100;
A = 16'h001C; B = 16'h00C9; #100;
A = 16'h001C; B = 16'h00CA; #100;
A = 16'h001C; B = 16'h00CB; #100;
A = 16'h001C; B = 16'h00CC; #100;
A = 16'h001C; B = 16'h00CD; #100;
A = 16'h001C; B = 16'h00CE; #100;
A = 16'h001C; B = 16'h00CF; #100;
A = 16'h001C; B = 16'h00D0; #100;
A = 16'h001C; B = 16'h00D1; #100;
A = 16'h001C; B = 16'h00D2; #100;
A = 16'h001C; B = 16'h00D3; #100;
A = 16'h001C; B = 16'h00D4; #100;
A = 16'h001C; B = 16'h00D5; #100;
A = 16'h001C; B = 16'h00D6; #100;
A = 16'h001C; B = 16'h00D7; #100;
A = 16'h001C; B = 16'h00D8; #100;
A = 16'h001C; B = 16'h00D9; #100;
A = 16'h001C; B = 16'h00DA; #100;
A = 16'h001C; B = 16'h00DB; #100;
A = 16'h001C; B = 16'h00DC; #100;
A = 16'h001C; B = 16'h00DD; #100;
A = 16'h001C; B = 16'h00DE; #100;
A = 16'h001C; B = 16'h00DF; #100;
A = 16'h001C; B = 16'h00E0; #100;
A = 16'h001C; B = 16'h00E1; #100;
A = 16'h001C; B = 16'h00E2; #100;
A = 16'h001C; B = 16'h00E3; #100;
A = 16'h001C; B = 16'h00E4; #100;
A = 16'h001C; B = 16'h00E5; #100;
A = 16'h001C; B = 16'h00E6; #100;
A = 16'h001C; B = 16'h00E7; #100;
A = 16'h001C; B = 16'h00E8; #100;
A = 16'h001C; B = 16'h00E9; #100;
A = 16'h001C; B = 16'h00EA; #100;
A = 16'h001C; B = 16'h00EB; #100;
A = 16'h001C; B = 16'h00EC; #100;
A = 16'h001C; B = 16'h00ED; #100;
A = 16'h001C; B = 16'h00EE; #100;
A = 16'h001C; B = 16'h00EF; #100;
A = 16'h001C; B = 16'h00F0; #100;
A = 16'h001C; B = 16'h00F1; #100;
A = 16'h001C; B = 16'h00F2; #100;
A = 16'h001C; B = 16'h00F3; #100;
A = 16'h001C; B = 16'h00F4; #100;
A = 16'h001C; B = 16'h00F5; #100;
A = 16'h001C; B = 16'h00F6; #100;
A = 16'h001C; B = 16'h00F7; #100;
A = 16'h001C; B = 16'h00F8; #100;
A = 16'h001C; B = 16'h00F9; #100;
A = 16'h001C; B = 16'h00FA; #100;
A = 16'h001C; B = 16'h00FB; #100;
A = 16'h001C; B = 16'h00FC; #100;
A = 16'h001C; B = 16'h00FD; #100;
A = 16'h001C; B = 16'h00FE; #100;
A = 16'h001C; B = 16'h00FF; #100;
A = 16'h001D; B = 16'h000; #100;
A = 16'h001D; B = 16'h001; #100;
A = 16'h001D; B = 16'h002; #100;
A = 16'h001D; B = 16'h003; #100;
A = 16'h001D; B = 16'h004; #100;
A = 16'h001D; B = 16'h005; #100;
A = 16'h001D; B = 16'h006; #100;
A = 16'h001D; B = 16'h007; #100;
A = 16'h001D; B = 16'h008; #100;
A = 16'h001D; B = 16'h009; #100;
A = 16'h001D; B = 16'h00A; #100;
A = 16'h001D; B = 16'h00B; #100;
A = 16'h001D; B = 16'h00C; #100;
A = 16'h001D; B = 16'h00D; #100;
A = 16'h001D; B = 16'h00E; #100;
A = 16'h001D; B = 16'h00F; #100;
A = 16'h001D; B = 16'h0010; #100;
A = 16'h001D; B = 16'h0011; #100;
A = 16'h001D; B = 16'h0012; #100;
A = 16'h001D; B = 16'h0013; #100;
A = 16'h001D; B = 16'h0014; #100;
A = 16'h001D; B = 16'h0015; #100;
A = 16'h001D; B = 16'h0016; #100;
A = 16'h001D; B = 16'h0017; #100;
A = 16'h001D; B = 16'h0018; #100;
A = 16'h001D; B = 16'h0019; #100;
A = 16'h001D; B = 16'h001A; #100;
A = 16'h001D; B = 16'h001B; #100;
A = 16'h001D; B = 16'h001C; #100;
A = 16'h001D; B = 16'h001D; #100;
A = 16'h001D; B = 16'h001E; #100;
A = 16'h001D; B = 16'h001F; #100;
A = 16'h001D; B = 16'h0020; #100;
A = 16'h001D; B = 16'h0021; #100;
A = 16'h001D; B = 16'h0022; #100;
A = 16'h001D; B = 16'h0023; #100;
A = 16'h001D; B = 16'h0024; #100;
A = 16'h001D; B = 16'h0025; #100;
A = 16'h001D; B = 16'h0026; #100;
A = 16'h001D; B = 16'h0027; #100;
A = 16'h001D; B = 16'h0028; #100;
A = 16'h001D; B = 16'h0029; #100;
A = 16'h001D; B = 16'h002A; #100;
A = 16'h001D; B = 16'h002B; #100;
A = 16'h001D; B = 16'h002C; #100;
A = 16'h001D; B = 16'h002D; #100;
A = 16'h001D; B = 16'h002E; #100;
A = 16'h001D; B = 16'h002F; #100;
A = 16'h001D; B = 16'h0030; #100;
A = 16'h001D; B = 16'h0031; #100;
A = 16'h001D; B = 16'h0032; #100;
A = 16'h001D; B = 16'h0033; #100;
A = 16'h001D; B = 16'h0034; #100;
A = 16'h001D; B = 16'h0035; #100;
A = 16'h001D; B = 16'h0036; #100;
A = 16'h001D; B = 16'h0037; #100;
A = 16'h001D; B = 16'h0038; #100;
A = 16'h001D; B = 16'h0039; #100;
A = 16'h001D; B = 16'h003A; #100;
A = 16'h001D; B = 16'h003B; #100;
A = 16'h001D; B = 16'h003C; #100;
A = 16'h001D; B = 16'h003D; #100;
A = 16'h001D; B = 16'h003E; #100;
A = 16'h001D; B = 16'h003F; #100;
A = 16'h001D; B = 16'h0040; #100;
A = 16'h001D; B = 16'h0041; #100;
A = 16'h001D; B = 16'h0042; #100;
A = 16'h001D; B = 16'h0043; #100;
A = 16'h001D; B = 16'h0044; #100;
A = 16'h001D; B = 16'h0045; #100;
A = 16'h001D; B = 16'h0046; #100;
A = 16'h001D; B = 16'h0047; #100;
A = 16'h001D; B = 16'h0048; #100;
A = 16'h001D; B = 16'h0049; #100;
A = 16'h001D; B = 16'h004A; #100;
A = 16'h001D; B = 16'h004B; #100;
A = 16'h001D; B = 16'h004C; #100;
A = 16'h001D; B = 16'h004D; #100;
A = 16'h001D; B = 16'h004E; #100;
A = 16'h001D; B = 16'h004F; #100;
A = 16'h001D; B = 16'h0050; #100;
A = 16'h001D; B = 16'h0051; #100;
A = 16'h001D; B = 16'h0052; #100;
A = 16'h001D; B = 16'h0053; #100;
A = 16'h001D; B = 16'h0054; #100;
A = 16'h001D; B = 16'h0055; #100;
A = 16'h001D; B = 16'h0056; #100;
A = 16'h001D; B = 16'h0057; #100;
A = 16'h001D; B = 16'h0058; #100;
A = 16'h001D; B = 16'h0059; #100;
A = 16'h001D; B = 16'h005A; #100;
A = 16'h001D; B = 16'h005B; #100;
A = 16'h001D; B = 16'h005C; #100;
A = 16'h001D; B = 16'h005D; #100;
A = 16'h001D; B = 16'h005E; #100;
A = 16'h001D; B = 16'h005F; #100;
A = 16'h001D; B = 16'h0060; #100;
A = 16'h001D; B = 16'h0061; #100;
A = 16'h001D; B = 16'h0062; #100;
A = 16'h001D; B = 16'h0063; #100;
A = 16'h001D; B = 16'h0064; #100;
A = 16'h001D; B = 16'h0065; #100;
A = 16'h001D; B = 16'h0066; #100;
A = 16'h001D; B = 16'h0067; #100;
A = 16'h001D; B = 16'h0068; #100;
A = 16'h001D; B = 16'h0069; #100;
A = 16'h001D; B = 16'h006A; #100;
A = 16'h001D; B = 16'h006B; #100;
A = 16'h001D; B = 16'h006C; #100;
A = 16'h001D; B = 16'h006D; #100;
A = 16'h001D; B = 16'h006E; #100;
A = 16'h001D; B = 16'h006F; #100;
A = 16'h001D; B = 16'h0070; #100;
A = 16'h001D; B = 16'h0071; #100;
A = 16'h001D; B = 16'h0072; #100;
A = 16'h001D; B = 16'h0073; #100;
A = 16'h001D; B = 16'h0074; #100;
A = 16'h001D; B = 16'h0075; #100;
A = 16'h001D; B = 16'h0076; #100;
A = 16'h001D; B = 16'h0077; #100;
A = 16'h001D; B = 16'h0078; #100;
A = 16'h001D; B = 16'h0079; #100;
A = 16'h001D; B = 16'h007A; #100;
A = 16'h001D; B = 16'h007B; #100;
A = 16'h001D; B = 16'h007C; #100;
A = 16'h001D; B = 16'h007D; #100;
A = 16'h001D; B = 16'h007E; #100;
A = 16'h001D; B = 16'h007F; #100;
A = 16'h001D; B = 16'h0080; #100;
A = 16'h001D; B = 16'h0081; #100;
A = 16'h001D; B = 16'h0082; #100;
A = 16'h001D; B = 16'h0083; #100;
A = 16'h001D; B = 16'h0084; #100;
A = 16'h001D; B = 16'h0085; #100;
A = 16'h001D; B = 16'h0086; #100;
A = 16'h001D; B = 16'h0087; #100;
A = 16'h001D; B = 16'h0088; #100;
A = 16'h001D; B = 16'h0089; #100;
A = 16'h001D; B = 16'h008A; #100;
A = 16'h001D; B = 16'h008B; #100;
A = 16'h001D; B = 16'h008C; #100;
A = 16'h001D; B = 16'h008D; #100;
A = 16'h001D; B = 16'h008E; #100;
A = 16'h001D; B = 16'h008F; #100;
A = 16'h001D; B = 16'h0090; #100;
A = 16'h001D; B = 16'h0091; #100;
A = 16'h001D; B = 16'h0092; #100;
A = 16'h001D; B = 16'h0093; #100;
A = 16'h001D; B = 16'h0094; #100;
A = 16'h001D; B = 16'h0095; #100;
A = 16'h001D; B = 16'h0096; #100;
A = 16'h001D; B = 16'h0097; #100;
A = 16'h001D; B = 16'h0098; #100;
A = 16'h001D; B = 16'h0099; #100;
A = 16'h001D; B = 16'h009A; #100;
A = 16'h001D; B = 16'h009B; #100;
A = 16'h001D; B = 16'h009C; #100;
A = 16'h001D; B = 16'h009D; #100;
A = 16'h001D; B = 16'h009E; #100;
A = 16'h001D; B = 16'h009F; #100;
A = 16'h001D; B = 16'h00A0; #100;
A = 16'h001D; B = 16'h00A1; #100;
A = 16'h001D; B = 16'h00A2; #100;
A = 16'h001D; B = 16'h00A3; #100;
A = 16'h001D; B = 16'h00A4; #100;
A = 16'h001D; B = 16'h00A5; #100;
A = 16'h001D; B = 16'h00A6; #100;
A = 16'h001D; B = 16'h00A7; #100;
A = 16'h001D; B = 16'h00A8; #100;
A = 16'h001D; B = 16'h00A9; #100;
A = 16'h001D; B = 16'h00AA; #100;
A = 16'h001D; B = 16'h00AB; #100;
A = 16'h001D; B = 16'h00AC; #100;
A = 16'h001D; B = 16'h00AD; #100;
A = 16'h001D; B = 16'h00AE; #100;
A = 16'h001D; B = 16'h00AF; #100;
A = 16'h001D; B = 16'h00B0; #100;
A = 16'h001D; B = 16'h00B1; #100;
A = 16'h001D; B = 16'h00B2; #100;
A = 16'h001D; B = 16'h00B3; #100;
A = 16'h001D; B = 16'h00B4; #100;
A = 16'h001D; B = 16'h00B5; #100;
A = 16'h001D; B = 16'h00B6; #100;
A = 16'h001D; B = 16'h00B7; #100;
A = 16'h001D; B = 16'h00B8; #100;
A = 16'h001D; B = 16'h00B9; #100;
A = 16'h001D; B = 16'h00BA; #100;
A = 16'h001D; B = 16'h00BB; #100;
A = 16'h001D; B = 16'h00BC; #100;
A = 16'h001D; B = 16'h00BD; #100;
A = 16'h001D; B = 16'h00BE; #100;
A = 16'h001D; B = 16'h00BF; #100;
A = 16'h001D; B = 16'h00C0; #100;
A = 16'h001D; B = 16'h00C1; #100;
A = 16'h001D; B = 16'h00C2; #100;
A = 16'h001D; B = 16'h00C3; #100;
A = 16'h001D; B = 16'h00C4; #100;
A = 16'h001D; B = 16'h00C5; #100;
A = 16'h001D; B = 16'h00C6; #100;
A = 16'h001D; B = 16'h00C7; #100;
A = 16'h001D; B = 16'h00C8; #100;
A = 16'h001D; B = 16'h00C9; #100;
A = 16'h001D; B = 16'h00CA; #100;
A = 16'h001D; B = 16'h00CB; #100;
A = 16'h001D; B = 16'h00CC; #100;
A = 16'h001D; B = 16'h00CD; #100;
A = 16'h001D; B = 16'h00CE; #100;
A = 16'h001D; B = 16'h00CF; #100;
A = 16'h001D; B = 16'h00D0; #100;
A = 16'h001D; B = 16'h00D1; #100;
A = 16'h001D; B = 16'h00D2; #100;
A = 16'h001D; B = 16'h00D3; #100;
A = 16'h001D; B = 16'h00D4; #100;
A = 16'h001D; B = 16'h00D5; #100;
A = 16'h001D; B = 16'h00D6; #100;
A = 16'h001D; B = 16'h00D7; #100;
A = 16'h001D; B = 16'h00D8; #100;
A = 16'h001D; B = 16'h00D9; #100;
A = 16'h001D; B = 16'h00DA; #100;
A = 16'h001D; B = 16'h00DB; #100;
A = 16'h001D; B = 16'h00DC; #100;
A = 16'h001D; B = 16'h00DD; #100;
A = 16'h001D; B = 16'h00DE; #100;
A = 16'h001D; B = 16'h00DF; #100;
A = 16'h001D; B = 16'h00E0; #100;
A = 16'h001D; B = 16'h00E1; #100;
A = 16'h001D; B = 16'h00E2; #100;
A = 16'h001D; B = 16'h00E3; #100;
A = 16'h001D; B = 16'h00E4; #100;
A = 16'h001D; B = 16'h00E5; #100;
A = 16'h001D; B = 16'h00E6; #100;
A = 16'h001D; B = 16'h00E7; #100;
A = 16'h001D; B = 16'h00E8; #100;
A = 16'h001D; B = 16'h00E9; #100;
A = 16'h001D; B = 16'h00EA; #100;
A = 16'h001D; B = 16'h00EB; #100;
A = 16'h001D; B = 16'h00EC; #100;
A = 16'h001D; B = 16'h00ED; #100;
A = 16'h001D; B = 16'h00EE; #100;
A = 16'h001D; B = 16'h00EF; #100;
A = 16'h001D; B = 16'h00F0; #100;
A = 16'h001D; B = 16'h00F1; #100;
A = 16'h001D; B = 16'h00F2; #100;
A = 16'h001D; B = 16'h00F3; #100;
A = 16'h001D; B = 16'h00F4; #100;
A = 16'h001D; B = 16'h00F5; #100;
A = 16'h001D; B = 16'h00F6; #100;
A = 16'h001D; B = 16'h00F7; #100;
A = 16'h001D; B = 16'h00F8; #100;
A = 16'h001D; B = 16'h00F9; #100;
A = 16'h001D; B = 16'h00FA; #100;
A = 16'h001D; B = 16'h00FB; #100;
A = 16'h001D; B = 16'h00FC; #100;
A = 16'h001D; B = 16'h00FD; #100;
A = 16'h001D; B = 16'h00FE; #100;
A = 16'h001D; B = 16'h00FF; #100;
A = 16'h001E; B = 16'h000; #100;
A = 16'h001E; B = 16'h001; #100;
A = 16'h001E; B = 16'h002; #100;
A = 16'h001E; B = 16'h003; #100;
A = 16'h001E; B = 16'h004; #100;
A = 16'h001E; B = 16'h005; #100;
A = 16'h001E; B = 16'h006; #100;
A = 16'h001E; B = 16'h007; #100;
A = 16'h001E; B = 16'h008; #100;
A = 16'h001E; B = 16'h009; #100;
A = 16'h001E; B = 16'h00A; #100;
A = 16'h001E; B = 16'h00B; #100;
A = 16'h001E; B = 16'h00C; #100;
A = 16'h001E; B = 16'h00D; #100;
A = 16'h001E; B = 16'h00E; #100;
A = 16'h001E; B = 16'h00F; #100;
A = 16'h001E; B = 16'h0010; #100;
A = 16'h001E; B = 16'h0011; #100;
A = 16'h001E; B = 16'h0012; #100;
A = 16'h001E; B = 16'h0013; #100;
A = 16'h001E; B = 16'h0014; #100;
A = 16'h001E; B = 16'h0015; #100;
A = 16'h001E; B = 16'h0016; #100;
A = 16'h001E; B = 16'h0017; #100;
A = 16'h001E; B = 16'h0018; #100;
A = 16'h001E; B = 16'h0019; #100;
A = 16'h001E; B = 16'h001A; #100;
A = 16'h001E; B = 16'h001B; #100;
A = 16'h001E; B = 16'h001C; #100;
A = 16'h001E; B = 16'h001D; #100;
A = 16'h001E; B = 16'h001E; #100;
A = 16'h001E; B = 16'h001F; #100;
A = 16'h001E; B = 16'h0020; #100;
A = 16'h001E; B = 16'h0021; #100;
A = 16'h001E; B = 16'h0022; #100;
A = 16'h001E; B = 16'h0023; #100;
A = 16'h001E; B = 16'h0024; #100;
A = 16'h001E; B = 16'h0025; #100;
A = 16'h001E; B = 16'h0026; #100;
A = 16'h001E; B = 16'h0027; #100;
A = 16'h001E; B = 16'h0028; #100;
A = 16'h001E; B = 16'h0029; #100;
A = 16'h001E; B = 16'h002A; #100;
A = 16'h001E; B = 16'h002B; #100;
A = 16'h001E; B = 16'h002C; #100;
A = 16'h001E; B = 16'h002D; #100;
A = 16'h001E; B = 16'h002E; #100;
A = 16'h001E; B = 16'h002F; #100;
A = 16'h001E; B = 16'h0030; #100;
A = 16'h001E; B = 16'h0031; #100;
A = 16'h001E; B = 16'h0032; #100;
A = 16'h001E; B = 16'h0033; #100;
A = 16'h001E; B = 16'h0034; #100;
A = 16'h001E; B = 16'h0035; #100;
A = 16'h001E; B = 16'h0036; #100;
A = 16'h001E; B = 16'h0037; #100;
A = 16'h001E; B = 16'h0038; #100;
A = 16'h001E; B = 16'h0039; #100;
A = 16'h001E; B = 16'h003A; #100;
A = 16'h001E; B = 16'h003B; #100;
A = 16'h001E; B = 16'h003C; #100;
A = 16'h001E; B = 16'h003D; #100;
A = 16'h001E; B = 16'h003E; #100;
A = 16'h001E; B = 16'h003F; #100;
A = 16'h001E; B = 16'h0040; #100;
A = 16'h001E; B = 16'h0041; #100;
A = 16'h001E; B = 16'h0042; #100;
A = 16'h001E; B = 16'h0043; #100;
A = 16'h001E; B = 16'h0044; #100;
A = 16'h001E; B = 16'h0045; #100;
A = 16'h001E; B = 16'h0046; #100;
A = 16'h001E; B = 16'h0047; #100;
A = 16'h001E; B = 16'h0048; #100;
A = 16'h001E; B = 16'h0049; #100;
A = 16'h001E; B = 16'h004A; #100;
A = 16'h001E; B = 16'h004B; #100;
A = 16'h001E; B = 16'h004C; #100;
A = 16'h001E; B = 16'h004D; #100;
A = 16'h001E; B = 16'h004E; #100;
A = 16'h001E; B = 16'h004F; #100;
A = 16'h001E; B = 16'h0050; #100;
A = 16'h001E; B = 16'h0051; #100;
A = 16'h001E; B = 16'h0052; #100;
A = 16'h001E; B = 16'h0053; #100;
A = 16'h001E; B = 16'h0054; #100;
A = 16'h001E; B = 16'h0055; #100;
A = 16'h001E; B = 16'h0056; #100;
A = 16'h001E; B = 16'h0057; #100;
A = 16'h001E; B = 16'h0058; #100;
A = 16'h001E; B = 16'h0059; #100;
A = 16'h001E; B = 16'h005A; #100;
A = 16'h001E; B = 16'h005B; #100;
A = 16'h001E; B = 16'h005C; #100;
A = 16'h001E; B = 16'h005D; #100;
A = 16'h001E; B = 16'h005E; #100;
A = 16'h001E; B = 16'h005F; #100;
A = 16'h001E; B = 16'h0060; #100;
A = 16'h001E; B = 16'h0061; #100;
A = 16'h001E; B = 16'h0062; #100;
A = 16'h001E; B = 16'h0063; #100;
A = 16'h001E; B = 16'h0064; #100;
A = 16'h001E; B = 16'h0065; #100;
A = 16'h001E; B = 16'h0066; #100;
A = 16'h001E; B = 16'h0067; #100;
A = 16'h001E; B = 16'h0068; #100;
A = 16'h001E; B = 16'h0069; #100;
A = 16'h001E; B = 16'h006A; #100;
A = 16'h001E; B = 16'h006B; #100;
A = 16'h001E; B = 16'h006C; #100;
A = 16'h001E; B = 16'h006D; #100;
A = 16'h001E; B = 16'h006E; #100;
A = 16'h001E; B = 16'h006F; #100;
A = 16'h001E; B = 16'h0070; #100;
A = 16'h001E; B = 16'h0071; #100;
A = 16'h001E; B = 16'h0072; #100;
A = 16'h001E; B = 16'h0073; #100;
A = 16'h001E; B = 16'h0074; #100;
A = 16'h001E; B = 16'h0075; #100;
A = 16'h001E; B = 16'h0076; #100;
A = 16'h001E; B = 16'h0077; #100;
A = 16'h001E; B = 16'h0078; #100;
A = 16'h001E; B = 16'h0079; #100;
A = 16'h001E; B = 16'h007A; #100;
A = 16'h001E; B = 16'h007B; #100;
A = 16'h001E; B = 16'h007C; #100;
A = 16'h001E; B = 16'h007D; #100;
A = 16'h001E; B = 16'h007E; #100;
A = 16'h001E; B = 16'h007F; #100;
A = 16'h001E; B = 16'h0080; #100;
A = 16'h001E; B = 16'h0081; #100;
A = 16'h001E; B = 16'h0082; #100;
A = 16'h001E; B = 16'h0083; #100;
A = 16'h001E; B = 16'h0084; #100;
A = 16'h001E; B = 16'h0085; #100;
A = 16'h001E; B = 16'h0086; #100;
A = 16'h001E; B = 16'h0087; #100;
A = 16'h001E; B = 16'h0088; #100;
A = 16'h001E; B = 16'h0089; #100;
A = 16'h001E; B = 16'h008A; #100;
A = 16'h001E; B = 16'h008B; #100;
A = 16'h001E; B = 16'h008C; #100;
A = 16'h001E; B = 16'h008D; #100;
A = 16'h001E; B = 16'h008E; #100;
A = 16'h001E; B = 16'h008F; #100;
A = 16'h001E; B = 16'h0090; #100;
A = 16'h001E; B = 16'h0091; #100;
A = 16'h001E; B = 16'h0092; #100;
A = 16'h001E; B = 16'h0093; #100;
A = 16'h001E; B = 16'h0094; #100;
A = 16'h001E; B = 16'h0095; #100;
A = 16'h001E; B = 16'h0096; #100;
A = 16'h001E; B = 16'h0097; #100;
A = 16'h001E; B = 16'h0098; #100;
A = 16'h001E; B = 16'h0099; #100;
A = 16'h001E; B = 16'h009A; #100;
A = 16'h001E; B = 16'h009B; #100;
A = 16'h001E; B = 16'h009C; #100;
A = 16'h001E; B = 16'h009D; #100;
A = 16'h001E; B = 16'h009E; #100;
A = 16'h001E; B = 16'h009F; #100;
A = 16'h001E; B = 16'h00A0; #100;
A = 16'h001E; B = 16'h00A1; #100;
A = 16'h001E; B = 16'h00A2; #100;
A = 16'h001E; B = 16'h00A3; #100;
A = 16'h001E; B = 16'h00A4; #100;
A = 16'h001E; B = 16'h00A5; #100;
A = 16'h001E; B = 16'h00A6; #100;
A = 16'h001E; B = 16'h00A7; #100;
A = 16'h001E; B = 16'h00A8; #100;
A = 16'h001E; B = 16'h00A9; #100;
A = 16'h001E; B = 16'h00AA; #100;
A = 16'h001E; B = 16'h00AB; #100;
A = 16'h001E; B = 16'h00AC; #100;
A = 16'h001E; B = 16'h00AD; #100;
A = 16'h001E; B = 16'h00AE; #100;
A = 16'h001E; B = 16'h00AF; #100;
A = 16'h001E; B = 16'h00B0; #100;
A = 16'h001E; B = 16'h00B1; #100;
A = 16'h001E; B = 16'h00B2; #100;
A = 16'h001E; B = 16'h00B3; #100;
A = 16'h001E; B = 16'h00B4; #100;
A = 16'h001E; B = 16'h00B5; #100;
A = 16'h001E; B = 16'h00B6; #100;
A = 16'h001E; B = 16'h00B7; #100;
A = 16'h001E; B = 16'h00B8; #100;
A = 16'h001E; B = 16'h00B9; #100;
A = 16'h001E; B = 16'h00BA; #100;
A = 16'h001E; B = 16'h00BB; #100;
A = 16'h001E; B = 16'h00BC; #100;
A = 16'h001E; B = 16'h00BD; #100;
A = 16'h001E; B = 16'h00BE; #100;
A = 16'h001E; B = 16'h00BF; #100;
A = 16'h001E; B = 16'h00C0; #100;
A = 16'h001E; B = 16'h00C1; #100;
A = 16'h001E; B = 16'h00C2; #100;
A = 16'h001E; B = 16'h00C3; #100;
A = 16'h001E; B = 16'h00C4; #100;
A = 16'h001E; B = 16'h00C5; #100;
A = 16'h001E; B = 16'h00C6; #100;
A = 16'h001E; B = 16'h00C7; #100;
A = 16'h001E; B = 16'h00C8; #100;
A = 16'h001E; B = 16'h00C9; #100;
A = 16'h001E; B = 16'h00CA; #100;
A = 16'h001E; B = 16'h00CB; #100;
A = 16'h001E; B = 16'h00CC; #100;
A = 16'h001E; B = 16'h00CD; #100;
A = 16'h001E; B = 16'h00CE; #100;
A = 16'h001E; B = 16'h00CF; #100;
A = 16'h001E; B = 16'h00D0; #100;
A = 16'h001E; B = 16'h00D1; #100;
A = 16'h001E; B = 16'h00D2; #100;
A = 16'h001E; B = 16'h00D3; #100;
A = 16'h001E; B = 16'h00D4; #100;
A = 16'h001E; B = 16'h00D5; #100;
A = 16'h001E; B = 16'h00D6; #100;
A = 16'h001E; B = 16'h00D7; #100;
A = 16'h001E; B = 16'h00D8; #100;
A = 16'h001E; B = 16'h00D9; #100;
A = 16'h001E; B = 16'h00DA; #100;
A = 16'h001E; B = 16'h00DB; #100;
A = 16'h001E; B = 16'h00DC; #100;
A = 16'h001E; B = 16'h00DD; #100;
A = 16'h001E; B = 16'h00DE; #100;
A = 16'h001E; B = 16'h00DF; #100;
A = 16'h001E; B = 16'h00E0; #100;
A = 16'h001E; B = 16'h00E1; #100;
A = 16'h001E; B = 16'h00E2; #100;
A = 16'h001E; B = 16'h00E3; #100;
A = 16'h001E; B = 16'h00E4; #100;
A = 16'h001E; B = 16'h00E5; #100;
A = 16'h001E; B = 16'h00E6; #100;
A = 16'h001E; B = 16'h00E7; #100;
A = 16'h001E; B = 16'h00E8; #100;
A = 16'h001E; B = 16'h00E9; #100;
A = 16'h001E; B = 16'h00EA; #100;
A = 16'h001E; B = 16'h00EB; #100;
A = 16'h001E; B = 16'h00EC; #100;
A = 16'h001E; B = 16'h00ED; #100;
A = 16'h001E; B = 16'h00EE; #100;
A = 16'h001E; B = 16'h00EF; #100;
A = 16'h001E; B = 16'h00F0; #100;
A = 16'h001E; B = 16'h00F1; #100;
A = 16'h001E; B = 16'h00F2; #100;
A = 16'h001E; B = 16'h00F3; #100;
A = 16'h001E; B = 16'h00F4; #100;
A = 16'h001E; B = 16'h00F5; #100;
A = 16'h001E; B = 16'h00F6; #100;
A = 16'h001E; B = 16'h00F7; #100;
A = 16'h001E; B = 16'h00F8; #100;
A = 16'h001E; B = 16'h00F9; #100;
A = 16'h001E; B = 16'h00FA; #100;
A = 16'h001E; B = 16'h00FB; #100;
A = 16'h001E; B = 16'h00FC; #100;
A = 16'h001E; B = 16'h00FD; #100;
A = 16'h001E; B = 16'h00FE; #100;
A = 16'h001E; B = 16'h00FF; #100;
A = 16'h001F; B = 16'h000; #100;
A = 16'h001F; B = 16'h001; #100;
A = 16'h001F; B = 16'h002; #100;
A = 16'h001F; B = 16'h003; #100;
A = 16'h001F; B = 16'h004; #100;
A = 16'h001F; B = 16'h005; #100;
A = 16'h001F; B = 16'h006; #100;
A = 16'h001F; B = 16'h007; #100;
A = 16'h001F; B = 16'h008; #100;
A = 16'h001F; B = 16'h009; #100;
A = 16'h001F; B = 16'h00A; #100;
A = 16'h001F; B = 16'h00B; #100;
A = 16'h001F; B = 16'h00C; #100;
A = 16'h001F; B = 16'h00D; #100;
A = 16'h001F; B = 16'h00E; #100;
A = 16'h001F; B = 16'h00F; #100;
A = 16'h001F; B = 16'h0010; #100;
A = 16'h001F; B = 16'h0011; #100;
A = 16'h001F; B = 16'h0012; #100;
A = 16'h001F; B = 16'h0013; #100;
A = 16'h001F; B = 16'h0014; #100;
A = 16'h001F; B = 16'h0015; #100;
A = 16'h001F; B = 16'h0016; #100;
A = 16'h001F; B = 16'h0017; #100;
A = 16'h001F; B = 16'h0018; #100;
A = 16'h001F; B = 16'h0019; #100;
A = 16'h001F; B = 16'h001A; #100;
A = 16'h001F; B = 16'h001B; #100;
A = 16'h001F; B = 16'h001C; #100;
A = 16'h001F; B = 16'h001D; #100;
A = 16'h001F; B = 16'h001E; #100;
A = 16'h001F; B = 16'h001F; #100;
A = 16'h001F; B = 16'h0020; #100;
A = 16'h001F; B = 16'h0021; #100;
A = 16'h001F; B = 16'h0022; #100;
A = 16'h001F; B = 16'h0023; #100;
A = 16'h001F; B = 16'h0024; #100;
A = 16'h001F; B = 16'h0025; #100;
A = 16'h001F; B = 16'h0026; #100;
A = 16'h001F; B = 16'h0027; #100;
A = 16'h001F; B = 16'h0028; #100;
A = 16'h001F; B = 16'h0029; #100;
A = 16'h001F; B = 16'h002A; #100;
A = 16'h001F; B = 16'h002B; #100;
A = 16'h001F; B = 16'h002C; #100;
A = 16'h001F; B = 16'h002D; #100;
A = 16'h001F; B = 16'h002E; #100;
A = 16'h001F; B = 16'h002F; #100;
A = 16'h001F; B = 16'h0030; #100;
A = 16'h001F; B = 16'h0031; #100;
A = 16'h001F; B = 16'h0032; #100;
A = 16'h001F; B = 16'h0033; #100;
A = 16'h001F; B = 16'h0034; #100;
A = 16'h001F; B = 16'h0035; #100;
A = 16'h001F; B = 16'h0036; #100;
A = 16'h001F; B = 16'h0037; #100;
A = 16'h001F; B = 16'h0038; #100;
A = 16'h001F; B = 16'h0039; #100;
A = 16'h001F; B = 16'h003A; #100;
A = 16'h001F; B = 16'h003B; #100;
A = 16'h001F; B = 16'h003C; #100;
A = 16'h001F; B = 16'h003D; #100;
A = 16'h001F; B = 16'h003E; #100;
A = 16'h001F; B = 16'h003F; #100;
A = 16'h001F; B = 16'h0040; #100;
A = 16'h001F; B = 16'h0041; #100;
A = 16'h001F; B = 16'h0042; #100;
A = 16'h001F; B = 16'h0043; #100;
A = 16'h001F; B = 16'h0044; #100;
A = 16'h001F; B = 16'h0045; #100;
A = 16'h001F; B = 16'h0046; #100;
A = 16'h001F; B = 16'h0047; #100;
A = 16'h001F; B = 16'h0048; #100;
A = 16'h001F; B = 16'h0049; #100;
A = 16'h001F; B = 16'h004A; #100;
A = 16'h001F; B = 16'h004B; #100;
A = 16'h001F; B = 16'h004C; #100;
A = 16'h001F; B = 16'h004D; #100;
A = 16'h001F; B = 16'h004E; #100;
A = 16'h001F; B = 16'h004F; #100;
A = 16'h001F; B = 16'h0050; #100;
A = 16'h001F; B = 16'h0051; #100;
A = 16'h001F; B = 16'h0052; #100;
A = 16'h001F; B = 16'h0053; #100;
A = 16'h001F; B = 16'h0054; #100;
A = 16'h001F; B = 16'h0055; #100;
A = 16'h001F; B = 16'h0056; #100;
A = 16'h001F; B = 16'h0057; #100;
A = 16'h001F; B = 16'h0058; #100;
A = 16'h001F; B = 16'h0059; #100;
A = 16'h001F; B = 16'h005A; #100;
A = 16'h001F; B = 16'h005B; #100;
A = 16'h001F; B = 16'h005C; #100;
A = 16'h001F; B = 16'h005D; #100;
A = 16'h001F; B = 16'h005E; #100;
A = 16'h001F; B = 16'h005F; #100;
A = 16'h001F; B = 16'h0060; #100;
A = 16'h001F; B = 16'h0061; #100;
A = 16'h001F; B = 16'h0062; #100;
A = 16'h001F; B = 16'h0063; #100;
A = 16'h001F; B = 16'h0064; #100;
A = 16'h001F; B = 16'h0065; #100;
A = 16'h001F; B = 16'h0066; #100;
A = 16'h001F; B = 16'h0067; #100;
A = 16'h001F; B = 16'h0068; #100;
A = 16'h001F; B = 16'h0069; #100;
A = 16'h001F; B = 16'h006A; #100;
A = 16'h001F; B = 16'h006B; #100;
A = 16'h001F; B = 16'h006C; #100;
A = 16'h001F; B = 16'h006D; #100;
A = 16'h001F; B = 16'h006E; #100;
A = 16'h001F; B = 16'h006F; #100;
A = 16'h001F; B = 16'h0070; #100;
A = 16'h001F; B = 16'h0071; #100;
A = 16'h001F; B = 16'h0072; #100;
A = 16'h001F; B = 16'h0073; #100;
A = 16'h001F; B = 16'h0074; #100;
A = 16'h001F; B = 16'h0075; #100;
A = 16'h001F; B = 16'h0076; #100;
A = 16'h001F; B = 16'h0077; #100;
A = 16'h001F; B = 16'h0078; #100;
A = 16'h001F; B = 16'h0079; #100;
A = 16'h001F; B = 16'h007A; #100;
A = 16'h001F; B = 16'h007B; #100;
A = 16'h001F; B = 16'h007C; #100;
A = 16'h001F; B = 16'h007D; #100;
A = 16'h001F; B = 16'h007E; #100;
A = 16'h001F; B = 16'h007F; #100;
A = 16'h001F; B = 16'h0080; #100;
A = 16'h001F; B = 16'h0081; #100;
A = 16'h001F; B = 16'h0082; #100;
A = 16'h001F; B = 16'h0083; #100;
A = 16'h001F; B = 16'h0084; #100;
A = 16'h001F; B = 16'h0085; #100;
A = 16'h001F; B = 16'h0086; #100;
A = 16'h001F; B = 16'h0087; #100;
A = 16'h001F; B = 16'h0088; #100;
A = 16'h001F; B = 16'h0089; #100;
A = 16'h001F; B = 16'h008A; #100;
A = 16'h001F; B = 16'h008B; #100;
A = 16'h001F; B = 16'h008C; #100;
A = 16'h001F; B = 16'h008D; #100;
A = 16'h001F; B = 16'h008E; #100;
A = 16'h001F; B = 16'h008F; #100;
A = 16'h001F; B = 16'h0090; #100;
A = 16'h001F; B = 16'h0091; #100;
A = 16'h001F; B = 16'h0092; #100;
A = 16'h001F; B = 16'h0093; #100;
A = 16'h001F; B = 16'h0094; #100;
A = 16'h001F; B = 16'h0095; #100;
A = 16'h001F; B = 16'h0096; #100;
A = 16'h001F; B = 16'h0097; #100;
A = 16'h001F; B = 16'h0098; #100;
A = 16'h001F; B = 16'h0099; #100;
A = 16'h001F; B = 16'h009A; #100;
A = 16'h001F; B = 16'h009B; #100;
A = 16'h001F; B = 16'h009C; #100;
A = 16'h001F; B = 16'h009D; #100;
A = 16'h001F; B = 16'h009E; #100;
A = 16'h001F; B = 16'h009F; #100;
A = 16'h001F; B = 16'h00A0; #100;
A = 16'h001F; B = 16'h00A1; #100;
A = 16'h001F; B = 16'h00A2; #100;
A = 16'h001F; B = 16'h00A3; #100;
A = 16'h001F; B = 16'h00A4; #100;
A = 16'h001F; B = 16'h00A5; #100;
A = 16'h001F; B = 16'h00A6; #100;
A = 16'h001F; B = 16'h00A7; #100;
A = 16'h001F; B = 16'h00A8; #100;
A = 16'h001F; B = 16'h00A9; #100;
A = 16'h001F; B = 16'h00AA; #100;
A = 16'h001F; B = 16'h00AB; #100;
A = 16'h001F; B = 16'h00AC; #100;
A = 16'h001F; B = 16'h00AD; #100;
A = 16'h001F; B = 16'h00AE; #100;
A = 16'h001F; B = 16'h00AF; #100;
A = 16'h001F; B = 16'h00B0; #100;
A = 16'h001F; B = 16'h00B1; #100;
A = 16'h001F; B = 16'h00B2; #100;
A = 16'h001F; B = 16'h00B3; #100;
A = 16'h001F; B = 16'h00B4; #100;
A = 16'h001F; B = 16'h00B5; #100;
A = 16'h001F; B = 16'h00B6; #100;
A = 16'h001F; B = 16'h00B7; #100;
A = 16'h001F; B = 16'h00B8; #100;
A = 16'h001F; B = 16'h00B9; #100;
A = 16'h001F; B = 16'h00BA; #100;
A = 16'h001F; B = 16'h00BB; #100;
A = 16'h001F; B = 16'h00BC; #100;
A = 16'h001F; B = 16'h00BD; #100;
A = 16'h001F; B = 16'h00BE; #100;
A = 16'h001F; B = 16'h00BF; #100;
A = 16'h001F; B = 16'h00C0; #100;
A = 16'h001F; B = 16'h00C1; #100;
A = 16'h001F; B = 16'h00C2; #100;
A = 16'h001F; B = 16'h00C3; #100;
A = 16'h001F; B = 16'h00C4; #100;
A = 16'h001F; B = 16'h00C5; #100;
A = 16'h001F; B = 16'h00C6; #100;
A = 16'h001F; B = 16'h00C7; #100;
A = 16'h001F; B = 16'h00C8; #100;
A = 16'h001F; B = 16'h00C9; #100;
A = 16'h001F; B = 16'h00CA; #100;
A = 16'h001F; B = 16'h00CB; #100;
A = 16'h001F; B = 16'h00CC; #100;
A = 16'h001F; B = 16'h00CD; #100;
A = 16'h001F; B = 16'h00CE; #100;
A = 16'h001F; B = 16'h00CF; #100;
A = 16'h001F; B = 16'h00D0; #100;
A = 16'h001F; B = 16'h00D1; #100;
A = 16'h001F; B = 16'h00D2; #100;
A = 16'h001F; B = 16'h00D3; #100;
A = 16'h001F; B = 16'h00D4; #100;
A = 16'h001F; B = 16'h00D5; #100;
A = 16'h001F; B = 16'h00D6; #100;
A = 16'h001F; B = 16'h00D7; #100;
A = 16'h001F; B = 16'h00D8; #100;
A = 16'h001F; B = 16'h00D9; #100;
A = 16'h001F; B = 16'h00DA; #100;
A = 16'h001F; B = 16'h00DB; #100;
A = 16'h001F; B = 16'h00DC; #100;
A = 16'h001F; B = 16'h00DD; #100;
A = 16'h001F; B = 16'h00DE; #100;
A = 16'h001F; B = 16'h00DF; #100;
A = 16'h001F; B = 16'h00E0; #100;
A = 16'h001F; B = 16'h00E1; #100;
A = 16'h001F; B = 16'h00E2; #100;
A = 16'h001F; B = 16'h00E3; #100;
A = 16'h001F; B = 16'h00E4; #100;
A = 16'h001F; B = 16'h00E5; #100;
A = 16'h001F; B = 16'h00E6; #100;
A = 16'h001F; B = 16'h00E7; #100;
A = 16'h001F; B = 16'h00E8; #100;
A = 16'h001F; B = 16'h00E9; #100;
A = 16'h001F; B = 16'h00EA; #100;
A = 16'h001F; B = 16'h00EB; #100;
A = 16'h001F; B = 16'h00EC; #100;
A = 16'h001F; B = 16'h00ED; #100;
A = 16'h001F; B = 16'h00EE; #100;
A = 16'h001F; B = 16'h00EF; #100;
A = 16'h001F; B = 16'h00F0; #100;
A = 16'h001F; B = 16'h00F1; #100;
A = 16'h001F; B = 16'h00F2; #100;
A = 16'h001F; B = 16'h00F3; #100;
A = 16'h001F; B = 16'h00F4; #100;
A = 16'h001F; B = 16'h00F5; #100;
A = 16'h001F; B = 16'h00F6; #100;
A = 16'h001F; B = 16'h00F7; #100;
A = 16'h001F; B = 16'h00F8; #100;
A = 16'h001F; B = 16'h00F9; #100;
A = 16'h001F; B = 16'h00FA; #100;
A = 16'h001F; B = 16'h00FB; #100;
A = 16'h001F; B = 16'h00FC; #100;
A = 16'h001F; B = 16'h00FD; #100;
A = 16'h001F; B = 16'h00FE; #100;
A = 16'h001F; B = 16'h00FF; #100;
A = 16'h0020; B = 16'h000; #100;
A = 16'h0020; B = 16'h001; #100;
A = 16'h0020; B = 16'h002; #100;
A = 16'h0020; B = 16'h003; #100;
A = 16'h0020; B = 16'h004; #100;
A = 16'h0020; B = 16'h005; #100;
A = 16'h0020; B = 16'h006; #100;
A = 16'h0020; B = 16'h007; #100;
A = 16'h0020; B = 16'h008; #100;
A = 16'h0020; B = 16'h009; #100;
A = 16'h0020; B = 16'h00A; #100;
A = 16'h0020; B = 16'h00B; #100;
A = 16'h0020; B = 16'h00C; #100;
A = 16'h0020; B = 16'h00D; #100;
A = 16'h0020; B = 16'h00E; #100;
A = 16'h0020; B = 16'h00F; #100;
A = 16'h0020; B = 16'h0010; #100;
A = 16'h0020; B = 16'h0011; #100;
A = 16'h0020; B = 16'h0012; #100;
A = 16'h0020; B = 16'h0013; #100;
A = 16'h0020; B = 16'h0014; #100;
A = 16'h0020; B = 16'h0015; #100;
A = 16'h0020; B = 16'h0016; #100;
A = 16'h0020; B = 16'h0017; #100;
A = 16'h0020; B = 16'h0018; #100;
A = 16'h0020; B = 16'h0019; #100;
A = 16'h0020; B = 16'h001A; #100;
A = 16'h0020; B = 16'h001B; #100;
A = 16'h0020; B = 16'h001C; #100;
A = 16'h0020; B = 16'h001D; #100;
A = 16'h0020; B = 16'h001E; #100;
A = 16'h0020; B = 16'h001F; #100;
A = 16'h0020; B = 16'h0020; #100;
A = 16'h0020; B = 16'h0021; #100;
A = 16'h0020; B = 16'h0022; #100;
A = 16'h0020; B = 16'h0023; #100;
A = 16'h0020; B = 16'h0024; #100;
A = 16'h0020; B = 16'h0025; #100;
A = 16'h0020; B = 16'h0026; #100;
A = 16'h0020; B = 16'h0027; #100;
A = 16'h0020; B = 16'h0028; #100;
A = 16'h0020; B = 16'h0029; #100;
A = 16'h0020; B = 16'h002A; #100;
A = 16'h0020; B = 16'h002B; #100;
A = 16'h0020; B = 16'h002C; #100;
A = 16'h0020; B = 16'h002D; #100;
A = 16'h0020; B = 16'h002E; #100;
A = 16'h0020; B = 16'h002F; #100;
A = 16'h0020; B = 16'h0030; #100;
A = 16'h0020; B = 16'h0031; #100;
A = 16'h0020; B = 16'h0032; #100;
A = 16'h0020; B = 16'h0033; #100;
A = 16'h0020; B = 16'h0034; #100;
A = 16'h0020; B = 16'h0035; #100;
A = 16'h0020; B = 16'h0036; #100;
A = 16'h0020; B = 16'h0037; #100;
A = 16'h0020; B = 16'h0038; #100;
A = 16'h0020; B = 16'h0039; #100;
A = 16'h0020; B = 16'h003A; #100;
A = 16'h0020; B = 16'h003B; #100;
A = 16'h0020; B = 16'h003C; #100;
A = 16'h0020; B = 16'h003D; #100;
A = 16'h0020; B = 16'h003E; #100;
A = 16'h0020; B = 16'h003F; #100;
A = 16'h0020; B = 16'h0040; #100;
A = 16'h0020; B = 16'h0041; #100;
A = 16'h0020; B = 16'h0042; #100;
A = 16'h0020; B = 16'h0043; #100;
A = 16'h0020; B = 16'h0044; #100;
A = 16'h0020; B = 16'h0045; #100;
A = 16'h0020; B = 16'h0046; #100;
A = 16'h0020; B = 16'h0047; #100;
A = 16'h0020; B = 16'h0048; #100;
A = 16'h0020; B = 16'h0049; #100;
A = 16'h0020; B = 16'h004A; #100;
A = 16'h0020; B = 16'h004B; #100;
A = 16'h0020; B = 16'h004C; #100;
A = 16'h0020; B = 16'h004D; #100;
A = 16'h0020; B = 16'h004E; #100;
A = 16'h0020; B = 16'h004F; #100;
A = 16'h0020; B = 16'h0050; #100;
A = 16'h0020; B = 16'h0051; #100;
A = 16'h0020; B = 16'h0052; #100;
A = 16'h0020; B = 16'h0053; #100;
A = 16'h0020; B = 16'h0054; #100;
A = 16'h0020; B = 16'h0055; #100;
A = 16'h0020; B = 16'h0056; #100;
A = 16'h0020; B = 16'h0057; #100;
A = 16'h0020; B = 16'h0058; #100;
A = 16'h0020; B = 16'h0059; #100;
A = 16'h0020; B = 16'h005A; #100;
A = 16'h0020; B = 16'h005B; #100;
A = 16'h0020; B = 16'h005C; #100;
A = 16'h0020; B = 16'h005D; #100;
A = 16'h0020; B = 16'h005E; #100;
A = 16'h0020; B = 16'h005F; #100;
A = 16'h0020; B = 16'h0060; #100;
A = 16'h0020; B = 16'h0061; #100;
A = 16'h0020; B = 16'h0062; #100;
A = 16'h0020; B = 16'h0063; #100;
A = 16'h0020; B = 16'h0064; #100;
A = 16'h0020; B = 16'h0065; #100;
A = 16'h0020; B = 16'h0066; #100;
A = 16'h0020; B = 16'h0067; #100;
A = 16'h0020; B = 16'h0068; #100;
A = 16'h0020; B = 16'h0069; #100;
A = 16'h0020; B = 16'h006A; #100;
A = 16'h0020; B = 16'h006B; #100;
A = 16'h0020; B = 16'h006C; #100;
A = 16'h0020; B = 16'h006D; #100;
A = 16'h0020; B = 16'h006E; #100;
A = 16'h0020; B = 16'h006F; #100;
A = 16'h0020; B = 16'h0070; #100;
A = 16'h0020; B = 16'h0071; #100;
A = 16'h0020; B = 16'h0072; #100;
A = 16'h0020; B = 16'h0073; #100;
A = 16'h0020; B = 16'h0074; #100;
A = 16'h0020; B = 16'h0075; #100;
A = 16'h0020; B = 16'h0076; #100;
A = 16'h0020; B = 16'h0077; #100;
A = 16'h0020; B = 16'h0078; #100;
A = 16'h0020; B = 16'h0079; #100;
A = 16'h0020; B = 16'h007A; #100;
A = 16'h0020; B = 16'h007B; #100;
A = 16'h0020; B = 16'h007C; #100;
A = 16'h0020; B = 16'h007D; #100;
A = 16'h0020; B = 16'h007E; #100;
A = 16'h0020; B = 16'h007F; #100;
A = 16'h0020; B = 16'h0080; #100;
A = 16'h0020; B = 16'h0081; #100;
A = 16'h0020; B = 16'h0082; #100;
A = 16'h0020; B = 16'h0083; #100;
A = 16'h0020; B = 16'h0084; #100;
A = 16'h0020; B = 16'h0085; #100;
A = 16'h0020; B = 16'h0086; #100;
A = 16'h0020; B = 16'h0087; #100;
A = 16'h0020; B = 16'h0088; #100;
A = 16'h0020; B = 16'h0089; #100;
A = 16'h0020; B = 16'h008A; #100;
A = 16'h0020; B = 16'h008B; #100;
A = 16'h0020; B = 16'h008C; #100;
A = 16'h0020; B = 16'h008D; #100;
A = 16'h0020; B = 16'h008E; #100;
A = 16'h0020; B = 16'h008F; #100;
A = 16'h0020; B = 16'h0090; #100;
A = 16'h0020; B = 16'h0091; #100;
A = 16'h0020; B = 16'h0092; #100;
A = 16'h0020; B = 16'h0093; #100;
A = 16'h0020; B = 16'h0094; #100;
A = 16'h0020; B = 16'h0095; #100;
A = 16'h0020; B = 16'h0096; #100;
A = 16'h0020; B = 16'h0097; #100;
A = 16'h0020; B = 16'h0098; #100;
A = 16'h0020; B = 16'h0099; #100;
A = 16'h0020; B = 16'h009A; #100;
A = 16'h0020; B = 16'h009B; #100;
A = 16'h0020; B = 16'h009C; #100;
A = 16'h0020; B = 16'h009D; #100;
A = 16'h0020; B = 16'h009E; #100;
A = 16'h0020; B = 16'h009F; #100;
A = 16'h0020; B = 16'h00A0; #100;
A = 16'h0020; B = 16'h00A1; #100;
A = 16'h0020; B = 16'h00A2; #100;
A = 16'h0020; B = 16'h00A3; #100;
A = 16'h0020; B = 16'h00A4; #100;
A = 16'h0020; B = 16'h00A5; #100;
A = 16'h0020; B = 16'h00A6; #100;
A = 16'h0020; B = 16'h00A7; #100;
A = 16'h0020; B = 16'h00A8; #100;
A = 16'h0020; B = 16'h00A9; #100;
A = 16'h0020; B = 16'h00AA; #100;
A = 16'h0020; B = 16'h00AB; #100;
A = 16'h0020; B = 16'h00AC; #100;
A = 16'h0020; B = 16'h00AD; #100;
A = 16'h0020; B = 16'h00AE; #100;
A = 16'h0020; B = 16'h00AF; #100;
A = 16'h0020; B = 16'h00B0; #100;
A = 16'h0020; B = 16'h00B1; #100;
A = 16'h0020; B = 16'h00B2; #100;
A = 16'h0020; B = 16'h00B3; #100;
A = 16'h0020; B = 16'h00B4; #100;
A = 16'h0020; B = 16'h00B5; #100;
A = 16'h0020; B = 16'h00B6; #100;
A = 16'h0020; B = 16'h00B7; #100;
A = 16'h0020; B = 16'h00B8; #100;
A = 16'h0020; B = 16'h00B9; #100;
A = 16'h0020; B = 16'h00BA; #100;
A = 16'h0020; B = 16'h00BB; #100;
A = 16'h0020; B = 16'h00BC; #100;
A = 16'h0020; B = 16'h00BD; #100;
A = 16'h0020; B = 16'h00BE; #100;
A = 16'h0020; B = 16'h00BF; #100;
A = 16'h0020; B = 16'h00C0; #100;
A = 16'h0020; B = 16'h00C1; #100;
A = 16'h0020; B = 16'h00C2; #100;
A = 16'h0020; B = 16'h00C3; #100;
A = 16'h0020; B = 16'h00C4; #100;
A = 16'h0020; B = 16'h00C5; #100;
A = 16'h0020; B = 16'h00C6; #100;
A = 16'h0020; B = 16'h00C7; #100;
A = 16'h0020; B = 16'h00C8; #100;
A = 16'h0020; B = 16'h00C9; #100;
A = 16'h0020; B = 16'h00CA; #100;
A = 16'h0020; B = 16'h00CB; #100;
A = 16'h0020; B = 16'h00CC; #100;
A = 16'h0020; B = 16'h00CD; #100;
A = 16'h0020; B = 16'h00CE; #100;
A = 16'h0020; B = 16'h00CF; #100;
A = 16'h0020; B = 16'h00D0; #100;
A = 16'h0020; B = 16'h00D1; #100;
A = 16'h0020; B = 16'h00D2; #100;
A = 16'h0020; B = 16'h00D3; #100;
A = 16'h0020; B = 16'h00D4; #100;
A = 16'h0020; B = 16'h00D5; #100;
A = 16'h0020; B = 16'h00D6; #100;
A = 16'h0020; B = 16'h00D7; #100;
A = 16'h0020; B = 16'h00D8; #100;
A = 16'h0020; B = 16'h00D9; #100;
A = 16'h0020; B = 16'h00DA; #100;
A = 16'h0020; B = 16'h00DB; #100;
A = 16'h0020; B = 16'h00DC; #100;
A = 16'h0020; B = 16'h00DD; #100;
A = 16'h0020; B = 16'h00DE; #100;
A = 16'h0020; B = 16'h00DF; #100;
A = 16'h0020; B = 16'h00E0; #100;
A = 16'h0020; B = 16'h00E1; #100;
A = 16'h0020; B = 16'h00E2; #100;
A = 16'h0020; B = 16'h00E3; #100;
A = 16'h0020; B = 16'h00E4; #100;
A = 16'h0020; B = 16'h00E5; #100;
A = 16'h0020; B = 16'h00E6; #100;
A = 16'h0020; B = 16'h00E7; #100;
A = 16'h0020; B = 16'h00E8; #100;
A = 16'h0020; B = 16'h00E9; #100;
A = 16'h0020; B = 16'h00EA; #100;
A = 16'h0020; B = 16'h00EB; #100;
A = 16'h0020; B = 16'h00EC; #100;
A = 16'h0020; B = 16'h00ED; #100;
A = 16'h0020; B = 16'h00EE; #100;
A = 16'h0020; B = 16'h00EF; #100;
A = 16'h0020; B = 16'h00F0; #100;
A = 16'h0020; B = 16'h00F1; #100;
A = 16'h0020; B = 16'h00F2; #100;
A = 16'h0020; B = 16'h00F3; #100;
A = 16'h0020; B = 16'h00F4; #100;
A = 16'h0020; B = 16'h00F5; #100;
A = 16'h0020; B = 16'h00F6; #100;
A = 16'h0020; B = 16'h00F7; #100;
A = 16'h0020; B = 16'h00F8; #100;
A = 16'h0020; B = 16'h00F9; #100;
A = 16'h0020; B = 16'h00FA; #100;
A = 16'h0020; B = 16'h00FB; #100;
A = 16'h0020; B = 16'h00FC; #100;
A = 16'h0020; B = 16'h00FD; #100;
A = 16'h0020; B = 16'h00FE; #100;
A = 16'h0020; B = 16'h00FF; #100;
A = 16'h0021; B = 16'h000; #100;
A = 16'h0021; B = 16'h001; #100;
A = 16'h0021; B = 16'h002; #100;
A = 16'h0021; B = 16'h003; #100;
A = 16'h0021; B = 16'h004; #100;
A = 16'h0021; B = 16'h005; #100;
A = 16'h0021; B = 16'h006; #100;
A = 16'h0021; B = 16'h007; #100;
A = 16'h0021; B = 16'h008; #100;
A = 16'h0021; B = 16'h009; #100;
A = 16'h0021; B = 16'h00A; #100;
A = 16'h0021; B = 16'h00B; #100;
A = 16'h0021; B = 16'h00C; #100;
A = 16'h0021; B = 16'h00D; #100;
A = 16'h0021; B = 16'h00E; #100;
A = 16'h0021; B = 16'h00F; #100;
A = 16'h0021; B = 16'h0010; #100;
A = 16'h0021; B = 16'h0011; #100;
A = 16'h0021; B = 16'h0012; #100;
A = 16'h0021; B = 16'h0013; #100;
A = 16'h0021; B = 16'h0014; #100;
A = 16'h0021; B = 16'h0015; #100;
A = 16'h0021; B = 16'h0016; #100;
A = 16'h0021; B = 16'h0017; #100;
A = 16'h0021; B = 16'h0018; #100;
A = 16'h0021; B = 16'h0019; #100;
A = 16'h0021; B = 16'h001A; #100;
A = 16'h0021; B = 16'h001B; #100;
A = 16'h0021; B = 16'h001C; #100;
A = 16'h0021; B = 16'h001D; #100;
A = 16'h0021; B = 16'h001E; #100;
A = 16'h0021; B = 16'h001F; #100;
A = 16'h0021; B = 16'h0020; #100;
A = 16'h0021; B = 16'h0021; #100;
A = 16'h0021; B = 16'h0022; #100;
A = 16'h0021; B = 16'h0023; #100;
A = 16'h0021; B = 16'h0024; #100;
A = 16'h0021; B = 16'h0025; #100;
A = 16'h0021; B = 16'h0026; #100;
A = 16'h0021; B = 16'h0027; #100;
A = 16'h0021; B = 16'h0028; #100;
A = 16'h0021; B = 16'h0029; #100;
A = 16'h0021; B = 16'h002A; #100;
A = 16'h0021; B = 16'h002B; #100;
A = 16'h0021; B = 16'h002C; #100;
A = 16'h0021; B = 16'h002D; #100;
A = 16'h0021; B = 16'h002E; #100;
A = 16'h0021; B = 16'h002F; #100;
A = 16'h0021; B = 16'h0030; #100;
A = 16'h0021; B = 16'h0031; #100;
A = 16'h0021; B = 16'h0032; #100;
A = 16'h0021; B = 16'h0033; #100;
A = 16'h0021; B = 16'h0034; #100;
A = 16'h0021; B = 16'h0035; #100;
A = 16'h0021; B = 16'h0036; #100;
A = 16'h0021; B = 16'h0037; #100;
A = 16'h0021; B = 16'h0038; #100;
A = 16'h0021; B = 16'h0039; #100;
A = 16'h0021; B = 16'h003A; #100;
A = 16'h0021; B = 16'h003B; #100;
A = 16'h0021; B = 16'h003C; #100;
A = 16'h0021; B = 16'h003D; #100;
A = 16'h0021; B = 16'h003E; #100;
A = 16'h0021; B = 16'h003F; #100;
A = 16'h0021; B = 16'h0040; #100;
A = 16'h0021; B = 16'h0041; #100;
A = 16'h0021; B = 16'h0042; #100;
A = 16'h0021; B = 16'h0043; #100;
A = 16'h0021; B = 16'h0044; #100;
A = 16'h0021; B = 16'h0045; #100;
A = 16'h0021; B = 16'h0046; #100;
A = 16'h0021; B = 16'h0047; #100;
A = 16'h0021; B = 16'h0048; #100;
A = 16'h0021; B = 16'h0049; #100;
A = 16'h0021; B = 16'h004A; #100;
A = 16'h0021; B = 16'h004B; #100;
A = 16'h0021; B = 16'h004C; #100;
A = 16'h0021; B = 16'h004D; #100;
A = 16'h0021; B = 16'h004E; #100;
A = 16'h0021; B = 16'h004F; #100;
A = 16'h0021; B = 16'h0050; #100;
A = 16'h0021; B = 16'h0051; #100;
A = 16'h0021; B = 16'h0052; #100;
A = 16'h0021; B = 16'h0053; #100;
A = 16'h0021; B = 16'h0054; #100;
A = 16'h0021; B = 16'h0055; #100;
A = 16'h0021; B = 16'h0056; #100;
A = 16'h0021; B = 16'h0057; #100;
A = 16'h0021; B = 16'h0058; #100;
A = 16'h0021; B = 16'h0059; #100;
A = 16'h0021; B = 16'h005A; #100;
A = 16'h0021; B = 16'h005B; #100;
A = 16'h0021; B = 16'h005C; #100;
A = 16'h0021; B = 16'h005D; #100;
A = 16'h0021; B = 16'h005E; #100;
A = 16'h0021; B = 16'h005F; #100;
A = 16'h0021; B = 16'h0060; #100;
A = 16'h0021; B = 16'h0061; #100;
A = 16'h0021; B = 16'h0062; #100;
A = 16'h0021; B = 16'h0063; #100;
A = 16'h0021; B = 16'h0064; #100;
A = 16'h0021; B = 16'h0065; #100;
A = 16'h0021; B = 16'h0066; #100;
A = 16'h0021; B = 16'h0067; #100;
A = 16'h0021; B = 16'h0068; #100;
A = 16'h0021; B = 16'h0069; #100;
A = 16'h0021; B = 16'h006A; #100;
A = 16'h0021; B = 16'h006B; #100;
A = 16'h0021; B = 16'h006C; #100;
A = 16'h0021; B = 16'h006D; #100;
A = 16'h0021; B = 16'h006E; #100;
A = 16'h0021; B = 16'h006F; #100;
A = 16'h0021; B = 16'h0070; #100;
A = 16'h0021; B = 16'h0071; #100;
A = 16'h0021; B = 16'h0072; #100;
A = 16'h0021; B = 16'h0073; #100;
A = 16'h0021; B = 16'h0074; #100;
A = 16'h0021; B = 16'h0075; #100;
A = 16'h0021; B = 16'h0076; #100;
A = 16'h0021; B = 16'h0077; #100;
A = 16'h0021; B = 16'h0078; #100;
A = 16'h0021; B = 16'h0079; #100;
A = 16'h0021; B = 16'h007A; #100;
A = 16'h0021; B = 16'h007B; #100;
A = 16'h0021; B = 16'h007C; #100;
A = 16'h0021; B = 16'h007D; #100;
A = 16'h0021; B = 16'h007E; #100;
A = 16'h0021; B = 16'h007F; #100;
A = 16'h0021; B = 16'h0080; #100;
A = 16'h0021; B = 16'h0081; #100;
A = 16'h0021; B = 16'h0082; #100;
A = 16'h0021; B = 16'h0083; #100;
A = 16'h0021; B = 16'h0084; #100;
A = 16'h0021; B = 16'h0085; #100;
A = 16'h0021; B = 16'h0086; #100;
A = 16'h0021; B = 16'h0087; #100;
A = 16'h0021; B = 16'h0088; #100;
A = 16'h0021; B = 16'h0089; #100;
A = 16'h0021; B = 16'h008A; #100;
A = 16'h0021; B = 16'h008B; #100;
A = 16'h0021; B = 16'h008C; #100;
A = 16'h0021; B = 16'h008D; #100;
A = 16'h0021; B = 16'h008E; #100;
A = 16'h0021; B = 16'h008F; #100;
A = 16'h0021; B = 16'h0090; #100;
A = 16'h0021; B = 16'h0091; #100;
A = 16'h0021; B = 16'h0092; #100;
A = 16'h0021; B = 16'h0093; #100;
A = 16'h0021; B = 16'h0094; #100;
A = 16'h0021; B = 16'h0095; #100;
A = 16'h0021; B = 16'h0096; #100;
A = 16'h0021; B = 16'h0097; #100;
A = 16'h0021; B = 16'h0098; #100;
A = 16'h0021; B = 16'h0099; #100;
A = 16'h0021; B = 16'h009A; #100;
A = 16'h0021; B = 16'h009B; #100;
A = 16'h0021; B = 16'h009C; #100;
A = 16'h0021; B = 16'h009D; #100;
A = 16'h0021; B = 16'h009E; #100;
A = 16'h0021; B = 16'h009F; #100;
A = 16'h0021; B = 16'h00A0; #100;
A = 16'h0021; B = 16'h00A1; #100;
A = 16'h0021; B = 16'h00A2; #100;
A = 16'h0021; B = 16'h00A3; #100;
A = 16'h0021; B = 16'h00A4; #100;
A = 16'h0021; B = 16'h00A5; #100;
A = 16'h0021; B = 16'h00A6; #100;
A = 16'h0021; B = 16'h00A7; #100;
A = 16'h0021; B = 16'h00A8; #100;
A = 16'h0021; B = 16'h00A9; #100;
A = 16'h0021; B = 16'h00AA; #100;
A = 16'h0021; B = 16'h00AB; #100;
A = 16'h0021; B = 16'h00AC; #100;
A = 16'h0021; B = 16'h00AD; #100;
A = 16'h0021; B = 16'h00AE; #100;
A = 16'h0021; B = 16'h00AF; #100;
A = 16'h0021; B = 16'h00B0; #100;
A = 16'h0021; B = 16'h00B1; #100;
A = 16'h0021; B = 16'h00B2; #100;
A = 16'h0021; B = 16'h00B3; #100;
A = 16'h0021; B = 16'h00B4; #100;
A = 16'h0021; B = 16'h00B5; #100;
A = 16'h0021; B = 16'h00B6; #100;
A = 16'h0021; B = 16'h00B7; #100;
A = 16'h0021; B = 16'h00B8; #100;
A = 16'h0021; B = 16'h00B9; #100;
A = 16'h0021; B = 16'h00BA; #100;
A = 16'h0021; B = 16'h00BB; #100;
A = 16'h0021; B = 16'h00BC; #100;
A = 16'h0021; B = 16'h00BD; #100;
A = 16'h0021; B = 16'h00BE; #100;
A = 16'h0021; B = 16'h00BF; #100;
A = 16'h0021; B = 16'h00C0; #100;
A = 16'h0021; B = 16'h00C1; #100;
A = 16'h0021; B = 16'h00C2; #100;
A = 16'h0021; B = 16'h00C3; #100;
A = 16'h0021; B = 16'h00C4; #100;
A = 16'h0021; B = 16'h00C5; #100;
A = 16'h0021; B = 16'h00C6; #100;
A = 16'h0021; B = 16'h00C7; #100;
A = 16'h0021; B = 16'h00C8; #100;
A = 16'h0021; B = 16'h00C9; #100;
A = 16'h0021; B = 16'h00CA; #100;
A = 16'h0021; B = 16'h00CB; #100;
A = 16'h0021; B = 16'h00CC; #100;
A = 16'h0021; B = 16'h00CD; #100;
A = 16'h0021; B = 16'h00CE; #100;
A = 16'h0021; B = 16'h00CF; #100;
A = 16'h0021; B = 16'h00D0; #100;
A = 16'h0021; B = 16'h00D1; #100;
A = 16'h0021; B = 16'h00D2; #100;
A = 16'h0021; B = 16'h00D3; #100;
A = 16'h0021; B = 16'h00D4; #100;
A = 16'h0021; B = 16'h00D5; #100;
A = 16'h0021; B = 16'h00D6; #100;
A = 16'h0021; B = 16'h00D7; #100;
A = 16'h0021; B = 16'h00D8; #100;
A = 16'h0021; B = 16'h00D9; #100;
A = 16'h0021; B = 16'h00DA; #100;
A = 16'h0021; B = 16'h00DB; #100;
A = 16'h0021; B = 16'h00DC; #100;
A = 16'h0021; B = 16'h00DD; #100;
A = 16'h0021; B = 16'h00DE; #100;
A = 16'h0021; B = 16'h00DF; #100;
A = 16'h0021; B = 16'h00E0; #100;
A = 16'h0021; B = 16'h00E1; #100;
A = 16'h0021; B = 16'h00E2; #100;
A = 16'h0021; B = 16'h00E3; #100;
A = 16'h0021; B = 16'h00E4; #100;
A = 16'h0021; B = 16'h00E5; #100;
A = 16'h0021; B = 16'h00E6; #100;
A = 16'h0021; B = 16'h00E7; #100;
A = 16'h0021; B = 16'h00E8; #100;
A = 16'h0021; B = 16'h00E9; #100;
A = 16'h0021; B = 16'h00EA; #100;
A = 16'h0021; B = 16'h00EB; #100;
A = 16'h0021; B = 16'h00EC; #100;
A = 16'h0021; B = 16'h00ED; #100;
A = 16'h0021; B = 16'h00EE; #100;
A = 16'h0021; B = 16'h00EF; #100;
A = 16'h0021; B = 16'h00F0; #100;
A = 16'h0021; B = 16'h00F1; #100;
A = 16'h0021; B = 16'h00F2; #100;
A = 16'h0021; B = 16'h00F3; #100;
A = 16'h0021; B = 16'h00F4; #100;
A = 16'h0021; B = 16'h00F5; #100;
A = 16'h0021; B = 16'h00F6; #100;
A = 16'h0021; B = 16'h00F7; #100;
A = 16'h0021; B = 16'h00F8; #100;
A = 16'h0021; B = 16'h00F9; #100;
A = 16'h0021; B = 16'h00FA; #100;
A = 16'h0021; B = 16'h00FB; #100;
A = 16'h0021; B = 16'h00FC; #100;
A = 16'h0021; B = 16'h00FD; #100;
A = 16'h0021; B = 16'h00FE; #100;
A = 16'h0021; B = 16'h00FF; #100;
A = 16'h0022; B = 16'h000; #100;
A = 16'h0022; B = 16'h001; #100;
A = 16'h0022; B = 16'h002; #100;
A = 16'h0022; B = 16'h003; #100;
A = 16'h0022; B = 16'h004; #100;
A = 16'h0022; B = 16'h005; #100;
A = 16'h0022; B = 16'h006; #100;
A = 16'h0022; B = 16'h007; #100;
A = 16'h0022; B = 16'h008; #100;
A = 16'h0022; B = 16'h009; #100;
A = 16'h0022; B = 16'h00A; #100;
A = 16'h0022; B = 16'h00B; #100;
A = 16'h0022; B = 16'h00C; #100;
A = 16'h0022; B = 16'h00D; #100;
A = 16'h0022; B = 16'h00E; #100;
A = 16'h0022; B = 16'h00F; #100;
A = 16'h0022; B = 16'h0010; #100;
A = 16'h0022; B = 16'h0011; #100;
A = 16'h0022; B = 16'h0012; #100;
A = 16'h0022; B = 16'h0013; #100;
A = 16'h0022; B = 16'h0014; #100;
A = 16'h0022; B = 16'h0015; #100;
A = 16'h0022; B = 16'h0016; #100;
A = 16'h0022; B = 16'h0017; #100;
A = 16'h0022; B = 16'h0018; #100;
A = 16'h0022; B = 16'h0019; #100;
A = 16'h0022; B = 16'h001A; #100;
A = 16'h0022; B = 16'h001B; #100;
A = 16'h0022; B = 16'h001C; #100;
A = 16'h0022; B = 16'h001D; #100;
A = 16'h0022; B = 16'h001E; #100;
A = 16'h0022; B = 16'h001F; #100;
A = 16'h0022; B = 16'h0020; #100;
A = 16'h0022; B = 16'h0021; #100;
A = 16'h0022; B = 16'h0022; #100;
A = 16'h0022; B = 16'h0023; #100;
A = 16'h0022; B = 16'h0024; #100;
A = 16'h0022; B = 16'h0025; #100;
A = 16'h0022; B = 16'h0026; #100;
A = 16'h0022; B = 16'h0027; #100;
A = 16'h0022; B = 16'h0028; #100;
A = 16'h0022; B = 16'h0029; #100;
A = 16'h0022; B = 16'h002A; #100;
A = 16'h0022; B = 16'h002B; #100;
A = 16'h0022; B = 16'h002C; #100;
A = 16'h0022; B = 16'h002D; #100;
A = 16'h0022; B = 16'h002E; #100;
A = 16'h0022; B = 16'h002F; #100;
A = 16'h0022; B = 16'h0030; #100;
A = 16'h0022; B = 16'h0031; #100;
A = 16'h0022; B = 16'h0032; #100;
A = 16'h0022; B = 16'h0033; #100;
A = 16'h0022; B = 16'h0034; #100;
A = 16'h0022; B = 16'h0035; #100;
A = 16'h0022; B = 16'h0036; #100;
A = 16'h0022; B = 16'h0037; #100;
A = 16'h0022; B = 16'h0038; #100;
A = 16'h0022; B = 16'h0039; #100;
A = 16'h0022; B = 16'h003A; #100;
A = 16'h0022; B = 16'h003B; #100;
A = 16'h0022; B = 16'h003C; #100;
A = 16'h0022; B = 16'h003D; #100;
A = 16'h0022; B = 16'h003E; #100;
A = 16'h0022; B = 16'h003F; #100;
A = 16'h0022; B = 16'h0040; #100;
A = 16'h0022; B = 16'h0041; #100;
A = 16'h0022; B = 16'h0042; #100;
A = 16'h0022; B = 16'h0043; #100;
A = 16'h0022; B = 16'h0044; #100;
A = 16'h0022; B = 16'h0045; #100;
A = 16'h0022; B = 16'h0046; #100;
A = 16'h0022; B = 16'h0047; #100;
A = 16'h0022; B = 16'h0048; #100;
A = 16'h0022; B = 16'h0049; #100;
A = 16'h0022; B = 16'h004A; #100;
A = 16'h0022; B = 16'h004B; #100;
A = 16'h0022; B = 16'h004C; #100;
A = 16'h0022; B = 16'h004D; #100;
A = 16'h0022; B = 16'h004E; #100;
A = 16'h0022; B = 16'h004F; #100;
A = 16'h0022; B = 16'h0050; #100;
A = 16'h0022; B = 16'h0051; #100;
A = 16'h0022; B = 16'h0052; #100;
A = 16'h0022; B = 16'h0053; #100;
A = 16'h0022; B = 16'h0054; #100;
A = 16'h0022; B = 16'h0055; #100;
A = 16'h0022; B = 16'h0056; #100;
A = 16'h0022; B = 16'h0057; #100;
A = 16'h0022; B = 16'h0058; #100;
A = 16'h0022; B = 16'h0059; #100;
A = 16'h0022; B = 16'h005A; #100;
A = 16'h0022; B = 16'h005B; #100;
A = 16'h0022; B = 16'h005C; #100;
A = 16'h0022; B = 16'h005D; #100;
A = 16'h0022; B = 16'h005E; #100;
A = 16'h0022; B = 16'h005F; #100;
A = 16'h0022; B = 16'h0060; #100;
A = 16'h0022; B = 16'h0061; #100;
A = 16'h0022; B = 16'h0062; #100;
A = 16'h0022; B = 16'h0063; #100;
A = 16'h0022; B = 16'h0064; #100;
A = 16'h0022; B = 16'h0065; #100;
A = 16'h0022; B = 16'h0066; #100;
A = 16'h0022; B = 16'h0067; #100;
A = 16'h0022; B = 16'h0068; #100;
A = 16'h0022; B = 16'h0069; #100;
A = 16'h0022; B = 16'h006A; #100;
A = 16'h0022; B = 16'h006B; #100;
A = 16'h0022; B = 16'h006C; #100;
A = 16'h0022; B = 16'h006D; #100;
A = 16'h0022; B = 16'h006E; #100;
A = 16'h0022; B = 16'h006F; #100;
A = 16'h0022; B = 16'h0070; #100;
A = 16'h0022; B = 16'h0071; #100;
A = 16'h0022; B = 16'h0072; #100;
A = 16'h0022; B = 16'h0073; #100;
A = 16'h0022; B = 16'h0074; #100;
A = 16'h0022; B = 16'h0075; #100;
A = 16'h0022; B = 16'h0076; #100;
A = 16'h0022; B = 16'h0077; #100;
A = 16'h0022; B = 16'h0078; #100;
A = 16'h0022; B = 16'h0079; #100;
A = 16'h0022; B = 16'h007A; #100;
A = 16'h0022; B = 16'h007B; #100;
A = 16'h0022; B = 16'h007C; #100;
A = 16'h0022; B = 16'h007D; #100;
A = 16'h0022; B = 16'h007E; #100;
A = 16'h0022; B = 16'h007F; #100;
A = 16'h0022; B = 16'h0080; #100;
A = 16'h0022; B = 16'h0081; #100;
A = 16'h0022; B = 16'h0082; #100;
A = 16'h0022; B = 16'h0083; #100;
A = 16'h0022; B = 16'h0084; #100;
A = 16'h0022; B = 16'h0085; #100;
A = 16'h0022; B = 16'h0086; #100;
A = 16'h0022; B = 16'h0087; #100;
A = 16'h0022; B = 16'h0088; #100;
A = 16'h0022; B = 16'h0089; #100;
A = 16'h0022; B = 16'h008A; #100;
A = 16'h0022; B = 16'h008B; #100;
A = 16'h0022; B = 16'h008C; #100;
A = 16'h0022; B = 16'h008D; #100;
A = 16'h0022; B = 16'h008E; #100;
A = 16'h0022; B = 16'h008F; #100;
A = 16'h0022; B = 16'h0090; #100;
A = 16'h0022; B = 16'h0091; #100;
A = 16'h0022; B = 16'h0092; #100;
A = 16'h0022; B = 16'h0093; #100;
A = 16'h0022; B = 16'h0094; #100;
A = 16'h0022; B = 16'h0095; #100;
A = 16'h0022; B = 16'h0096; #100;
A = 16'h0022; B = 16'h0097; #100;
A = 16'h0022; B = 16'h0098; #100;
A = 16'h0022; B = 16'h0099; #100;
A = 16'h0022; B = 16'h009A; #100;
A = 16'h0022; B = 16'h009B; #100;
A = 16'h0022; B = 16'h009C; #100;
A = 16'h0022; B = 16'h009D; #100;
A = 16'h0022; B = 16'h009E; #100;
A = 16'h0022; B = 16'h009F; #100;
A = 16'h0022; B = 16'h00A0; #100;
A = 16'h0022; B = 16'h00A1; #100;
A = 16'h0022; B = 16'h00A2; #100;
A = 16'h0022; B = 16'h00A3; #100;
A = 16'h0022; B = 16'h00A4; #100;
A = 16'h0022; B = 16'h00A5; #100;
A = 16'h0022; B = 16'h00A6; #100;
A = 16'h0022; B = 16'h00A7; #100;
A = 16'h0022; B = 16'h00A8; #100;
A = 16'h0022; B = 16'h00A9; #100;
A = 16'h0022; B = 16'h00AA; #100;
A = 16'h0022; B = 16'h00AB; #100;
A = 16'h0022; B = 16'h00AC; #100;
A = 16'h0022; B = 16'h00AD; #100;
A = 16'h0022; B = 16'h00AE; #100;
A = 16'h0022; B = 16'h00AF; #100;
A = 16'h0022; B = 16'h00B0; #100;
A = 16'h0022; B = 16'h00B1; #100;
A = 16'h0022; B = 16'h00B2; #100;
A = 16'h0022; B = 16'h00B3; #100;
A = 16'h0022; B = 16'h00B4; #100;
A = 16'h0022; B = 16'h00B5; #100;
A = 16'h0022; B = 16'h00B6; #100;
A = 16'h0022; B = 16'h00B7; #100;
A = 16'h0022; B = 16'h00B8; #100;
A = 16'h0022; B = 16'h00B9; #100;
A = 16'h0022; B = 16'h00BA; #100;
A = 16'h0022; B = 16'h00BB; #100;
A = 16'h0022; B = 16'h00BC; #100;
A = 16'h0022; B = 16'h00BD; #100;
A = 16'h0022; B = 16'h00BE; #100;
A = 16'h0022; B = 16'h00BF; #100;
A = 16'h0022; B = 16'h00C0; #100;
A = 16'h0022; B = 16'h00C1; #100;
A = 16'h0022; B = 16'h00C2; #100;
A = 16'h0022; B = 16'h00C3; #100;
A = 16'h0022; B = 16'h00C4; #100;
A = 16'h0022; B = 16'h00C5; #100;
A = 16'h0022; B = 16'h00C6; #100;
A = 16'h0022; B = 16'h00C7; #100;
A = 16'h0022; B = 16'h00C8; #100;
A = 16'h0022; B = 16'h00C9; #100;
A = 16'h0022; B = 16'h00CA; #100;
A = 16'h0022; B = 16'h00CB; #100;
A = 16'h0022; B = 16'h00CC; #100;
A = 16'h0022; B = 16'h00CD; #100;
A = 16'h0022; B = 16'h00CE; #100;
A = 16'h0022; B = 16'h00CF; #100;
A = 16'h0022; B = 16'h00D0; #100;
A = 16'h0022; B = 16'h00D1; #100;
A = 16'h0022; B = 16'h00D2; #100;
A = 16'h0022; B = 16'h00D3; #100;
A = 16'h0022; B = 16'h00D4; #100;
A = 16'h0022; B = 16'h00D5; #100;
A = 16'h0022; B = 16'h00D6; #100;
A = 16'h0022; B = 16'h00D7; #100;
A = 16'h0022; B = 16'h00D8; #100;
A = 16'h0022; B = 16'h00D9; #100;
A = 16'h0022; B = 16'h00DA; #100;
A = 16'h0022; B = 16'h00DB; #100;
A = 16'h0022; B = 16'h00DC; #100;
A = 16'h0022; B = 16'h00DD; #100;
A = 16'h0022; B = 16'h00DE; #100;
A = 16'h0022; B = 16'h00DF; #100;
A = 16'h0022; B = 16'h00E0; #100;
A = 16'h0022; B = 16'h00E1; #100;
A = 16'h0022; B = 16'h00E2; #100;
A = 16'h0022; B = 16'h00E3; #100;
A = 16'h0022; B = 16'h00E4; #100;
A = 16'h0022; B = 16'h00E5; #100;
A = 16'h0022; B = 16'h00E6; #100;
A = 16'h0022; B = 16'h00E7; #100;
A = 16'h0022; B = 16'h00E8; #100;
A = 16'h0022; B = 16'h00E9; #100;
A = 16'h0022; B = 16'h00EA; #100;
A = 16'h0022; B = 16'h00EB; #100;
A = 16'h0022; B = 16'h00EC; #100;
A = 16'h0022; B = 16'h00ED; #100;
A = 16'h0022; B = 16'h00EE; #100;
A = 16'h0022; B = 16'h00EF; #100;
A = 16'h0022; B = 16'h00F0; #100;
A = 16'h0022; B = 16'h00F1; #100;
A = 16'h0022; B = 16'h00F2; #100;
A = 16'h0022; B = 16'h00F3; #100;
A = 16'h0022; B = 16'h00F4; #100;
A = 16'h0022; B = 16'h00F5; #100;
A = 16'h0022; B = 16'h00F6; #100;
A = 16'h0022; B = 16'h00F7; #100;
A = 16'h0022; B = 16'h00F8; #100;
A = 16'h0022; B = 16'h00F9; #100;
A = 16'h0022; B = 16'h00FA; #100;
A = 16'h0022; B = 16'h00FB; #100;
A = 16'h0022; B = 16'h00FC; #100;
A = 16'h0022; B = 16'h00FD; #100;
A = 16'h0022; B = 16'h00FE; #100;
A = 16'h0022; B = 16'h00FF; #100;
A = 16'h0023; B = 16'h000; #100;
A = 16'h0023; B = 16'h001; #100;
A = 16'h0023; B = 16'h002; #100;
A = 16'h0023; B = 16'h003; #100;
A = 16'h0023; B = 16'h004; #100;
A = 16'h0023; B = 16'h005; #100;
A = 16'h0023; B = 16'h006; #100;
A = 16'h0023; B = 16'h007; #100;
A = 16'h0023; B = 16'h008; #100;
A = 16'h0023; B = 16'h009; #100;
A = 16'h0023; B = 16'h00A; #100;
A = 16'h0023; B = 16'h00B; #100;
A = 16'h0023; B = 16'h00C; #100;
A = 16'h0023; B = 16'h00D; #100;
A = 16'h0023; B = 16'h00E; #100;
A = 16'h0023; B = 16'h00F; #100;
A = 16'h0023; B = 16'h0010; #100;
A = 16'h0023; B = 16'h0011; #100;
A = 16'h0023; B = 16'h0012; #100;
A = 16'h0023; B = 16'h0013; #100;
A = 16'h0023; B = 16'h0014; #100;
A = 16'h0023; B = 16'h0015; #100;
A = 16'h0023; B = 16'h0016; #100;
A = 16'h0023; B = 16'h0017; #100;
A = 16'h0023; B = 16'h0018; #100;
A = 16'h0023; B = 16'h0019; #100;
A = 16'h0023; B = 16'h001A; #100;
A = 16'h0023; B = 16'h001B; #100;
A = 16'h0023; B = 16'h001C; #100;
A = 16'h0023; B = 16'h001D; #100;
A = 16'h0023; B = 16'h001E; #100;
A = 16'h0023; B = 16'h001F; #100;
A = 16'h0023; B = 16'h0020; #100;
A = 16'h0023; B = 16'h0021; #100;
A = 16'h0023; B = 16'h0022; #100;
A = 16'h0023; B = 16'h0023; #100;
A = 16'h0023; B = 16'h0024; #100;
A = 16'h0023; B = 16'h0025; #100;
A = 16'h0023; B = 16'h0026; #100;
A = 16'h0023; B = 16'h0027; #100;
A = 16'h0023; B = 16'h0028; #100;
A = 16'h0023; B = 16'h0029; #100;
A = 16'h0023; B = 16'h002A; #100;
A = 16'h0023; B = 16'h002B; #100;
A = 16'h0023; B = 16'h002C; #100;
A = 16'h0023; B = 16'h002D; #100;
A = 16'h0023; B = 16'h002E; #100;
A = 16'h0023; B = 16'h002F; #100;
A = 16'h0023; B = 16'h0030; #100;
A = 16'h0023; B = 16'h0031; #100;
A = 16'h0023; B = 16'h0032; #100;
A = 16'h0023; B = 16'h0033; #100;
A = 16'h0023; B = 16'h0034; #100;
A = 16'h0023; B = 16'h0035; #100;
A = 16'h0023; B = 16'h0036; #100;
A = 16'h0023; B = 16'h0037; #100;
A = 16'h0023; B = 16'h0038; #100;
A = 16'h0023; B = 16'h0039; #100;
A = 16'h0023; B = 16'h003A; #100;
A = 16'h0023; B = 16'h003B; #100;
A = 16'h0023; B = 16'h003C; #100;
A = 16'h0023; B = 16'h003D; #100;
A = 16'h0023; B = 16'h003E; #100;
A = 16'h0023; B = 16'h003F; #100;
A = 16'h0023; B = 16'h0040; #100;
A = 16'h0023; B = 16'h0041; #100;
A = 16'h0023; B = 16'h0042; #100;
A = 16'h0023; B = 16'h0043; #100;
A = 16'h0023; B = 16'h0044; #100;
A = 16'h0023; B = 16'h0045; #100;
A = 16'h0023; B = 16'h0046; #100;
A = 16'h0023; B = 16'h0047; #100;
A = 16'h0023; B = 16'h0048; #100;
A = 16'h0023; B = 16'h0049; #100;
A = 16'h0023; B = 16'h004A; #100;
A = 16'h0023; B = 16'h004B; #100;
A = 16'h0023; B = 16'h004C; #100;
A = 16'h0023; B = 16'h004D; #100;
A = 16'h0023; B = 16'h004E; #100;
A = 16'h0023; B = 16'h004F; #100;
A = 16'h0023; B = 16'h0050; #100;
A = 16'h0023; B = 16'h0051; #100;
A = 16'h0023; B = 16'h0052; #100;
A = 16'h0023; B = 16'h0053; #100;
A = 16'h0023; B = 16'h0054; #100;
A = 16'h0023; B = 16'h0055; #100;
A = 16'h0023; B = 16'h0056; #100;
A = 16'h0023; B = 16'h0057; #100;
A = 16'h0023; B = 16'h0058; #100;
A = 16'h0023; B = 16'h0059; #100;
A = 16'h0023; B = 16'h005A; #100;
A = 16'h0023; B = 16'h005B; #100;
A = 16'h0023; B = 16'h005C; #100;
A = 16'h0023; B = 16'h005D; #100;
A = 16'h0023; B = 16'h005E; #100;
A = 16'h0023; B = 16'h005F; #100;
A = 16'h0023; B = 16'h0060; #100;
A = 16'h0023; B = 16'h0061; #100;
A = 16'h0023; B = 16'h0062; #100;
A = 16'h0023; B = 16'h0063; #100;
A = 16'h0023; B = 16'h0064; #100;
A = 16'h0023; B = 16'h0065; #100;
A = 16'h0023; B = 16'h0066; #100;
A = 16'h0023; B = 16'h0067; #100;
A = 16'h0023; B = 16'h0068; #100;
A = 16'h0023; B = 16'h0069; #100;
A = 16'h0023; B = 16'h006A; #100;
A = 16'h0023; B = 16'h006B; #100;
A = 16'h0023; B = 16'h006C; #100;
A = 16'h0023; B = 16'h006D; #100;
A = 16'h0023; B = 16'h006E; #100;
A = 16'h0023; B = 16'h006F; #100;
A = 16'h0023; B = 16'h0070; #100;
A = 16'h0023; B = 16'h0071; #100;
A = 16'h0023; B = 16'h0072; #100;
A = 16'h0023; B = 16'h0073; #100;
A = 16'h0023; B = 16'h0074; #100;
A = 16'h0023; B = 16'h0075; #100;
A = 16'h0023; B = 16'h0076; #100;
A = 16'h0023; B = 16'h0077; #100;
A = 16'h0023; B = 16'h0078; #100;
A = 16'h0023; B = 16'h0079; #100;
A = 16'h0023; B = 16'h007A; #100;
A = 16'h0023; B = 16'h007B; #100;
A = 16'h0023; B = 16'h007C; #100;
A = 16'h0023; B = 16'h007D; #100;
A = 16'h0023; B = 16'h007E; #100;
A = 16'h0023; B = 16'h007F; #100;
A = 16'h0023; B = 16'h0080; #100;
A = 16'h0023; B = 16'h0081; #100;
A = 16'h0023; B = 16'h0082; #100;
A = 16'h0023; B = 16'h0083; #100;
A = 16'h0023; B = 16'h0084; #100;
A = 16'h0023; B = 16'h0085; #100;
A = 16'h0023; B = 16'h0086; #100;
A = 16'h0023; B = 16'h0087; #100;
A = 16'h0023; B = 16'h0088; #100;
A = 16'h0023; B = 16'h0089; #100;
A = 16'h0023; B = 16'h008A; #100;
A = 16'h0023; B = 16'h008B; #100;
A = 16'h0023; B = 16'h008C; #100;
A = 16'h0023; B = 16'h008D; #100;
A = 16'h0023; B = 16'h008E; #100;
A = 16'h0023; B = 16'h008F; #100;
A = 16'h0023; B = 16'h0090; #100;
A = 16'h0023; B = 16'h0091; #100;
A = 16'h0023; B = 16'h0092; #100;
A = 16'h0023; B = 16'h0093; #100;
A = 16'h0023; B = 16'h0094; #100;
A = 16'h0023; B = 16'h0095; #100;
A = 16'h0023; B = 16'h0096; #100;
A = 16'h0023; B = 16'h0097; #100;
A = 16'h0023; B = 16'h0098; #100;
A = 16'h0023; B = 16'h0099; #100;
A = 16'h0023; B = 16'h009A; #100;
A = 16'h0023; B = 16'h009B; #100;
A = 16'h0023; B = 16'h009C; #100;
A = 16'h0023; B = 16'h009D; #100;
A = 16'h0023; B = 16'h009E; #100;
A = 16'h0023; B = 16'h009F; #100;
A = 16'h0023; B = 16'h00A0; #100;
A = 16'h0023; B = 16'h00A1; #100;
A = 16'h0023; B = 16'h00A2; #100;
A = 16'h0023; B = 16'h00A3; #100;
A = 16'h0023; B = 16'h00A4; #100;
A = 16'h0023; B = 16'h00A5; #100;
A = 16'h0023; B = 16'h00A6; #100;
A = 16'h0023; B = 16'h00A7; #100;
A = 16'h0023; B = 16'h00A8; #100;
A = 16'h0023; B = 16'h00A9; #100;
A = 16'h0023; B = 16'h00AA; #100;
A = 16'h0023; B = 16'h00AB; #100;
A = 16'h0023; B = 16'h00AC; #100;
A = 16'h0023; B = 16'h00AD; #100;
A = 16'h0023; B = 16'h00AE; #100;
A = 16'h0023; B = 16'h00AF; #100;
A = 16'h0023; B = 16'h00B0; #100;
A = 16'h0023; B = 16'h00B1; #100;
A = 16'h0023; B = 16'h00B2; #100;
A = 16'h0023; B = 16'h00B3; #100;
A = 16'h0023; B = 16'h00B4; #100;
A = 16'h0023; B = 16'h00B5; #100;
A = 16'h0023; B = 16'h00B6; #100;
A = 16'h0023; B = 16'h00B7; #100;
A = 16'h0023; B = 16'h00B8; #100;
A = 16'h0023; B = 16'h00B9; #100;
A = 16'h0023; B = 16'h00BA; #100;
A = 16'h0023; B = 16'h00BB; #100;
A = 16'h0023; B = 16'h00BC; #100;
A = 16'h0023; B = 16'h00BD; #100;
A = 16'h0023; B = 16'h00BE; #100;
A = 16'h0023; B = 16'h00BF; #100;
A = 16'h0023; B = 16'h00C0; #100;
A = 16'h0023; B = 16'h00C1; #100;
A = 16'h0023; B = 16'h00C2; #100;
A = 16'h0023; B = 16'h00C3; #100;
A = 16'h0023; B = 16'h00C4; #100;
A = 16'h0023; B = 16'h00C5; #100;
A = 16'h0023; B = 16'h00C6; #100;
A = 16'h0023; B = 16'h00C7; #100;
A = 16'h0023; B = 16'h00C8; #100;
A = 16'h0023; B = 16'h00C9; #100;
A = 16'h0023; B = 16'h00CA; #100;
A = 16'h0023; B = 16'h00CB; #100;
A = 16'h0023; B = 16'h00CC; #100;
A = 16'h0023; B = 16'h00CD; #100;
A = 16'h0023; B = 16'h00CE; #100;
A = 16'h0023; B = 16'h00CF; #100;
A = 16'h0023; B = 16'h00D0; #100;
A = 16'h0023; B = 16'h00D1; #100;
A = 16'h0023; B = 16'h00D2; #100;
A = 16'h0023; B = 16'h00D3; #100;
A = 16'h0023; B = 16'h00D4; #100;
A = 16'h0023; B = 16'h00D5; #100;
A = 16'h0023; B = 16'h00D6; #100;
A = 16'h0023; B = 16'h00D7; #100;
A = 16'h0023; B = 16'h00D8; #100;
A = 16'h0023; B = 16'h00D9; #100;
A = 16'h0023; B = 16'h00DA; #100;
A = 16'h0023; B = 16'h00DB; #100;
A = 16'h0023; B = 16'h00DC; #100;
A = 16'h0023; B = 16'h00DD; #100;
A = 16'h0023; B = 16'h00DE; #100;
A = 16'h0023; B = 16'h00DF; #100;
A = 16'h0023; B = 16'h00E0; #100;
A = 16'h0023; B = 16'h00E1; #100;
A = 16'h0023; B = 16'h00E2; #100;
A = 16'h0023; B = 16'h00E3; #100;
A = 16'h0023; B = 16'h00E4; #100;
A = 16'h0023; B = 16'h00E5; #100;
A = 16'h0023; B = 16'h00E6; #100;
A = 16'h0023; B = 16'h00E7; #100;
A = 16'h0023; B = 16'h00E8; #100;
A = 16'h0023; B = 16'h00E9; #100;
A = 16'h0023; B = 16'h00EA; #100;
A = 16'h0023; B = 16'h00EB; #100;
A = 16'h0023; B = 16'h00EC; #100;
A = 16'h0023; B = 16'h00ED; #100;
A = 16'h0023; B = 16'h00EE; #100;
A = 16'h0023; B = 16'h00EF; #100;
A = 16'h0023; B = 16'h00F0; #100;
A = 16'h0023; B = 16'h00F1; #100;
A = 16'h0023; B = 16'h00F2; #100;
A = 16'h0023; B = 16'h00F3; #100;
A = 16'h0023; B = 16'h00F4; #100;
A = 16'h0023; B = 16'h00F5; #100;
A = 16'h0023; B = 16'h00F6; #100;
A = 16'h0023; B = 16'h00F7; #100;
A = 16'h0023; B = 16'h00F8; #100;
A = 16'h0023; B = 16'h00F9; #100;
A = 16'h0023; B = 16'h00FA; #100;
A = 16'h0023; B = 16'h00FB; #100;
A = 16'h0023; B = 16'h00FC; #100;
A = 16'h0023; B = 16'h00FD; #100;
A = 16'h0023; B = 16'h00FE; #100;
A = 16'h0023; B = 16'h00FF; #100;
A = 16'h0024; B = 16'h000; #100;
A = 16'h0024; B = 16'h001; #100;
A = 16'h0024; B = 16'h002; #100;
A = 16'h0024; B = 16'h003; #100;
A = 16'h0024; B = 16'h004; #100;
A = 16'h0024; B = 16'h005; #100;
A = 16'h0024; B = 16'h006; #100;
A = 16'h0024; B = 16'h007; #100;
A = 16'h0024; B = 16'h008; #100;
A = 16'h0024; B = 16'h009; #100;
A = 16'h0024; B = 16'h00A; #100;
A = 16'h0024; B = 16'h00B; #100;
A = 16'h0024; B = 16'h00C; #100;
A = 16'h0024; B = 16'h00D; #100;
A = 16'h0024; B = 16'h00E; #100;
A = 16'h0024; B = 16'h00F; #100;
A = 16'h0024; B = 16'h0010; #100;
A = 16'h0024; B = 16'h0011; #100;
A = 16'h0024; B = 16'h0012; #100;
A = 16'h0024; B = 16'h0013; #100;
A = 16'h0024; B = 16'h0014; #100;
A = 16'h0024; B = 16'h0015; #100;
A = 16'h0024; B = 16'h0016; #100;
A = 16'h0024; B = 16'h0017; #100;
A = 16'h0024; B = 16'h0018; #100;
A = 16'h0024; B = 16'h0019; #100;
A = 16'h0024; B = 16'h001A; #100;
A = 16'h0024; B = 16'h001B; #100;
A = 16'h0024; B = 16'h001C; #100;
A = 16'h0024; B = 16'h001D; #100;
A = 16'h0024; B = 16'h001E; #100;
A = 16'h0024; B = 16'h001F; #100;
A = 16'h0024; B = 16'h0020; #100;
A = 16'h0024; B = 16'h0021; #100;
A = 16'h0024; B = 16'h0022; #100;
A = 16'h0024; B = 16'h0023; #100;
A = 16'h0024; B = 16'h0024; #100;
A = 16'h0024; B = 16'h0025; #100;
A = 16'h0024; B = 16'h0026; #100;
A = 16'h0024; B = 16'h0027; #100;
A = 16'h0024; B = 16'h0028; #100;
A = 16'h0024; B = 16'h0029; #100;
A = 16'h0024; B = 16'h002A; #100;
A = 16'h0024; B = 16'h002B; #100;
A = 16'h0024; B = 16'h002C; #100;
A = 16'h0024; B = 16'h002D; #100;
A = 16'h0024; B = 16'h002E; #100;
A = 16'h0024; B = 16'h002F; #100;
A = 16'h0024; B = 16'h0030; #100;
A = 16'h0024; B = 16'h0031; #100;
A = 16'h0024; B = 16'h0032; #100;
A = 16'h0024; B = 16'h0033; #100;
A = 16'h0024; B = 16'h0034; #100;
A = 16'h0024; B = 16'h0035; #100;
A = 16'h0024; B = 16'h0036; #100;
A = 16'h0024; B = 16'h0037; #100;
A = 16'h0024; B = 16'h0038; #100;
A = 16'h0024; B = 16'h0039; #100;
A = 16'h0024; B = 16'h003A; #100;
A = 16'h0024; B = 16'h003B; #100;
A = 16'h0024; B = 16'h003C; #100;
A = 16'h0024; B = 16'h003D; #100;
A = 16'h0024; B = 16'h003E; #100;
A = 16'h0024; B = 16'h003F; #100;
A = 16'h0024; B = 16'h0040; #100;
A = 16'h0024; B = 16'h0041; #100;
A = 16'h0024; B = 16'h0042; #100;
A = 16'h0024; B = 16'h0043; #100;
A = 16'h0024; B = 16'h0044; #100;
A = 16'h0024; B = 16'h0045; #100;
A = 16'h0024; B = 16'h0046; #100;
A = 16'h0024; B = 16'h0047; #100;
A = 16'h0024; B = 16'h0048; #100;
A = 16'h0024; B = 16'h0049; #100;
A = 16'h0024; B = 16'h004A; #100;
A = 16'h0024; B = 16'h004B; #100;
A = 16'h0024; B = 16'h004C; #100;
A = 16'h0024; B = 16'h004D; #100;
A = 16'h0024; B = 16'h004E; #100;
A = 16'h0024; B = 16'h004F; #100;
A = 16'h0024; B = 16'h0050; #100;
A = 16'h0024; B = 16'h0051; #100;
A = 16'h0024; B = 16'h0052; #100;
A = 16'h0024; B = 16'h0053; #100;
A = 16'h0024; B = 16'h0054; #100;
A = 16'h0024; B = 16'h0055; #100;
A = 16'h0024; B = 16'h0056; #100;
A = 16'h0024; B = 16'h0057; #100;
A = 16'h0024; B = 16'h0058; #100;
A = 16'h0024; B = 16'h0059; #100;
A = 16'h0024; B = 16'h005A; #100;
A = 16'h0024; B = 16'h005B; #100;
A = 16'h0024; B = 16'h005C; #100;
A = 16'h0024; B = 16'h005D; #100;
A = 16'h0024; B = 16'h005E; #100;
A = 16'h0024; B = 16'h005F; #100;
A = 16'h0024; B = 16'h0060; #100;
A = 16'h0024; B = 16'h0061; #100;
A = 16'h0024; B = 16'h0062; #100;
A = 16'h0024; B = 16'h0063; #100;
A = 16'h0024; B = 16'h0064; #100;
A = 16'h0024; B = 16'h0065; #100;
A = 16'h0024; B = 16'h0066; #100;
A = 16'h0024; B = 16'h0067; #100;
A = 16'h0024; B = 16'h0068; #100;
A = 16'h0024; B = 16'h0069; #100;
A = 16'h0024; B = 16'h006A; #100;
A = 16'h0024; B = 16'h006B; #100;
A = 16'h0024; B = 16'h006C; #100;
A = 16'h0024; B = 16'h006D; #100;
A = 16'h0024; B = 16'h006E; #100;
A = 16'h0024; B = 16'h006F; #100;
A = 16'h0024; B = 16'h0070; #100;
A = 16'h0024; B = 16'h0071; #100;
A = 16'h0024; B = 16'h0072; #100;
A = 16'h0024; B = 16'h0073; #100;
A = 16'h0024; B = 16'h0074; #100;
A = 16'h0024; B = 16'h0075; #100;
A = 16'h0024; B = 16'h0076; #100;
A = 16'h0024; B = 16'h0077; #100;
A = 16'h0024; B = 16'h0078; #100;
A = 16'h0024; B = 16'h0079; #100;
A = 16'h0024; B = 16'h007A; #100;
A = 16'h0024; B = 16'h007B; #100;
A = 16'h0024; B = 16'h007C; #100;
A = 16'h0024; B = 16'h007D; #100;
A = 16'h0024; B = 16'h007E; #100;
A = 16'h0024; B = 16'h007F; #100;
A = 16'h0024; B = 16'h0080; #100;
A = 16'h0024; B = 16'h0081; #100;
A = 16'h0024; B = 16'h0082; #100;
A = 16'h0024; B = 16'h0083; #100;
A = 16'h0024; B = 16'h0084; #100;
A = 16'h0024; B = 16'h0085; #100;
A = 16'h0024; B = 16'h0086; #100;
A = 16'h0024; B = 16'h0087; #100;
A = 16'h0024; B = 16'h0088; #100;
A = 16'h0024; B = 16'h0089; #100;
A = 16'h0024; B = 16'h008A; #100;
A = 16'h0024; B = 16'h008B; #100;
A = 16'h0024; B = 16'h008C; #100;
A = 16'h0024; B = 16'h008D; #100;
A = 16'h0024; B = 16'h008E; #100;
A = 16'h0024; B = 16'h008F; #100;
A = 16'h0024; B = 16'h0090; #100;
A = 16'h0024; B = 16'h0091; #100;
A = 16'h0024; B = 16'h0092; #100;
A = 16'h0024; B = 16'h0093; #100;
A = 16'h0024; B = 16'h0094; #100;
A = 16'h0024; B = 16'h0095; #100;
A = 16'h0024; B = 16'h0096; #100;
A = 16'h0024; B = 16'h0097; #100;
A = 16'h0024; B = 16'h0098; #100;
A = 16'h0024; B = 16'h0099; #100;
A = 16'h0024; B = 16'h009A; #100;
A = 16'h0024; B = 16'h009B; #100;
A = 16'h0024; B = 16'h009C; #100;
A = 16'h0024; B = 16'h009D; #100;
A = 16'h0024; B = 16'h009E; #100;
A = 16'h0024; B = 16'h009F; #100;
A = 16'h0024; B = 16'h00A0; #100;
A = 16'h0024; B = 16'h00A1; #100;
A = 16'h0024; B = 16'h00A2; #100;
A = 16'h0024; B = 16'h00A3; #100;
A = 16'h0024; B = 16'h00A4; #100;
A = 16'h0024; B = 16'h00A5; #100;
A = 16'h0024; B = 16'h00A6; #100;
A = 16'h0024; B = 16'h00A7; #100;
A = 16'h0024; B = 16'h00A8; #100;
A = 16'h0024; B = 16'h00A9; #100;
A = 16'h0024; B = 16'h00AA; #100;
A = 16'h0024; B = 16'h00AB; #100;
A = 16'h0024; B = 16'h00AC; #100;
A = 16'h0024; B = 16'h00AD; #100;
A = 16'h0024; B = 16'h00AE; #100;
A = 16'h0024; B = 16'h00AF; #100;
A = 16'h0024; B = 16'h00B0; #100;
A = 16'h0024; B = 16'h00B1; #100;
A = 16'h0024; B = 16'h00B2; #100;
A = 16'h0024; B = 16'h00B3; #100;
A = 16'h0024; B = 16'h00B4; #100;
A = 16'h0024; B = 16'h00B5; #100;
A = 16'h0024; B = 16'h00B6; #100;
A = 16'h0024; B = 16'h00B7; #100;
A = 16'h0024; B = 16'h00B8; #100;
A = 16'h0024; B = 16'h00B9; #100;
A = 16'h0024; B = 16'h00BA; #100;
A = 16'h0024; B = 16'h00BB; #100;
A = 16'h0024; B = 16'h00BC; #100;
A = 16'h0024; B = 16'h00BD; #100;
A = 16'h0024; B = 16'h00BE; #100;
A = 16'h0024; B = 16'h00BF; #100;
A = 16'h0024; B = 16'h00C0; #100;
A = 16'h0024; B = 16'h00C1; #100;
A = 16'h0024; B = 16'h00C2; #100;
A = 16'h0024; B = 16'h00C3; #100;
A = 16'h0024; B = 16'h00C4; #100;
A = 16'h0024; B = 16'h00C5; #100;
A = 16'h0024; B = 16'h00C6; #100;
A = 16'h0024; B = 16'h00C7; #100;
A = 16'h0024; B = 16'h00C8; #100;
A = 16'h0024; B = 16'h00C9; #100;
A = 16'h0024; B = 16'h00CA; #100;
A = 16'h0024; B = 16'h00CB; #100;
A = 16'h0024; B = 16'h00CC; #100;
A = 16'h0024; B = 16'h00CD; #100;
A = 16'h0024; B = 16'h00CE; #100;
A = 16'h0024; B = 16'h00CF; #100;
A = 16'h0024; B = 16'h00D0; #100;
A = 16'h0024; B = 16'h00D1; #100;
A = 16'h0024; B = 16'h00D2; #100;
A = 16'h0024; B = 16'h00D3; #100;
A = 16'h0024; B = 16'h00D4; #100;
A = 16'h0024; B = 16'h00D5; #100;
A = 16'h0024; B = 16'h00D6; #100;
A = 16'h0024; B = 16'h00D7; #100;
A = 16'h0024; B = 16'h00D8; #100;
A = 16'h0024; B = 16'h00D9; #100;
A = 16'h0024; B = 16'h00DA; #100;
A = 16'h0024; B = 16'h00DB; #100;
A = 16'h0024; B = 16'h00DC; #100;
A = 16'h0024; B = 16'h00DD; #100;
A = 16'h0024; B = 16'h00DE; #100;
A = 16'h0024; B = 16'h00DF; #100;
A = 16'h0024; B = 16'h00E0; #100;
A = 16'h0024; B = 16'h00E1; #100;
A = 16'h0024; B = 16'h00E2; #100;
A = 16'h0024; B = 16'h00E3; #100;
A = 16'h0024; B = 16'h00E4; #100;
A = 16'h0024; B = 16'h00E5; #100;
A = 16'h0024; B = 16'h00E6; #100;
A = 16'h0024; B = 16'h00E7; #100;
A = 16'h0024; B = 16'h00E8; #100;
A = 16'h0024; B = 16'h00E9; #100;
A = 16'h0024; B = 16'h00EA; #100;
A = 16'h0024; B = 16'h00EB; #100;
A = 16'h0024; B = 16'h00EC; #100;
A = 16'h0024; B = 16'h00ED; #100;
A = 16'h0024; B = 16'h00EE; #100;
A = 16'h0024; B = 16'h00EF; #100;
A = 16'h0024; B = 16'h00F0; #100;
A = 16'h0024; B = 16'h00F1; #100;
A = 16'h0024; B = 16'h00F2; #100;
A = 16'h0024; B = 16'h00F3; #100;
A = 16'h0024; B = 16'h00F4; #100;
A = 16'h0024; B = 16'h00F5; #100;
A = 16'h0024; B = 16'h00F6; #100;
A = 16'h0024; B = 16'h00F7; #100;
A = 16'h0024; B = 16'h00F8; #100;
A = 16'h0024; B = 16'h00F9; #100;
A = 16'h0024; B = 16'h00FA; #100;
A = 16'h0024; B = 16'h00FB; #100;
A = 16'h0024; B = 16'h00FC; #100;
A = 16'h0024; B = 16'h00FD; #100;
A = 16'h0024; B = 16'h00FE; #100;
A = 16'h0024; B = 16'h00FF; #100;
A = 16'h0025; B = 16'h000; #100;
A = 16'h0025; B = 16'h001; #100;
A = 16'h0025; B = 16'h002; #100;
A = 16'h0025; B = 16'h003; #100;
A = 16'h0025; B = 16'h004; #100;
A = 16'h0025; B = 16'h005; #100;
A = 16'h0025; B = 16'h006; #100;
A = 16'h0025; B = 16'h007; #100;
A = 16'h0025; B = 16'h008; #100;
A = 16'h0025; B = 16'h009; #100;
A = 16'h0025; B = 16'h00A; #100;
A = 16'h0025; B = 16'h00B; #100;
A = 16'h0025; B = 16'h00C; #100;
A = 16'h0025; B = 16'h00D; #100;
A = 16'h0025; B = 16'h00E; #100;
A = 16'h0025; B = 16'h00F; #100;
A = 16'h0025; B = 16'h0010; #100;
A = 16'h0025; B = 16'h0011; #100;
A = 16'h0025; B = 16'h0012; #100;
A = 16'h0025; B = 16'h0013; #100;
A = 16'h0025; B = 16'h0014; #100;
A = 16'h0025; B = 16'h0015; #100;
A = 16'h0025; B = 16'h0016; #100;
A = 16'h0025; B = 16'h0017; #100;
A = 16'h0025; B = 16'h0018; #100;
A = 16'h0025; B = 16'h0019; #100;
A = 16'h0025; B = 16'h001A; #100;
A = 16'h0025; B = 16'h001B; #100;
A = 16'h0025; B = 16'h001C; #100;
A = 16'h0025; B = 16'h001D; #100;
A = 16'h0025; B = 16'h001E; #100;
A = 16'h0025; B = 16'h001F; #100;
A = 16'h0025; B = 16'h0020; #100;
A = 16'h0025; B = 16'h0021; #100;
A = 16'h0025; B = 16'h0022; #100;
A = 16'h0025; B = 16'h0023; #100;
A = 16'h0025; B = 16'h0024; #100;
A = 16'h0025; B = 16'h0025; #100;
A = 16'h0025; B = 16'h0026; #100;
A = 16'h0025; B = 16'h0027; #100;
A = 16'h0025; B = 16'h0028; #100;
A = 16'h0025; B = 16'h0029; #100;
A = 16'h0025; B = 16'h002A; #100;
A = 16'h0025; B = 16'h002B; #100;
A = 16'h0025; B = 16'h002C; #100;
A = 16'h0025; B = 16'h002D; #100;
A = 16'h0025; B = 16'h002E; #100;
A = 16'h0025; B = 16'h002F; #100;
A = 16'h0025; B = 16'h0030; #100;
A = 16'h0025; B = 16'h0031; #100;
A = 16'h0025; B = 16'h0032; #100;
A = 16'h0025; B = 16'h0033; #100;
A = 16'h0025; B = 16'h0034; #100;
A = 16'h0025; B = 16'h0035; #100;
A = 16'h0025; B = 16'h0036; #100;
A = 16'h0025; B = 16'h0037; #100;
A = 16'h0025; B = 16'h0038; #100;
A = 16'h0025; B = 16'h0039; #100;
A = 16'h0025; B = 16'h003A; #100;
A = 16'h0025; B = 16'h003B; #100;
A = 16'h0025; B = 16'h003C; #100;
A = 16'h0025; B = 16'h003D; #100;
A = 16'h0025; B = 16'h003E; #100;
A = 16'h0025; B = 16'h003F; #100;
A = 16'h0025; B = 16'h0040; #100;
A = 16'h0025; B = 16'h0041; #100;
A = 16'h0025; B = 16'h0042; #100;
A = 16'h0025; B = 16'h0043; #100;
A = 16'h0025; B = 16'h0044; #100;
A = 16'h0025; B = 16'h0045; #100;
A = 16'h0025; B = 16'h0046; #100;
A = 16'h0025; B = 16'h0047; #100;
A = 16'h0025; B = 16'h0048; #100;
A = 16'h0025; B = 16'h0049; #100;
A = 16'h0025; B = 16'h004A; #100;
A = 16'h0025; B = 16'h004B; #100;
A = 16'h0025; B = 16'h004C; #100;
A = 16'h0025; B = 16'h004D; #100;
A = 16'h0025; B = 16'h004E; #100;
A = 16'h0025; B = 16'h004F; #100;
A = 16'h0025; B = 16'h0050; #100;
A = 16'h0025; B = 16'h0051; #100;
A = 16'h0025; B = 16'h0052; #100;
A = 16'h0025; B = 16'h0053; #100;
A = 16'h0025; B = 16'h0054; #100;
A = 16'h0025; B = 16'h0055; #100;
A = 16'h0025; B = 16'h0056; #100;
A = 16'h0025; B = 16'h0057; #100;
A = 16'h0025; B = 16'h0058; #100;
A = 16'h0025; B = 16'h0059; #100;
A = 16'h0025; B = 16'h005A; #100;
A = 16'h0025; B = 16'h005B; #100;
A = 16'h0025; B = 16'h005C; #100;
A = 16'h0025; B = 16'h005D; #100;
A = 16'h0025; B = 16'h005E; #100;
A = 16'h0025; B = 16'h005F; #100;
A = 16'h0025; B = 16'h0060; #100;
A = 16'h0025; B = 16'h0061; #100;
A = 16'h0025; B = 16'h0062; #100;
A = 16'h0025; B = 16'h0063; #100;
A = 16'h0025; B = 16'h0064; #100;
A = 16'h0025; B = 16'h0065; #100;
A = 16'h0025; B = 16'h0066; #100;
A = 16'h0025; B = 16'h0067; #100;
A = 16'h0025; B = 16'h0068; #100;
A = 16'h0025; B = 16'h0069; #100;
A = 16'h0025; B = 16'h006A; #100;
A = 16'h0025; B = 16'h006B; #100;
A = 16'h0025; B = 16'h006C; #100;
A = 16'h0025; B = 16'h006D; #100;
A = 16'h0025; B = 16'h006E; #100;
A = 16'h0025; B = 16'h006F; #100;
A = 16'h0025; B = 16'h0070; #100;
A = 16'h0025; B = 16'h0071; #100;
A = 16'h0025; B = 16'h0072; #100;
A = 16'h0025; B = 16'h0073; #100;
A = 16'h0025; B = 16'h0074; #100;
A = 16'h0025; B = 16'h0075; #100;
A = 16'h0025; B = 16'h0076; #100;
A = 16'h0025; B = 16'h0077; #100;
A = 16'h0025; B = 16'h0078; #100;
A = 16'h0025; B = 16'h0079; #100;
A = 16'h0025; B = 16'h007A; #100;
A = 16'h0025; B = 16'h007B; #100;
A = 16'h0025; B = 16'h007C; #100;
A = 16'h0025; B = 16'h007D; #100;
A = 16'h0025; B = 16'h007E; #100;
A = 16'h0025; B = 16'h007F; #100;
A = 16'h0025; B = 16'h0080; #100;
A = 16'h0025; B = 16'h0081; #100;
A = 16'h0025; B = 16'h0082; #100;
A = 16'h0025; B = 16'h0083; #100;
A = 16'h0025; B = 16'h0084; #100;
A = 16'h0025; B = 16'h0085; #100;
A = 16'h0025; B = 16'h0086; #100;
A = 16'h0025; B = 16'h0087; #100;
A = 16'h0025; B = 16'h0088; #100;
A = 16'h0025; B = 16'h0089; #100;
A = 16'h0025; B = 16'h008A; #100;
A = 16'h0025; B = 16'h008B; #100;
A = 16'h0025; B = 16'h008C; #100;
A = 16'h0025; B = 16'h008D; #100;
A = 16'h0025; B = 16'h008E; #100;
A = 16'h0025; B = 16'h008F; #100;
A = 16'h0025; B = 16'h0090; #100;
A = 16'h0025; B = 16'h0091; #100;
A = 16'h0025; B = 16'h0092; #100;
A = 16'h0025; B = 16'h0093; #100;
A = 16'h0025; B = 16'h0094; #100;
A = 16'h0025; B = 16'h0095; #100;
A = 16'h0025; B = 16'h0096; #100;
A = 16'h0025; B = 16'h0097; #100;
A = 16'h0025; B = 16'h0098; #100;
A = 16'h0025; B = 16'h0099; #100;
A = 16'h0025; B = 16'h009A; #100;
A = 16'h0025; B = 16'h009B; #100;
A = 16'h0025; B = 16'h009C; #100;
A = 16'h0025; B = 16'h009D; #100;
A = 16'h0025; B = 16'h009E; #100;
A = 16'h0025; B = 16'h009F; #100;
A = 16'h0025; B = 16'h00A0; #100;
A = 16'h0025; B = 16'h00A1; #100;
A = 16'h0025; B = 16'h00A2; #100;
A = 16'h0025; B = 16'h00A3; #100;
A = 16'h0025; B = 16'h00A4; #100;
A = 16'h0025; B = 16'h00A5; #100;
A = 16'h0025; B = 16'h00A6; #100;
A = 16'h0025; B = 16'h00A7; #100;
A = 16'h0025; B = 16'h00A8; #100;
A = 16'h0025; B = 16'h00A9; #100;
A = 16'h0025; B = 16'h00AA; #100;
A = 16'h0025; B = 16'h00AB; #100;
A = 16'h0025; B = 16'h00AC; #100;
A = 16'h0025; B = 16'h00AD; #100;
A = 16'h0025; B = 16'h00AE; #100;
A = 16'h0025; B = 16'h00AF; #100;
A = 16'h0025; B = 16'h00B0; #100;
A = 16'h0025; B = 16'h00B1; #100;
A = 16'h0025; B = 16'h00B2; #100;
A = 16'h0025; B = 16'h00B3; #100;
A = 16'h0025; B = 16'h00B4; #100;
A = 16'h0025; B = 16'h00B5; #100;
A = 16'h0025; B = 16'h00B6; #100;
A = 16'h0025; B = 16'h00B7; #100;
A = 16'h0025; B = 16'h00B8; #100;
A = 16'h0025; B = 16'h00B9; #100;
A = 16'h0025; B = 16'h00BA; #100;
A = 16'h0025; B = 16'h00BB; #100;
A = 16'h0025; B = 16'h00BC; #100;
A = 16'h0025; B = 16'h00BD; #100;
A = 16'h0025; B = 16'h00BE; #100;
A = 16'h0025; B = 16'h00BF; #100;
A = 16'h0025; B = 16'h00C0; #100;
A = 16'h0025; B = 16'h00C1; #100;
A = 16'h0025; B = 16'h00C2; #100;
A = 16'h0025; B = 16'h00C3; #100;
A = 16'h0025; B = 16'h00C4; #100;
A = 16'h0025; B = 16'h00C5; #100;
A = 16'h0025; B = 16'h00C6; #100;
A = 16'h0025; B = 16'h00C7; #100;
A = 16'h0025; B = 16'h00C8; #100;
A = 16'h0025; B = 16'h00C9; #100;
A = 16'h0025; B = 16'h00CA; #100;
A = 16'h0025; B = 16'h00CB; #100;
A = 16'h0025; B = 16'h00CC; #100;
A = 16'h0025; B = 16'h00CD; #100;
A = 16'h0025; B = 16'h00CE; #100;
A = 16'h0025; B = 16'h00CF; #100;
A = 16'h0025; B = 16'h00D0; #100;
A = 16'h0025; B = 16'h00D1; #100;
A = 16'h0025; B = 16'h00D2; #100;
A = 16'h0025; B = 16'h00D3; #100;
A = 16'h0025; B = 16'h00D4; #100;
A = 16'h0025; B = 16'h00D5; #100;
A = 16'h0025; B = 16'h00D6; #100;
A = 16'h0025; B = 16'h00D7; #100;
A = 16'h0025; B = 16'h00D8; #100;
A = 16'h0025; B = 16'h00D9; #100;
A = 16'h0025; B = 16'h00DA; #100;
A = 16'h0025; B = 16'h00DB; #100;
A = 16'h0025; B = 16'h00DC; #100;
A = 16'h0025; B = 16'h00DD; #100;
A = 16'h0025; B = 16'h00DE; #100;
A = 16'h0025; B = 16'h00DF; #100;
A = 16'h0025; B = 16'h00E0; #100;
A = 16'h0025; B = 16'h00E1; #100;
A = 16'h0025; B = 16'h00E2; #100;
A = 16'h0025; B = 16'h00E3; #100;
A = 16'h0025; B = 16'h00E4; #100;
A = 16'h0025; B = 16'h00E5; #100;
A = 16'h0025; B = 16'h00E6; #100;
A = 16'h0025; B = 16'h00E7; #100;
A = 16'h0025; B = 16'h00E8; #100;
A = 16'h0025; B = 16'h00E9; #100;
A = 16'h0025; B = 16'h00EA; #100;
A = 16'h0025; B = 16'h00EB; #100;
A = 16'h0025; B = 16'h00EC; #100;
A = 16'h0025; B = 16'h00ED; #100;
A = 16'h0025; B = 16'h00EE; #100;
A = 16'h0025; B = 16'h00EF; #100;
A = 16'h0025; B = 16'h00F0; #100;
A = 16'h0025; B = 16'h00F1; #100;
A = 16'h0025; B = 16'h00F2; #100;
A = 16'h0025; B = 16'h00F3; #100;
A = 16'h0025; B = 16'h00F4; #100;
A = 16'h0025; B = 16'h00F5; #100;
A = 16'h0025; B = 16'h00F6; #100;
A = 16'h0025; B = 16'h00F7; #100;
A = 16'h0025; B = 16'h00F8; #100;
A = 16'h0025; B = 16'h00F9; #100;
A = 16'h0025; B = 16'h00FA; #100;
A = 16'h0025; B = 16'h00FB; #100;
A = 16'h0025; B = 16'h00FC; #100;
A = 16'h0025; B = 16'h00FD; #100;
A = 16'h0025; B = 16'h00FE; #100;
A = 16'h0025; B = 16'h00FF; #100;
A = 16'h0026; B = 16'h000; #100;
A = 16'h0026; B = 16'h001; #100;
A = 16'h0026; B = 16'h002; #100;
A = 16'h0026; B = 16'h003; #100;
A = 16'h0026; B = 16'h004; #100;
A = 16'h0026; B = 16'h005; #100;
A = 16'h0026; B = 16'h006; #100;
A = 16'h0026; B = 16'h007; #100;
A = 16'h0026; B = 16'h008; #100;
A = 16'h0026; B = 16'h009; #100;
A = 16'h0026; B = 16'h00A; #100;
A = 16'h0026; B = 16'h00B; #100;
A = 16'h0026; B = 16'h00C; #100;
A = 16'h0026; B = 16'h00D; #100;
A = 16'h0026; B = 16'h00E; #100;
A = 16'h0026; B = 16'h00F; #100;
A = 16'h0026; B = 16'h0010; #100;
A = 16'h0026; B = 16'h0011; #100;
A = 16'h0026; B = 16'h0012; #100;
A = 16'h0026; B = 16'h0013; #100;
A = 16'h0026; B = 16'h0014; #100;
A = 16'h0026; B = 16'h0015; #100;
A = 16'h0026; B = 16'h0016; #100;
A = 16'h0026; B = 16'h0017; #100;
A = 16'h0026; B = 16'h0018; #100;
A = 16'h0026; B = 16'h0019; #100;
A = 16'h0026; B = 16'h001A; #100;
A = 16'h0026; B = 16'h001B; #100;
A = 16'h0026; B = 16'h001C; #100;
A = 16'h0026; B = 16'h001D; #100;
A = 16'h0026; B = 16'h001E; #100;
A = 16'h0026; B = 16'h001F; #100;
A = 16'h0026; B = 16'h0020; #100;
A = 16'h0026; B = 16'h0021; #100;
A = 16'h0026; B = 16'h0022; #100;
A = 16'h0026; B = 16'h0023; #100;
A = 16'h0026; B = 16'h0024; #100;
A = 16'h0026; B = 16'h0025; #100;
A = 16'h0026; B = 16'h0026; #100;
A = 16'h0026; B = 16'h0027; #100;
A = 16'h0026; B = 16'h0028; #100;
A = 16'h0026; B = 16'h0029; #100;
A = 16'h0026; B = 16'h002A; #100;
A = 16'h0026; B = 16'h002B; #100;
A = 16'h0026; B = 16'h002C; #100;
A = 16'h0026; B = 16'h002D; #100;
A = 16'h0026; B = 16'h002E; #100;
A = 16'h0026; B = 16'h002F; #100;
A = 16'h0026; B = 16'h0030; #100;
A = 16'h0026; B = 16'h0031; #100;
A = 16'h0026; B = 16'h0032; #100;
A = 16'h0026; B = 16'h0033; #100;
A = 16'h0026; B = 16'h0034; #100;
A = 16'h0026; B = 16'h0035; #100;
A = 16'h0026; B = 16'h0036; #100;
A = 16'h0026; B = 16'h0037; #100;
A = 16'h0026; B = 16'h0038; #100;
A = 16'h0026; B = 16'h0039; #100;
A = 16'h0026; B = 16'h003A; #100;
A = 16'h0026; B = 16'h003B; #100;
A = 16'h0026; B = 16'h003C; #100;
A = 16'h0026; B = 16'h003D; #100;
A = 16'h0026; B = 16'h003E; #100;
A = 16'h0026; B = 16'h003F; #100;
A = 16'h0026; B = 16'h0040; #100;
A = 16'h0026; B = 16'h0041; #100;
A = 16'h0026; B = 16'h0042; #100;
A = 16'h0026; B = 16'h0043; #100;
A = 16'h0026; B = 16'h0044; #100;
A = 16'h0026; B = 16'h0045; #100;
A = 16'h0026; B = 16'h0046; #100;
A = 16'h0026; B = 16'h0047; #100;
A = 16'h0026; B = 16'h0048; #100;
A = 16'h0026; B = 16'h0049; #100;
A = 16'h0026; B = 16'h004A; #100;
A = 16'h0026; B = 16'h004B; #100;
A = 16'h0026; B = 16'h004C; #100;
A = 16'h0026; B = 16'h004D; #100;
A = 16'h0026; B = 16'h004E; #100;
A = 16'h0026; B = 16'h004F; #100;
A = 16'h0026; B = 16'h0050; #100;
A = 16'h0026; B = 16'h0051; #100;
A = 16'h0026; B = 16'h0052; #100;
A = 16'h0026; B = 16'h0053; #100;
A = 16'h0026; B = 16'h0054; #100;
A = 16'h0026; B = 16'h0055; #100;
A = 16'h0026; B = 16'h0056; #100;
A = 16'h0026; B = 16'h0057; #100;
A = 16'h0026; B = 16'h0058; #100;
A = 16'h0026; B = 16'h0059; #100;
A = 16'h0026; B = 16'h005A; #100;
A = 16'h0026; B = 16'h005B; #100;
A = 16'h0026; B = 16'h005C; #100;
A = 16'h0026; B = 16'h005D; #100;
A = 16'h0026; B = 16'h005E; #100;
A = 16'h0026; B = 16'h005F; #100;
A = 16'h0026; B = 16'h0060; #100;
A = 16'h0026; B = 16'h0061; #100;
A = 16'h0026; B = 16'h0062; #100;
A = 16'h0026; B = 16'h0063; #100;
A = 16'h0026; B = 16'h0064; #100;
A = 16'h0026; B = 16'h0065; #100;
A = 16'h0026; B = 16'h0066; #100;
A = 16'h0026; B = 16'h0067; #100;
A = 16'h0026; B = 16'h0068; #100;
A = 16'h0026; B = 16'h0069; #100;
A = 16'h0026; B = 16'h006A; #100;
A = 16'h0026; B = 16'h006B; #100;
A = 16'h0026; B = 16'h006C; #100;
A = 16'h0026; B = 16'h006D; #100;
A = 16'h0026; B = 16'h006E; #100;
A = 16'h0026; B = 16'h006F; #100;
A = 16'h0026; B = 16'h0070; #100;
A = 16'h0026; B = 16'h0071; #100;
A = 16'h0026; B = 16'h0072; #100;
A = 16'h0026; B = 16'h0073; #100;
A = 16'h0026; B = 16'h0074; #100;
A = 16'h0026; B = 16'h0075; #100;
A = 16'h0026; B = 16'h0076; #100;
A = 16'h0026; B = 16'h0077; #100;
A = 16'h0026; B = 16'h0078; #100;
A = 16'h0026; B = 16'h0079; #100;
A = 16'h0026; B = 16'h007A; #100;
A = 16'h0026; B = 16'h007B; #100;
A = 16'h0026; B = 16'h007C; #100;
A = 16'h0026; B = 16'h007D; #100;
A = 16'h0026; B = 16'h007E; #100;
A = 16'h0026; B = 16'h007F; #100;
A = 16'h0026; B = 16'h0080; #100;
A = 16'h0026; B = 16'h0081; #100;
A = 16'h0026; B = 16'h0082; #100;
A = 16'h0026; B = 16'h0083; #100;
A = 16'h0026; B = 16'h0084; #100;
A = 16'h0026; B = 16'h0085; #100;
A = 16'h0026; B = 16'h0086; #100;
A = 16'h0026; B = 16'h0087; #100;
A = 16'h0026; B = 16'h0088; #100;
A = 16'h0026; B = 16'h0089; #100;
A = 16'h0026; B = 16'h008A; #100;
A = 16'h0026; B = 16'h008B; #100;
A = 16'h0026; B = 16'h008C; #100;
A = 16'h0026; B = 16'h008D; #100;
A = 16'h0026; B = 16'h008E; #100;
A = 16'h0026; B = 16'h008F; #100;
A = 16'h0026; B = 16'h0090; #100;
A = 16'h0026; B = 16'h0091; #100;
A = 16'h0026; B = 16'h0092; #100;
A = 16'h0026; B = 16'h0093; #100;
A = 16'h0026; B = 16'h0094; #100;
A = 16'h0026; B = 16'h0095; #100;
A = 16'h0026; B = 16'h0096; #100;
A = 16'h0026; B = 16'h0097; #100;
A = 16'h0026; B = 16'h0098; #100;
A = 16'h0026; B = 16'h0099; #100;
A = 16'h0026; B = 16'h009A; #100;
A = 16'h0026; B = 16'h009B; #100;
A = 16'h0026; B = 16'h009C; #100;
A = 16'h0026; B = 16'h009D; #100;
A = 16'h0026; B = 16'h009E; #100;
A = 16'h0026; B = 16'h009F; #100;
A = 16'h0026; B = 16'h00A0; #100;
A = 16'h0026; B = 16'h00A1; #100;
A = 16'h0026; B = 16'h00A2; #100;
A = 16'h0026; B = 16'h00A3; #100;
A = 16'h0026; B = 16'h00A4; #100;
A = 16'h0026; B = 16'h00A5; #100;
A = 16'h0026; B = 16'h00A6; #100;
A = 16'h0026; B = 16'h00A7; #100;
A = 16'h0026; B = 16'h00A8; #100;
A = 16'h0026; B = 16'h00A9; #100;
A = 16'h0026; B = 16'h00AA; #100;
A = 16'h0026; B = 16'h00AB; #100;
A = 16'h0026; B = 16'h00AC; #100;
A = 16'h0026; B = 16'h00AD; #100;
A = 16'h0026; B = 16'h00AE; #100;
A = 16'h0026; B = 16'h00AF; #100;
A = 16'h0026; B = 16'h00B0; #100;
A = 16'h0026; B = 16'h00B1; #100;
A = 16'h0026; B = 16'h00B2; #100;
A = 16'h0026; B = 16'h00B3; #100;
A = 16'h0026; B = 16'h00B4; #100;
A = 16'h0026; B = 16'h00B5; #100;
A = 16'h0026; B = 16'h00B6; #100;
A = 16'h0026; B = 16'h00B7; #100;
A = 16'h0026; B = 16'h00B8; #100;
A = 16'h0026; B = 16'h00B9; #100;
A = 16'h0026; B = 16'h00BA; #100;
A = 16'h0026; B = 16'h00BB; #100;
A = 16'h0026; B = 16'h00BC; #100;
A = 16'h0026; B = 16'h00BD; #100;
A = 16'h0026; B = 16'h00BE; #100;
A = 16'h0026; B = 16'h00BF; #100;
A = 16'h0026; B = 16'h00C0; #100;
A = 16'h0026; B = 16'h00C1; #100;
A = 16'h0026; B = 16'h00C2; #100;
A = 16'h0026; B = 16'h00C3; #100;
A = 16'h0026; B = 16'h00C4; #100;
A = 16'h0026; B = 16'h00C5; #100;
A = 16'h0026; B = 16'h00C6; #100;
A = 16'h0026; B = 16'h00C7; #100;
A = 16'h0026; B = 16'h00C8; #100;
A = 16'h0026; B = 16'h00C9; #100;
A = 16'h0026; B = 16'h00CA; #100;
A = 16'h0026; B = 16'h00CB; #100;
A = 16'h0026; B = 16'h00CC; #100;
A = 16'h0026; B = 16'h00CD; #100;
A = 16'h0026; B = 16'h00CE; #100;
A = 16'h0026; B = 16'h00CF; #100;
A = 16'h0026; B = 16'h00D0; #100;
A = 16'h0026; B = 16'h00D1; #100;
A = 16'h0026; B = 16'h00D2; #100;
A = 16'h0026; B = 16'h00D3; #100;
A = 16'h0026; B = 16'h00D4; #100;
A = 16'h0026; B = 16'h00D5; #100;
A = 16'h0026; B = 16'h00D6; #100;
A = 16'h0026; B = 16'h00D7; #100;
A = 16'h0026; B = 16'h00D8; #100;
A = 16'h0026; B = 16'h00D9; #100;
A = 16'h0026; B = 16'h00DA; #100;
A = 16'h0026; B = 16'h00DB; #100;
A = 16'h0026; B = 16'h00DC; #100;
A = 16'h0026; B = 16'h00DD; #100;
A = 16'h0026; B = 16'h00DE; #100;
A = 16'h0026; B = 16'h00DF; #100;
A = 16'h0026; B = 16'h00E0; #100;
A = 16'h0026; B = 16'h00E1; #100;
A = 16'h0026; B = 16'h00E2; #100;
A = 16'h0026; B = 16'h00E3; #100;
A = 16'h0026; B = 16'h00E4; #100;
A = 16'h0026; B = 16'h00E5; #100;
A = 16'h0026; B = 16'h00E6; #100;
A = 16'h0026; B = 16'h00E7; #100;
A = 16'h0026; B = 16'h00E8; #100;
A = 16'h0026; B = 16'h00E9; #100;
A = 16'h0026; B = 16'h00EA; #100;
A = 16'h0026; B = 16'h00EB; #100;
A = 16'h0026; B = 16'h00EC; #100;
A = 16'h0026; B = 16'h00ED; #100;
A = 16'h0026; B = 16'h00EE; #100;
A = 16'h0026; B = 16'h00EF; #100;
A = 16'h0026; B = 16'h00F0; #100;
A = 16'h0026; B = 16'h00F1; #100;
A = 16'h0026; B = 16'h00F2; #100;
A = 16'h0026; B = 16'h00F3; #100;
A = 16'h0026; B = 16'h00F4; #100;
A = 16'h0026; B = 16'h00F5; #100;
A = 16'h0026; B = 16'h00F6; #100;
A = 16'h0026; B = 16'h00F7; #100;
A = 16'h0026; B = 16'h00F8; #100;
A = 16'h0026; B = 16'h00F9; #100;
A = 16'h0026; B = 16'h00FA; #100;
A = 16'h0026; B = 16'h00FB; #100;
A = 16'h0026; B = 16'h00FC; #100;
A = 16'h0026; B = 16'h00FD; #100;
A = 16'h0026; B = 16'h00FE; #100;
A = 16'h0026; B = 16'h00FF; #100;
A = 16'h0027; B = 16'h000; #100;
A = 16'h0027; B = 16'h001; #100;
A = 16'h0027; B = 16'h002; #100;
A = 16'h0027; B = 16'h003; #100;
A = 16'h0027; B = 16'h004; #100;
A = 16'h0027; B = 16'h005; #100;
A = 16'h0027; B = 16'h006; #100;
A = 16'h0027; B = 16'h007; #100;
A = 16'h0027; B = 16'h008; #100;
A = 16'h0027; B = 16'h009; #100;
A = 16'h0027; B = 16'h00A; #100;
A = 16'h0027; B = 16'h00B; #100;
A = 16'h0027; B = 16'h00C; #100;
A = 16'h0027; B = 16'h00D; #100;
A = 16'h0027; B = 16'h00E; #100;
A = 16'h0027; B = 16'h00F; #100;
A = 16'h0027; B = 16'h0010; #100;
A = 16'h0027; B = 16'h0011; #100;
A = 16'h0027; B = 16'h0012; #100;
A = 16'h0027; B = 16'h0013; #100;
A = 16'h0027; B = 16'h0014; #100;
A = 16'h0027; B = 16'h0015; #100;
A = 16'h0027; B = 16'h0016; #100;
A = 16'h0027; B = 16'h0017; #100;
A = 16'h0027; B = 16'h0018; #100;
A = 16'h0027; B = 16'h0019; #100;
A = 16'h0027; B = 16'h001A; #100;
A = 16'h0027; B = 16'h001B; #100;
A = 16'h0027; B = 16'h001C; #100;
A = 16'h0027; B = 16'h001D; #100;
A = 16'h0027; B = 16'h001E; #100;
A = 16'h0027; B = 16'h001F; #100;
A = 16'h0027; B = 16'h0020; #100;
A = 16'h0027; B = 16'h0021; #100;
A = 16'h0027; B = 16'h0022; #100;
A = 16'h0027; B = 16'h0023; #100;
A = 16'h0027; B = 16'h0024; #100;
A = 16'h0027; B = 16'h0025; #100;
A = 16'h0027; B = 16'h0026; #100;
A = 16'h0027; B = 16'h0027; #100;
A = 16'h0027; B = 16'h0028; #100;
A = 16'h0027; B = 16'h0029; #100;
A = 16'h0027; B = 16'h002A; #100;
A = 16'h0027; B = 16'h002B; #100;
A = 16'h0027; B = 16'h002C; #100;
A = 16'h0027; B = 16'h002D; #100;
A = 16'h0027; B = 16'h002E; #100;
A = 16'h0027; B = 16'h002F; #100;
A = 16'h0027; B = 16'h0030; #100;
A = 16'h0027; B = 16'h0031; #100;
A = 16'h0027; B = 16'h0032; #100;
A = 16'h0027; B = 16'h0033; #100;
A = 16'h0027; B = 16'h0034; #100;
A = 16'h0027; B = 16'h0035; #100;
A = 16'h0027; B = 16'h0036; #100;
A = 16'h0027; B = 16'h0037; #100;
A = 16'h0027; B = 16'h0038; #100;
A = 16'h0027; B = 16'h0039; #100;
A = 16'h0027; B = 16'h003A; #100;
A = 16'h0027; B = 16'h003B; #100;
A = 16'h0027; B = 16'h003C; #100;
A = 16'h0027; B = 16'h003D; #100;
A = 16'h0027; B = 16'h003E; #100;
A = 16'h0027; B = 16'h003F; #100;
A = 16'h0027; B = 16'h0040; #100;
A = 16'h0027; B = 16'h0041; #100;
A = 16'h0027; B = 16'h0042; #100;
A = 16'h0027; B = 16'h0043; #100;
A = 16'h0027; B = 16'h0044; #100;
A = 16'h0027; B = 16'h0045; #100;
A = 16'h0027; B = 16'h0046; #100;
A = 16'h0027; B = 16'h0047; #100;
A = 16'h0027; B = 16'h0048; #100;
A = 16'h0027; B = 16'h0049; #100;
A = 16'h0027; B = 16'h004A; #100;
A = 16'h0027; B = 16'h004B; #100;
A = 16'h0027; B = 16'h004C; #100;
A = 16'h0027; B = 16'h004D; #100;
A = 16'h0027; B = 16'h004E; #100;
A = 16'h0027; B = 16'h004F; #100;
A = 16'h0027; B = 16'h0050; #100;
A = 16'h0027; B = 16'h0051; #100;
A = 16'h0027; B = 16'h0052; #100;
A = 16'h0027; B = 16'h0053; #100;
A = 16'h0027; B = 16'h0054; #100;
A = 16'h0027; B = 16'h0055; #100;
A = 16'h0027; B = 16'h0056; #100;
A = 16'h0027; B = 16'h0057; #100;
A = 16'h0027; B = 16'h0058; #100;
A = 16'h0027; B = 16'h0059; #100;
A = 16'h0027; B = 16'h005A; #100;
A = 16'h0027; B = 16'h005B; #100;
A = 16'h0027; B = 16'h005C; #100;
A = 16'h0027; B = 16'h005D; #100;
A = 16'h0027; B = 16'h005E; #100;
A = 16'h0027; B = 16'h005F; #100;
A = 16'h0027; B = 16'h0060; #100;
A = 16'h0027; B = 16'h0061; #100;
A = 16'h0027; B = 16'h0062; #100;
A = 16'h0027; B = 16'h0063; #100;
A = 16'h0027; B = 16'h0064; #100;
A = 16'h0027; B = 16'h0065; #100;
A = 16'h0027; B = 16'h0066; #100;
A = 16'h0027; B = 16'h0067; #100;
A = 16'h0027; B = 16'h0068; #100;
A = 16'h0027; B = 16'h0069; #100;
A = 16'h0027; B = 16'h006A; #100;
A = 16'h0027; B = 16'h006B; #100;
A = 16'h0027; B = 16'h006C; #100;
A = 16'h0027; B = 16'h006D; #100;
A = 16'h0027; B = 16'h006E; #100;
A = 16'h0027; B = 16'h006F; #100;
A = 16'h0027; B = 16'h0070; #100;
A = 16'h0027; B = 16'h0071; #100;
A = 16'h0027; B = 16'h0072; #100;
A = 16'h0027; B = 16'h0073; #100;
A = 16'h0027; B = 16'h0074; #100;
A = 16'h0027; B = 16'h0075; #100;
A = 16'h0027; B = 16'h0076; #100;
A = 16'h0027; B = 16'h0077; #100;
A = 16'h0027; B = 16'h0078; #100;
A = 16'h0027; B = 16'h0079; #100;
A = 16'h0027; B = 16'h007A; #100;
A = 16'h0027; B = 16'h007B; #100;
A = 16'h0027; B = 16'h007C; #100;
A = 16'h0027; B = 16'h007D; #100;
A = 16'h0027; B = 16'h007E; #100;
A = 16'h0027; B = 16'h007F; #100;
A = 16'h0027; B = 16'h0080; #100;
A = 16'h0027; B = 16'h0081; #100;
A = 16'h0027; B = 16'h0082; #100;
A = 16'h0027; B = 16'h0083; #100;
A = 16'h0027; B = 16'h0084; #100;
A = 16'h0027; B = 16'h0085; #100;
A = 16'h0027; B = 16'h0086; #100;
A = 16'h0027; B = 16'h0087; #100;
A = 16'h0027; B = 16'h0088; #100;
A = 16'h0027; B = 16'h0089; #100;
A = 16'h0027; B = 16'h008A; #100;
A = 16'h0027; B = 16'h008B; #100;
A = 16'h0027; B = 16'h008C; #100;
A = 16'h0027; B = 16'h008D; #100;
A = 16'h0027; B = 16'h008E; #100;
A = 16'h0027; B = 16'h008F; #100;
A = 16'h0027; B = 16'h0090; #100;
A = 16'h0027; B = 16'h0091; #100;
A = 16'h0027; B = 16'h0092; #100;
A = 16'h0027; B = 16'h0093; #100;
A = 16'h0027; B = 16'h0094; #100;
A = 16'h0027; B = 16'h0095; #100;
A = 16'h0027; B = 16'h0096; #100;
A = 16'h0027; B = 16'h0097; #100;
A = 16'h0027; B = 16'h0098; #100;
A = 16'h0027; B = 16'h0099; #100;
A = 16'h0027; B = 16'h009A; #100;
A = 16'h0027; B = 16'h009B; #100;
A = 16'h0027; B = 16'h009C; #100;
A = 16'h0027; B = 16'h009D; #100;
A = 16'h0027; B = 16'h009E; #100;
A = 16'h0027; B = 16'h009F; #100;
A = 16'h0027; B = 16'h00A0; #100;
A = 16'h0027; B = 16'h00A1; #100;
A = 16'h0027; B = 16'h00A2; #100;
A = 16'h0027; B = 16'h00A3; #100;
A = 16'h0027; B = 16'h00A4; #100;
A = 16'h0027; B = 16'h00A5; #100;
A = 16'h0027; B = 16'h00A6; #100;
A = 16'h0027; B = 16'h00A7; #100;
A = 16'h0027; B = 16'h00A8; #100;
A = 16'h0027; B = 16'h00A9; #100;
A = 16'h0027; B = 16'h00AA; #100;
A = 16'h0027; B = 16'h00AB; #100;
A = 16'h0027; B = 16'h00AC; #100;
A = 16'h0027; B = 16'h00AD; #100;
A = 16'h0027; B = 16'h00AE; #100;
A = 16'h0027; B = 16'h00AF; #100;
A = 16'h0027; B = 16'h00B0; #100;
A = 16'h0027; B = 16'h00B1; #100;
A = 16'h0027; B = 16'h00B2; #100;
A = 16'h0027; B = 16'h00B3; #100;
A = 16'h0027; B = 16'h00B4; #100;
A = 16'h0027; B = 16'h00B5; #100;
A = 16'h0027; B = 16'h00B6; #100;
A = 16'h0027; B = 16'h00B7; #100;
A = 16'h0027; B = 16'h00B8; #100;
A = 16'h0027; B = 16'h00B9; #100;
A = 16'h0027; B = 16'h00BA; #100;
A = 16'h0027; B = 16'h00BB; #100;
A = 16'h0027; B = 16'h00BC; #100;
A = 16'h0027; B = 16'h00BD; #100;
A = 16'h0027; B = 16'h00BE; #100;
A = 16'h0027; B = 16'h00BF; #100;
A = 16'h0027; B = 16'h00C0; #100;
A = 16'h0027; B = 16'h00C1; #100;
A = 16'h0027; B = 16'h00C2; #100;
A = 16'h0027; B = 16'h00C3; #100;
A = 16'h0027; B = 16'h00C4; #100;
A = 16'h0027; B = 16'h00C5; #100;
A = 16'h0027; B = 16'h00C6; #100;
A = 16'h0027; B = 16'h00C7; #100;
A = 16'h0027; B = 16'h00C8; #100;
A = 16'h0027; B = 16'h00C9; #100;
A = 16'h0027; B = 16'h00CA; #100;
A = 16'h0027; B = 16'h00CB; #100;
A = 16'h0027; B = 16'h00CC; #100;
A = 16'h0027; B = 16'h00CD; #100;
A = 16'h0027; B = 16'h00CE; #100;
A = 16'h0027; B = 16'h00CF; #100;
A = 16'h0027; B = 16'h00D0; #100;
A = 16'h0027; B = 16'h00D1; #100;
A = 16'h0027; B = 16'h00D2; #100;
A = 16'h0027; B = 16'h00D3; #100;
A = 16'h0027; B = 16'h00D4; #100;
A = 16'h0027; B = 16'h00D5; #100;
A = 16'h0027; B = 16'h00D6; #100;
A = 16'h0027; B = 16'h00D7; #100;
A = 16'h0027; B = 16'h00D8; #100;
A = 16'h0027; B = 16'h00D9; #100;
A = 16'h0027; B = 16'h00DA; #100;
A = 16'h0027; B = 16'h00DB; #100;
A = 16'h0027; B = 16'h00DC; #100;
A = 16'h0027; B = 16'h00DD; #100;
A = 16'h0027; B = 16'h00DE; #100;
A = 16'h0027; B = 16'h00DF; #100;
A = 16'h0027; B = 16'h00E0; #100;
A = 16'h0027; B = 16'h00E1; #100;
A = 16'h0027; B = 16'h00E2; #100;
A = 16'h0027; B = 16'h00E3; #100;
A = 16'h0027; B = 16'h00E4; #100;
A = 16'h0027; B = 16'h00E5; #100;
A = 16'h0027; B = 16'h00E6; #100;
A = 16'h0027; B = 16'h00E7; #100;
A = 16'h0027; B = 16'h00E8; #100;
A = 16'h0027; B = 16'h00E9; #100;
A = 16'h0027; B = 16'h00EA; #100;
A = 16'h0027; B = 16'h00EB; #100;
A = 16'h0027; B = 16'h00EC; #100;
A = 16'h0027; B = 16'h00ED; #100;
A = 16'h0027; B = 16'h00EE; #100;
A = 16'h0027; B = 16'h00EF; #100;
A = 16'h0027; B = 16'h00F0; #100;
A = 16'h0027; B = 16'h00F1; #100;
A = 16'h0027; B = 16'h00F2; #100;
A = 16'h0027; B = 16'h00F3; #100;
A = 16'h0027; B = 16'h00F4; #100;
A = 16'h0027; B = 16'h00F5; #100;
A = 16'h0027; B = 16'h00F6; #100;
A = 16'h0027; B = 16'h00F7; #100;
A = 16'h0027; B = 16'h00F8; #100;
A = 16'h0027; B = 16'h00F9; #100;
A = 16'h0027; B = 16'h00FA; #100;
A = 16'h0027; B = 16'h00FB; #100;
A = 16'h0027; B = 16'h00FC; #100;
A = 16'h0027; B = 16'h00FD; #100;
A = 16'h0027; B = 16'h00FE; #100;
A = 16'h0027; B = 16'h00FF; #100;
A = 16'h0028; B = 16'h000; #100;
A = 16'h0028; B = 16'h001; #100;
A = 16'h0028; B = 16'h002; #100;
A = 16'h0028; B = 16'h003; #100;
A = 16'h0028; B = 16'h004; #100;
A = 16'h0028; B = 16'h005; #100;
A = 16'h0028; B = 16'h006; #100;
A = 16'h0028; B = 16'h007; #100;
A = 16'h0028; B = 16'h008; #100;
A = 16'h0028; B = 16'h009; #100;
A = 16'h0028; B = 16'h00A; #100;
A = 16'h0028; B = 16'h00B; #100;
A = 16'h0028; B = 16'h00C; #100;
A = 16'h0028; B = 16'h00D; #100;
A = 16'h0028; B = 16'h00E; #100;
A = 16'h0028; B = 16'h00F; #100;
A = 16'h0028; B = 16'h0010; #100;
A = 16'h0028; B = 16'h0011; #100;
A = 16'h0028; B = 16'h0012; #100;
A = 16'h0028; B = 16'h0013; #100;
A = 16'h0028; B = 16'h0014; #100;
A = 16'h0028; B = 16'h0015; #100;
A = 16'h0028; B = 16'h0016; #100;
A = 16'h0028; B = 16'h0017; #100;
A = 16'h0028; B = 16'h0018; #100;
A = 16'h0028; B = 16'h0019; #100;
A = 16'h0028; B = 16'h001A; #100;
A = 16'h0028; B = 16'h001B; #100;
A = 16'h0028; B = 16'h001C; #100;
A = 16'h0028; B = 16'h001D; #100;
A = 16'h0028; B = 16'h001E; #100;
A = 16'h0028; B = 16'h001F; #100;
A = 16'h0028; B = 16'h0020; #100;
A = 16'h0028; B = 16'h0021; #100;
A = 16'h0028; B = 16'h0022; #100;
A = 16'h0028; B = 16'h0023; #100;
A = 16'h0028; B = 16'h0024; #100;
A = 16'h0028; B = 16'h0025; #100;
A = 16'h0028; B = 16'h0026; #100;
A = 16'h0028; B = 16'h0027; #100;
A = 16'h0028; B = 16'h0028; #100;
A = 16'h0028; B = 16'h0029; #100;
A = 16'h0028; B = 16'h002A; #100;
A = 16'h0028; B = 16'h002B; #100;
A = 16'h0028; B = 16'h002C; #100;
A = 16'h0028; B = 16'h002D; #100;
A = 16'h0028; B = 16'h002E; #100;
A = 16'h0028; B = 16'h002F; #100;
A = 16'h0028; B = 16'h0030; #100;
A = 16'h0028; B = 16'h0031; #100;
A = 16'h0028; B = 16'h0032; #100;
A = 16'h0028; B = 16'h0033; #100;
A = 16'h0028; B = 16'h0034; #100;
A = 16'h0028; B = 16'h0035; #100;
A = 16'h0028; B = 16'h0036; #100;
A = 16'h0028; B = 16'h0037; #100;
A = 16'h0028; B = 16'h0038; #100;
A = 16'h0028; B = 16'h0039; #100;
A = 16'h0028; B = 16'h003A; #100;
A = 16'h0028; B = 16'h003B; #100;
A = 16'h0028; B = 16'h003C; #100;
A = 16'h0028; B = 16'h003D; #100;
A = 16'h0028; B = 16'h003E; #100;
A = 16'h0028; B = 16'h003F; #100;
A = 16'h0028; B = 16'h0040; #100;
A = 16'h0028; B = 16'h0041; #100;
A = 16'h0028; B = 16'h0042; #100;
A = 16'h0028; B = 16'h0043; #100;
A = 16'h0028; B = 16'h0044; #100;
A = 16'h0028; B = 16'h0045; #100;
A = 16'h0028; B = 16'h0046; #100;
A = 16'h0028; B = 16'h0047; #100;
A = 16'h0028; B = 16'h0048; #100;
A = 16'h0028; B = 16'h0049; #100;
A = 16'h0028; B = 16'h004A; #100;
A = 16'h0028; B = 16'h004B; #100;
A = 16'h0028; B = 16'h004C; #100;
A = 16'h0028; B = 16'h004D; #100;
A = 16'h0028; B = 16'h004E; #100;
A = 16'h0028; B = 16'h004F; #100;
A = 16'h0028; B = 16'h0050; #100;
A = 16'h0028; B = 16'h0051; #100;
A = 16'h0028; B = 16'h0052; #100;
A = 16'h0028; B = 16'h0053; #100;
A = 16'h0028; B = 16'h0054; #100;
A = 16'h0028; B = 16'h0055; #100;
A = 16'h0028; B = 16'h0056; #100;
A = 16'h0028; B = 16'h0057; #100;
A = 16'h0028; B = 16'h0058; #100;
A = 16'h0028; B = 16'h0059; #100;
A = 16'h0028; B = 16'h005A; #100;
A = 16'h0028; B = 16'h005B; #100;
A = 16'h0028; B = 16'h005C; #100;
A = 16'h0028; B = 16'h005D; #100;
A = 16'h0028; B = 16'h005E; #100;
A = 16'h0028; B = 16'h005F; #100;
A = 16'h0028; B = 16'h0060; #100;
A = 16'h0028; B = 16'h0061; #100;
A = 16'h0028; B = 16'h0062; #100;
A = 16'h0028; B = 16'h0063; #100;
A = 16'h0028; B = 16'h0064; #100;
A = 16'h0028; B = 16'h0065; #100;
A = 16'h0028; B = 16'h0066; #100;
A = 16'h0028; B = 16'h0067; #100;
A = 16'h0028; B = 16'h0068; #100;
A = 16'h0028; B = 16'h0069; #100;
A = 16'h0028; B = 16'h006A; #100;
A = 16'h0028; B = 16'h006B; #100;
A = 16'h0028; B = 16'h006C; #100;
A = 16'h0028; B = 16'h006D; #100;
A = 16'h0028; B = 16'h006E; #100;
A = 16'h0028; B = 16'h006F; #100;
A = 16'h0028; B = 16'h0070; #100;
A = 16'h0028; B = 16'h0071; #100;
A = 16'h0028; B = 16'h0072; #100;
A = 16'h0028; B = 16'h0073; #100;
A = 16'h0028; B = 16'h0074; #100;
A = 16'h0028; B = 16'h0075; #100;
A = 16'h0028; B = 16'h0076; #100;
A = 16'h0028; B = 16'h0077; #100;
A = 16'h0028; B = 16'h0078; #100;
A = 16'h0028; B = 16'h0079; #100;
A = 16'h0028; B = 16'h007A; #100;
A = 16'h0028; B = 16'h007B; #100;
A = 16'h0028; B = 16'h007C; #100;
A = 16'h0028; B = 16'h007D; #100;
A = 16'h0028; B = 16'h007E; #100;
A = 16'h0028; B = 16'h007F; #100;
A = 16'h0028; B = 16'h0080; #100;
A = 16'h0028; B = 16'h0081; #100;
A = 16'h0028; B = 16'h0082; #100;
A = 16'h0028; B = 16'h0083; #100;
A = 16'h0028; B = 16'h0084; #100;
A = 16'h0028; B = 16'h0085; #100;
A = 16'h0028; B = 16'h0086; #100;
A = 16'h0028; B = 16'h0087; #100;
A = 16'h0028; B = 16'h0088; #100;
A = 16'h0028; B = 16'h0089; #100;
A = 16'h0028; B = 16'h008A; #100;
A = 16'h0028; B = 16'h008B; #100;
A = 16'h0028; B = 16'h008C; #100;
A = 16'h0028; B = 16'h008D; #100;
A = 16'h0028; B = 16'h008E; #100;
A = 16'h0028; B = 16'h008F; #100;
A = 16'h0028; B = 16'h0090; #100;
A = 16'h0028; B = 16'h0091; #100;
A = 16'h0028; B = 16'h0092; #100;
A = 16'h0028; B = 16'h0093; #100;
A = 16'h0028; B = 16'h0094; #100;
A = 16'h0028; B = 16'h0095; #100;
A = 16'h0028; B = 16'h0096; #100;
A = 16'h0028; B = 16'h0097; #100;
A = 16'h0028; B = 16'h0098; #100;
A = 16'h0028; B = 16'h0099; #100;
A = 16'h0028; B = 16'h009A; #100;
A = 16'h0028; B = 16'h009B; #100;
A = 16'h0028; B = 16'h009C; #100;
A = 16'h0028; B = 16'h009D; #100;
A = 16'h0028; B = 16'h009E; #100;
A = 16'h0028; B = 16'h009F; #100;
A = 16'h0028; B = 16'h00A0; #100;
A = 16'h0028; B = 16'h00A1; #100;
A = 16'h0028; B = 16'h00A2; #100;
A = 16'h0028; B = 16'h00A3; #100;
A = 16'h0028; B = 16'h00A4; #100;
A = 16'h0028; B = 16'h00A5; #100;
A = 16'h0028; B = 16'h00A6; #100;
A = 16'h0028; B = 16'h00A7; #100;
A = 16'h0028; B = 16'h00A8; #100;
A = 16'h0028; B = 16'h00A9; #100;
A = 16'h0028; B = 16'h00AA; #100;
A = 16'h0028; B = 16'h00AB; #100;
A = 16'h0028; B = 16'h00AC; #100;
A = 16'h0028; B = 16'h00AD; #100;
A = 16'h0028; B = 16'h00AE; #100;
A = 16'h0028; B = 16'h00AF; #100;
A = 16'h0028; B = 16'h00B0; #100;
A = 16'h0028; B = 16'h00B1; #100;
A = 16'h0028; B = 16'h00B2; #100;
A = 16'h0028; B = 16'h00B3; #100;
A = 16'h0028; B = 16'h00B4; #100;
A = 16'h0028; B = 16'h00B5; #100;
A = 16'h0028; B = 16'h00B6; #100;
A = 16'h0028; B = 16'h00B7; #100;
A = 16'h0028; B = 16'h00B8; #100;
A = 16'h0028; B = 16'h00B9; #100;
A = 16'h0028; B = 16'h00BA; #100;
A = 16'h0028; B = 16'h00BB; #100;
A = 16'h0028; B = 16'h00BC; #100;
A = 16'h0028; B = 16'h00BD; #100;
A = 16'h0028; B = 16'h00BE; #100;
A = 16'h0028; B = 16'h00BF; #100;
A = 16'h0028; B = 16'h00C0; #100;
A = 16'h0028; B = 16'h00C1; #100;
A = 16'h0028; B = 16'h00C2; #100;
A = 16'h0028; B = 16'h00C3; #100;
A = 16'h0028; B = 16'h00C4; #100;
A = 16'h0028; B = 16'h00C5; #100;
A = 16'h0028; B = 16'h00C6; #100;
A = 16'h0028; B = 16'h00C7; #100;
A = 16'h0028; B = 16'h00C8; #100;
A = 16'h0028; B = 16'h00C9; #100;
A = 16'h0028; B = 16'h00CA; #100;
A = 16'h0028; B = 16'h00CB; #100;
A = 16'h0028; B = 16'h00CC; #100;
A = 16'h0028; B = 16'h00CD; #100;
A = 16'h0028; B = 16'h00CE; #100;
A = 16'h0028; B = 16'h00CF; #100;
A = 16'h0028; B = 16'h00D0; #100;
A = 16'h0028; B = 16'h00D1; #100;
A = 16'h0028; B = 16'h00D2; #100;
A = 16'h0028; B = 16'h00D3; #100;
A = 16'h0028; B = 16'h00D4; #100;
A = 16'h0028; B = 16'h00D5; #100;
A = 16'h0028; B = 16'h00D6; #100;
A = 16'h0028; B = 16'h00D7; #100;
A = 16'h0028; B = 16'h00D8; #100;
A = 16'h0028; B = 16'h00D9; #100;
A = 16'h0028; B = 16'h00DA; #100;
A = 16'h0028; B = 16'h00DB; #100;
A = 16'h0028; B = 16'h00DC; #100;
A = 16'h0028; B = 16'h00DD; #100;
A = 16'h0028; B = 16'h00DE; #100;
A = 16'h0028; B = 16'h00DF; #100;
A = 16'h0028; B = 16'h00E0; #100;
A = 16'h0028; B = 16'h00E1; #100;
A = 16'h0028; B = 16'h00E2; #100;
A = 16'h0028; B = 16'h00E3; #100;
A = 16'h0028; B = 16'h00E4; #100;
A = 16'h0028; B = 16'h00E5; #100;
A = 16'h0028; B = 16'h00E6; #100;
A = 16'h0028; B = 16'h00E7; #100;
A = 16'h0028; B = 16'h00E8; #100;
A = 16'h0028; B = 16'h00E9; #100;
A = 16'h0028; B = 16'h00EA; #100;
A = 16'h0028; B = 16'h00EB; #100;
A = 16'h0028; B = 16'h00EC; #100;
A = 16'h0028; B = 16'h00ED; #100;
A = 16'h0028; B = 16'h00EE; #100;
A = 16'h0028; B = 16'h00EF; #100;
A = 16'h0028; B = 16'h00F0; #100;
A = 16'h0028; B = 16'h00F1; #100;
A = 16'h0028; B = 16'h00F2; #100;
A = 16'h0028; B = 16'h00F3; #100;
A = 16'h0028; B = 16'h00F4; #100;
A = 16'h0028; B = 16'h00F5; #100;
A = 16'h0028; B = 16'h00F6; #100;
A = 16'h0028; B = 16'h00F7; #100;
A = 16'h0028; B = 16'h00F8; #100;
A = 16'h0028; B = 16'h00F9; #100;
A = 16'h0028; B = 16'h00FA; #100;
A = 16'h0028; B = 16'h00FB; #100;
A = 16'h0028; B = 16'h00FC; #100;
A = 16'h0028; B = 16'h00FD; #100;
A = 16'h0028; B = 16'h00FE; #100;
A = 16'h0028; B = 16'h00FF; #100;
A = 16'h0029; B = 16'h000; #100;
A = 16'h0029; B = 16'h001; #100;
A = 16'h0029; B = 16'h002; #100;
A = 16'h0029; B = 16'h003; #100;
A = 16'h0029; B = 16'h004; #100;
A = 16'h0029; B = 16'h005; #100;
A = 16'h0029; B = 16'h006; #100;
A = 16'h0029; B = 16'h007; #100;
A = 16'h0029; B = 16'h008; #100;
A = 16'h0029; B = 16'h009; #100;
A = 16'h0029; B = 16'h00A; #100;
A = 16'h0029; B = 16'h00B; #100;
A = 16'h0029; B = 16'h00C; #100;
A = 16'h0029; B = 16'h00D; #100;
A = 16'h0029; B = 16'h00E; #100;
A = 16'h0029; B = 16'h00F; #100;
A = 16'h0029; B = 16'h0010; #100;
A = 16'h0029; B = 16'h0011; #100;
A = 16'h0029; B = 16'h0012; #100;
A = 16'h0029; B = 16'h0013; #100;
A = 16'h0029; B = 16'h0014; #100;
A = 16'h0029; B = 16'h0015; #100;
A = 16'h0029; B = 16'h0016; #100;
A = 16'h0029; B = 16'h0017; #100;
A = 16'h0029; B = 16'h0018; #100;
A = 16'h0029; B = 16'h0019; #100;
A = 16'h0029; B = 16'h001A; #100;
A = 16'h0029; B = 16'h001B; #100;
A = 16'h0029; B = 16'h001C; #100;
A = 16'h0029; B = 16'h001D; #100;
A = 16'h0029; B = 16'h001E; #100;
A = 16'h0029; B = 16'h001F; #100;
A = 16'h0029; B = 16'h0020; #100;
A = 16'h0029; B = 16'h0021; #100;
A = 16'h0029; B = 16'h0022; #100;
A = 16'h0029; B = 16'h0023; #100;
A = 16'h0029; B = 16'h0024; #100;
A = 16'h0029; B = 16'h0025; #100;
A = 16'h0029; B = 16'h0026; #100;
A = 16'h0029; B = 16'h0027; #100;
A = 16'h0029; B = 16'h0028; #100;
A = 16'h0029; B = 16'h0029; #100;
A = 16'h0029; B = 16'h002A; #100;
A = 16'h0029; B = 16'h002B; #100;
A = 16'h0029; B = 16'h002C; #100;
A = 16'h0029; B = 16'h002D; #100;
A = 16'h0029; B = 16'h002E; #100;
A = 16'h0029; B = 16'h002F; #100;
A = 16'h0029; B = 16'h0030; #100;
A = 16'h0029; B = 16'h0031; #100;
A = 16'h0029; B = 16'h0032; #100;
A = 16'h0029; B = 16'h0033; #100;
A = 16'h0029; B = 16'h0034; #100;
A = 16'h0029; B = 16'h0035; #100;
A = 16'h0029; B = 16'h0036; #100;
A = 16'h0029; B = 16'h0037; #100;
A = 16'h0029; B = 16'h0038; #100;
A = 16'h0029; B = 16'h0039; #100;
A = 16'h0029; B = 16'h003A; #100;
A = 16'h0029; B = 16'h003B; #100;
A = 16'h0029; B = 16'h003C; #100;
A = 16'h0029; B = 16'h003D; #100;
A = 16'h0029; B = 16'h003E; #100;
A = 16'h0029; B = 16'h003F; #100;
A = 16'h0029; B = 16'h0040; #100;
A = 16'h0029; B = 16'h0041; #100;
A = 16'h0029; B = 16'h0042; #100;
A = 16'h0029; B = 16'h0043; #100;
A = 16'h0029; B = 16'h0044; #100;
A = 16'h0029; B = 16'h0045; #100;
A = 16'h0029; B = 16'h0046; #100;
A = 16'h0029; B = 16'h0047; #100;
A = 16'h0029; B = 16'h0048; #100;
A = 16'h0029; B = 16'h0049; #100;
A = 16'h0029; B = 16'h004A; #100;
A = 16'h0029; B = 16'h004B; #100;
A = 16'h0029; B = 16'h004C; #100;
A = 16'h0029; B = 16'h004D; #100;
A = 16'h0029; B = 16'h004E; #100;
A = 16'h0029; B = 16'h004F; #100;
A = 16'h0029; B = 16'h0050; #100;
A = 16'h0029; B = 16'h0051; #100;
A = 16'h0029; B = 16'h0052; #100;
A = 16'h0029; B = 16'h0053; #100;
A = 16'h0029; B = 16'h0054; #100;
A = 16'h0029; B = 16'h0055; #100;
A = 16'h0029; B = 16'h0056; #100;
A = 16'h0029; B = 16'h0057; #100;
A = 16'h0029; B = 16'h0058; #100;
A = 16'h0029; B = 16'h0059; #100;
A = 16'h0029; B = 16'h005A; #100;
A = 16'h0029; B = 16'h005B; #100;
A = 16'h0029; B = 16'h005C; #100;
A = 16'h0029; B = 16'h005D; #100;
A = 16'h0029; B = 16'h005E; #100;
A = 16'h0029; B = 16'h005F; #100;
A = 16'h0029; B = 16'h0060; #100;
A = 16'h0029; B = 16'h0061; #100;
A = 16'h0029; B = 16'h0062; #100;
A = 16'h0029; B = 16'h0063; #100;
A = 16'h0029; B = 16'h0064; #100;
A = 16'h0029; B = 16'h0065; #100;
A = 16'h0029; B = 16'h0066; #100;
A = 16'h0029; B = 16'h0067; #100;
A = 16'h0029; B = 16'h0068; #100;
A = 16'h0029; B = 16'h0069; #100;
A = 16'h0029; B = 16'h006A; #100;
A = 16'h0029; B = 16'h006B; #100;
A = 16'h0029; B = 16'h006C; #100;
A = 16'h0029; B = 16'h006D; #100;
A = 16'h0029; B = 16'h006E; #100;
A = 16'h0029; B = 16'h006F; #100;
A = 16'h0029; B = 16'h0070; #100;
A = 16'h0029; B = 16'h0071; #100;
A = 16'h0029; B = 16'h0072; #100;
A = 16'h0029; B = 16'h0073; #100;
A = 16'h0029; B = 16'h0074; #100;
A = 16'h0029; B = 16'h0075; #100;
A = 16'h0029; B = 16'h0076; #100;
A = 16'h0029; B = 16'h0077; #100;
A = 16'h0029; B = 16'h0078; #100;
A = 16'h0029; B = 16'h0079; #100;
A = 16'h0029; B = 16'h007A; #100;
A = 16'h0029; B = 16'h007B; #100;
A = 16'h0029; B = 16'h007C; #100;
A = 16'h0029; B = 16'h007D; #100;
A = 16'h0029; B = 16'h007E; #100;
A = 16'h0029; B = 16'h007F; #100;
A = 16'h0029; B = 16'h0080; #100;
A = 16'h0029; B = 16'h0081; #100;
A = 16'h0029; B = 16'h0082; #100;
A = 16'h0029; B = 16'h0083; #100;
A = 16'h0029; B = 16'h0084; #100;
A = 16'h0029; B = 16'h0085; #100;
A = 16'h0029; B = 16'h0086; #100;
A = 16'h0029; B = 16'h0087; #100;
A = 16'h0029; B = 16'h0088; #100;
A = 16'h0029; B = 16'h0089; #100;
A = 16'h0029; B = 16'h008A; #100;
A = 16'h0029; B = 16'h008B; #100;
A = 16'h0029; B = 16'h008C; #100;
A = 16'h0029; B = 16'h008D; #100;
A = 16'h0029; B = 16'h008E; #100;
A = 16'h0029; B = 16'h008F; #100;
A = 16'h0029; B = 16'h0090; #100;
A = 16'h0029; B = 16'h0091; #100;
A = 16'h0029; B = 16'h0092; #100;
A = 16'h0029; B = 16'h0093; #100;
A = 16'h0029; B = 16'h0094; #100;
A = 16'h0029; B = 16'h0095; #100;
A = 16'h0029; B = 16'h0096; #100;
A = 16'h0029; B = 16'h0097; #100;
A = 16'h0029; B = 16'h0098; #100;
A = 16'h0029; B = 16'h0099; #100;
A = 16'h0029; B = 16'h009A; #100;
A = 16'h0029; B = 16'h009B; #100;
A = 16'h0029; B = 16'h009C; #100;
A = 16'h0029; B = 16'h009D; #100;
A = 16'h0029; B = 16'h009E; #100;
A = 16'h0029; B = 16'h009F; #100;
A = 16'h0029; B = 16'h00A0; #100;
A = 16'h0029; B = 16'h00A1; #100;
A = 16'h0029; B = 16'h00A2; #100;
A = 16'h0029; B = 16'h00A3; #100;
A = 16'h0029; B = 16'h00A4; #100;
A = 16'h0029; B = 16'h00A5; #100;
A = 16'h0029; B = 16'h00A6; #100;
A = 16'h0029; B = 16'h00A7; #100;
A = 16'h0029; B = 16'h00A8; #100;
A = 16'h0029; B = 16'h00A9; #100;
A = 16'h0029; B = 16'h00AA; #100;
A = 16'h0029; B = 16'h00AB; #100;
A = 16'h0029; B = 16'h00AC; #100;
A = 16'h0029; B = 16'h00AD; #100;
A = 16'h0029; B = 16'h00AE; #100;
A = 16'h0029; B = 16'h00AF; #100;
A = 16'h0029; B = 16'h00B0; #100;
A = 16'h0029; B = 16'h00B1; #100;
A = 16'h0029; B = 16'h00B2; #100;
A = 16'h0029; B = 16'h00B3; #100;
A = 16'h0029; B = 16'h00B4; #100;
A = 16'h0029; B = 16'h00B5; #100;
A = 16'h0029; B = 16'h00B6; #100;
A = 16'h0029; B = 16'h00B7; #100;
A = 16'h0029; B = 16'h00B8; #100;
A = 16'h0029; B = 16'h00B9; #100;
A = 16'h0029; B = 16'h00BA; #100;
A = 16'h0029; B = 16'h00BB; #100;
A = 16'h0029; B = 16'h00BC; #100;
A = 16'h0029; B = 16'h00BD; #100;
A = 16'h0029; B = 16'h00BE; #100;
A = 16'h0029; B = 16'h00BF; #100;
A = 16'h0029; B = 16'h00C0; #100;
A = 16'h0029; B = 16'h00C1; #100;
A = 16'h0029; B = 16'h00C2; #100;
A = 16'h0029; B = 16'h00C3; #100;
A = 16'h0029; B = 16'h00C4; #100;
A = 16'h0029; B = 16'h00C5; #100;
A = 16'h0029; B = 16'h00C6; #100;
A = 16'h0029; B = 16'h00C7; #100;
A = 16'h0029; B = 16'h00C8; #100;
A = 16'h0029; B = 16'h00C9; #100;
A = 16'h0029; B = 16'h00CA; #100;
A = 16'h0029; B = 16'h00CB; #100;
A = 16'h0029; B = 16'h00CC; #100;
A = 16'h0029; B = 16'h00CD; #100;
A = 16'h0029; B = 16'h00CE; #100;
A = 16'h0029; B = 16'h00CF; #100;
A = 16'h0029; B = 16'h00D0; #100;
A = 16'h0029; B = 16'h00D1; #100;
A = 16'h0029; B = 16'h00D2; #100;
A = 16'h0029; B = 16'h00D3; #100;
A = 16'h0029; B = 16'h00D4; #100;
A = 16'h0029; B = 16'h00D5; #100;
A = 16'h0029; B = 16'h00D6; #100;
A = 16'h0029; B = 16'h00D7; #100;
A = 16'h0029; B = 16'h00D8; #100;
A = 16'h0029; B = 16'h00D9; #100;
A = 16'h0029; B = 16'h00DA; #100;
A = 16'h0029; B = 16'h00DB; #100;
A = 16'h0029; B = 16'h00DC; #100;
A = 16'h0029; B = 16'h00DD; #100;
A = 16'h0029; B = 16'h00DE; #100;
A = 16'h0029; B = 16'h00DF; #100;
A = 16'h0029; B = 16'h00E0; #100;
A = 16'h0029; B = 16'h00E1; #100;
A = 16'h0029; B = 16'h00E2; #100;
A = 16'h0029; B = 16'h00E3; #100;
A = 16'h0029; B = 16'h00E4; #100;
A = 16'h0029; B = 16'h00E5; #100;
A = 16'h0029; B = 16'h00E6; #100;
A = 16'h0029; B = 16'h00E7; #100;
A = 16'h0029; B = 16'h00E8; #100;
A = 16'h0029; B = 16'h00E9; #100;
A = 16'h0029; B = 16'h00EA; #100;
A = 16'h0029; B = 16'h00EB; #100;
A = 16'h0029; B = 16'h00EC; #100;
A = 16'h0029; B = 16'h00ED; #100;
A = 16'h0029; B = 16'h00EE; #100;
A = 16'h0029; B = 16'h00EF; #100;
A = 16'h0029; B = 16'h00F0; #100;
A = 16'h0029; B = 16'h00F1; #100;
A = 16'h0029; B = 16'h00F2; #100;
A = 16'h0029; B = 16'h00F3; #100;
A = 16'h0029; B = 16'h00F4; #100;
A = 16'h0029; B = 16'h00F5; #100;
A = 16'h0029; B = 16'h00F6; #100;
A = 16'h0029; B = 16'h00F7; #100;
A = 16'h0029; B = 16'h00F8; #100;
A = 16'h0029; B = 16'h00F9; #100;
A = 16'h0029; B = 16'h00FA; #100;
A = 16'h0029; B = 16'h00FB; #100;
A = 16'h0029; B = 16'h00FC; #100;
A = 16'h0029; B = 16'h00FD; #100;
A = 16'h0029; B = 16'h00FE; #100;
A = 16'h0029; B = 16'h00FF; #100;
A = 16'h002A; B = 16'h000; #100;
A = 16'h002A; B = 16'h001; #100;
A = 16'h002A; B = 16'h002; #100;
A = 16'h002A; B = 16'h003; #100;
A = 16'h002A; B = 16'h004; #100;
A = 16'h002A; B = 16'h005; #100;
A = 16'h002A; B = 16'h006; #100;
A = 16'h002A; B = 16'h007; #100;
A = 16'h002A; B = 16'h008; #100;
A = 16'h002A; B = 16'h009; #100;
A = 16'h002A; B = 16'h00A; #100;
A = 16'h002A; B = 16'h00B; #100;
A = 16'h002A; B = 16'h00C; #100;
A = 16'h002A; B = 16'h00D; #100;
A = 16'h002A; B = 16'h00E; #100;
A = 16'h002A; B = 16'h00F; #100;
A = 16'h002A; B = 16'h0010; #100;
A = 16'h002A; B = 16'h0011; #100;
A = 16'h002A; B = 16'h0012; #100;
A = 16'h002A; B = 16'h0013; #100;
A = 16'h002A; B = 16'h0014; #100;
A = 16'h002A; B = 16'h0015; #100;
A = 16'h002A; B = 16'h0016; #100;
A = 16'h002A; B = 16'h0017; #100;
A = 16'h002A; B = 16'h0018; #100;
A = 16'h002A; B = 16'h0019; #100;
A = 16'h002A; B = 16'h001A; #100;
A = 16'h002A; B = 16'h001B; #100;
A = 16'h002A; B = 16'h001C; #100;
A = 16'h002A; B = 16'h001D; #100;
A = 16'h002A; B = 16'h001E; #100;
A = 16'h002A; B = 16'h001F; #100;
A = 16'h002A; B = 16'h0020; #100;
A = 16'h002A; B = 16'h0021; #100;
A = 16'h002A; B = 16'h0022; #100;
A = 16'h002A; B = 16'h0023; #100;
A = 16'h002A; B = 16'h0024; #100;
A = 16'h002A; B = 16'h0025; #100;
A = 16'h002A; B = 16'h0026; #100;
A = 16'h002A; B = 16'h0027; #100;
A = 16'h002A; B = 16'h0028; #100;
A = 16'h002A; B = 16'h0029; #100;
A = 16'h002A; B = 16'h002A; #100;
A = 16'h002A; B = 16'h002B; #100;
A = 16'h002A; B = 16'h002C; #100;
A = 16'h002A; B = 16'h002D; #100;
A = 16'h002A; B = 16'h002E; #100;
A = 16'h002A; B = 16'h002F; #100;
A = 16'h002A; B = 16'h0030; #100;
A = 16'h002A; B = 16'h0031; #100;
A = 16'h002A; B = 16'h0032; #100;
A = 16'h002A; B = 16'h0033; #100;
A = 16'h002A; B = 16'h0034; #100;
A = 16'h002A; B = 16'h0035; #100;
A = 16'h002A; B = 16'h0036; #100;
A = 16'h002A; B = 16'h0037; #100;
A = 16'h002A; B = 16'h0038; #100;
A = 16'h002A; B = 16'h0039; #100;
A = 16'h002A; B = 16'h003A; #100;
A = 16'h002A; B = 16'h003B; #100;
A = 16'h002A; B = 16'h003C; #100;
A = 16'h002A; B = 16'h003D; #100;
A = 16'h002A; B = 16'h003E; #100;
A = 16'h002A; B = 16'h003F; #100;
A = 16'h002A; B = 16'h0040; #100;
A = 16'h002A; B = 16'h0041; #100;
A = 16'h002A; B = 16'h0042; #100;
A = 16'h002A; B = 16'h0043; #100;
A = 16'h002A; B = 16'h0044; #100;
A = 16'h002A; B = 16'h0045; #100;
A = 16'h002A; B = 16'h0046; #100;
A = 16'h002A; B = 16'h0047; #100;
A = 16'h002A; B = 16'h0048; #100;
A = 16'h002A; B = 16'h0049; #100;
A = 16'h002A; B = 16'h004A; #100;
A = 16'h002A; B = 16'h004B; #100;
A = 16'h002A; B = 16'h004C; #100;
A = 16'h002A; B = 16'h004D; #100;
A = 16'h002A; B = 16'h004E; #100;
A = 16'h002A; B = 16'h004F; #100;
A = 16'h002A; B = 16'h0050; #100;
A = 16'h002A; B = 16'h0051; #100;
A = 16'h002A; B = 16'h0052; #100;
A = 16'h002A; B = 16'h0053; #100;
A = 16'h002A; B = 16'h0054; #100;
A = 16'h002A; B = 16'h0055; #100;
A = 16'h002A; B = 16'h0056; #100;
A = 16'h002A; B = 16'h0057; #100;
A = 16'h002A; B = 16'h0058; #100;
A = 16'h002A; B = 16'h0059; #100;
A = 16'h002A; B = 16'h005A; #100;
A = 16'h002A; B = 16'h005B; #100;
A = 16'h002A; B = 16'h005C; #100;
A = 16'h002A; B = 16'h005D; #100;
A = 16'h002A; B = 16'h005E; #100;
A = 16'h002A; B = 16'h005F; #100;
A = 16'h002A; B = 16'h0060; #100;
A = 16'h002A; B = 16'h0061; #100;
A = 16'h002A; B = 16'h0062; #100;
A = 16'h002A; B = 16'h0063; #100;
A = 16'h002A; B = 16'h0064; #100;
A = 16'h002A; B = 16'h0065; #100;
A = 16'h002A; B = 16'h0066; #100;
A = 16'h002A; B = 16'h0067; #100;
A = 16'h002A; B = 16'h0068; #100;
A = 16'h002A; B = 16'h0069; #100;
A = 16'h002A; B = 16'h006A; #100;
A = 16'h002A; B = 16'h006B; #100;
A = 16'h002A; B = 16'h006C; #100;
A = 16'h002A; B = 16'h006D; #100;
A = 16'h002A; B = 16'h006E; #100;
A = 16'h002A; B = 16'h006F; #100;
A = 16'h002A; B = 16'h0070; #100;
A = 16'h002A; B = 16'h0071; #100;
A = 16'h002A; B = 16'h0072; #100;
A = 16'h002A; B = 16'h0073; #100;
A = 16'h002A; B = 16'h0074; #100;
A = 16'h002A; B = 16'h0075; #100;
A = 16'h002A; B = 16'h0076; #100;
A = 16'h002A; B = 16'h0077; #100;
A = 16'h002A; B = 16'h0078; #100;
A = 16'h002A; B = 16'h0079; #100;
A = 16'h002A; B = 16'h007A; #100;
A = 16'h002A; B = 16'h007B; #100;
A = 16'h002A; B = 16'h007C; #100;
A = 16'h002A; B = 16'h007D; #100;
A = 16'h002A; B = 16'h007E; #100;
A = 16'h002A; B = 16'h007F; #100;
A = 16'h002A; B = 16'h0080; #100;
A = 16'h002A; B = 16'h0081; #100;
A = 16'h002A; B = 16'h0082; #100;
A = 16'h002A; B = 16'h0083; #100;
A = 16'h002A; B = 16'h0084; #100;
A = 16'h002A; B = 16'h0085; #100;
A = 16'h002A; B = 16'h0086; #100;
A = 16'h002A; B = 16'h0087; #100;
A = 16'h002A; B = 16'h0088; #100;
A = 16'h002A; B = 16'h0089; #100;
A = 16'h002A; B = 16'h008A; #100;
A = 16'h002A; B = 16'h008B; #100;
A = 16'h002A; B = 16'h008C; #100;
A = 16'h002A; B = 16'h008D; #100;
A = 16'h002A; B = 16'h008E; #100;
A = 16'h002A; B = 16'h008F; #100;
A = 16'h002A; B = 16'h0090; #100;
A = 16'h002A; B = 16'h0091; #100;
A = 16'h002A; B = 16'h0092; #100;
A = 16'h002A; B = 16'h0093; #100;
A = 16'h002A; B = 16'h0094; #100;
A = 16'h002A; B = 16'h0095; #100;
A = 16'h002A; B = 16'h0096; #100;
A = 16'h002A; B = 16'h0097; #100;
A = 16'h002A; B = 16'h0098; #100;
A = 16'h002A; B = 16'h0099; #100;
A = 16'h002A; B = 16'h009A; #100;
A = 16'h002A; B = 16'h009B; #100;
A = 16'h002A; B = 16'h009C; #100;
A = 16'h002A; B = 16'h009D; #100;
A = 16'h002A; B = 16'h009E; #100;
A = 16'h002A; B = 16'h009F; #100;
A = 16'h002A; B = 16'h00A0; #100;
A = 16'h002A; B = 16'h00A1; #100;
A = 16'h002A; B = 16'h00A2; #100;
A = 16'h002A; B = 16'h00A3; #100;
A = 16'h002A; B = 16'h00A4; #100;
A = 16'h002A; B = 16'h00A5; #100;
A = 16'h002A; B = 16'h00A6; #100;
A = 16'h002A; B = 16'h00A7; #100;
A = 16'h002A; B = 16'h00A8; #100;
A = 16'h002A; B = 16'h00A9; #100;
A = 16'h002A; B = 16'h00AA; #100;
A = 16'h002A; B = 16'h00AB; #100;
A = 16'h002A; B = 16'h00AC; #100;
A = 16'h002A; B = 16'h00AD; #100;
A = 16'h002A; B = 16'h00AE; #100;
A = 16'h002A; B = 16'h00AF; #100;
A = 16'h002A; B = 16'h00B0; #100;
A = 16'h002A; B = 16'h00B1; #100;
A = 16'h002A; B = 16'h00B2; #100;
A = 16'h002A; B = 16'h00B3; #100;
A = 16'h002A; B = 16'h00B4; #100;
A = 16'h002A; B = 16'h00B5; #100;
A = 16'h002A; B = 16'h00B6; #100;
A = 16'h002A; B = 16'h00B7; #100;
A = 16'h002A; B = 16'h00B8; #100;
A = 16'h002A; B = 16'h00B9; #100;
A = 16'h002A; B = 16'h00BA; #100;
A = 16'h002A; B = 16'h00BB; #100;
A = 16'h002A; B = 16'h00BC; #100;
A = 16'h002A; B = 16'h00BD; #100;
A = 16'h002A; B = 16'h00BE; #100;
A = 16'h002A; B = 16'h00BF; #100;
A = 16'h002A; B = 16'h00C0; #100;
A = 16'h002A; B = 16'h00C1; #100;
A = 16'h002A; B = 16'h00C2; #100;
A = 16'h002A; B = 16'h00C3; #100;
A = 16'h002A; B = 16'h00C4; #100;
A = 16'h002A; B = 16'h00C5; #100;
A = 16'h002A; B = 16'h00C6; #100;
A = 16'h002A; B = 16'h00C7; #100;
A = 16'h002A; B = 16'h00C8; #100;
A = 16'h002A; B = 16'h00C9; #100;
A = 16'h002A; B = 16'h00CA; #100;
A = 16'h002A; B = 16'h00CB; #100;
A = 16'h002A; B = 16'h00CC; #100;
A = 16'h002A; B = 16'h00CD; #100;
A = 16'h002A; B = 16'h00CE; #100;
A = 16'h002A; B = 16'h00CF; #100;
A = 16'h002A; B = 16'h00D0; #100;
A = 16'h002A; B = 16'h00D1; #100;
A = 16'h002A; B = 16'h00D2; #100;
A = 16'h002A; B = 16'h00D3; #100;
A = 16'h002A; B = 16'h00D4; #100;
A = 16'h002A; B = 16'h00D5; #100;
A = 16'h002A; B = 16'h00D6; #100;
A = 16'h002A; B = 16'h00D7; #100;
A = 16'h002A; B = 16'h00D8; #100;
A = 16'h002A; B = 16'h00D9; #100;
A = 16'h002A; B = 16'h00DA; #100;
A = 16'h002A; B = 16'h00DB; #100;
A = 16'h002A; B = 16'h00DC; #100;
A = 16'h002A; B = 16'h00DD; #100;
A = 16'h002A; B = 16'h00DE; #100;
A = 16'h002A; B = 16'h00DF; #100;
A = 16'h002A; B = 16'h00E0; #100;
A = 16'h002A; B = 16'h00E1; #100;
A = 16'h002A; B = 16'h00E2; #100;
A = 16'h002A; B = 16'h00E3; #100;
A = 16'h002A; B = 16'h00E4; #100;
A = 16'h002A; B = 16'h00E5; #100;
A = 16'h002A; B = 16'h00E6; #100;
A = 16'h002A; B = 16'h00E7; #100;
A = 16'h002A; B = 16'h00E8; #100;
A = 16'h002A; B = 16'h00E9; #100;
A = 16'h002A; B = 16'h00EA; #100;
A = 16'h002A; B = 16'h00EB; #100;
A = 16'h002A; B = 16'h00EC; #100;
A = 16'h002A; B = 16'h00ED; #100;
A = 16'h002A; B = 16'h00EE; #100;
A = 16'h002A; B = 16'h00EF; #100;
A = 16'h002A; B = 16'h00F0; #100;
A = 16'h002A; B = 16'h00F1; #100;
A = 16'h002A; B = 16'h00F2; #100;
A = 16'h002A; B = 16'h00F3; #100;
A = 16'h002A; B = 16'h00F4; #100;
A = 16'h002A; B = 16'h00F5; #100;
A = 16'h002A; B = 16'h00F6; #100;
A = 16'h002A; B = 16'h00F7; #100;
A = 16'h002A; B = 16'h00F8; #100;
A = 16'h002A; B = 16'h00F9; #100;
A = 16'h002A; B = 16'h00FA; #100;
A = 16'h002A; B = 16'h00FB; #100;
A = 16'h002A; B = 16'h00FC; #100;
A = 16'h002A; B = 16'h00FD; #100;
A = 16'h002A; B = 16'h00FE; #100;
A = 16'h002A; B = 16'h00FF; #100;
A = 16'h002B; B = 16'h000; #100;
A = 16'h002B; B = 16'h001; #100;
A = 16'h002B; B = 16'h002; #100;
A = 16'h002B; B = 16'h003; #100;
A = 16'h002B; B = 16'h004; #100;
A = 16'h002B; B = 16'h005; #100;
A = 16'h002B; B = 16'h006; #100;
A = 16'h002B; B = 16'h007; #100;
A = 16'h002B; B = 16'h008; #100;
A = 16'h002B; B = 16'h009; #100;
A = 16'h002B; B = 16'h00A; #100;
A = 16'h002B; B = 16'h00B; #100;
A = 16'h002B; B = 16'h00C; #100;
A = 16'h002B; B = 16'h00D; #100;
A = 16'h002B; B = 16'h00E; #100;
A = 16'h002B; B = 16'h00F; #100;
A = 16'h002B; B = 16'h0010; #100;
A = 16'h002B; B = 16'h0011; #100;
A = 16'h002B; B = 16'h0012; #100;
A = 16'h002B; B = 16'h0013; #100;
A = 16'h002B; B = 16'h0014; #100;
A = 16'h002B; B = 16'h0015; #100;
A = 16'h002B; B = 16'h0016; #100;
A = 16'h002B; B = 16'h0017; #100;
A = 16'h002B; B = 16'h0018; #100;
A = 16'h002B; B = 16'h0019; #100;
A = 16'h002B; B = 16'h001A; #100;
A = 16'h002B; B = 16'h001B; #100;
A = 16'h002B; B = 16'h001C; #100;
A = 16'h002B; B = 16'h001D; #100;
A = 16'h002B; B = 16'h001E; #100;
A = 16'h002B; B = 16'h001F; #100;
A = 16'h002B; B = 16'h0020; #100;
A = 16'h002B; B = 16'h0021; #100;
A = 16'h002B; B = 16'h0022; #100;
A = 16'h002B; B = 16'h0023; #100;
A = 16'h002B; B = 16'h0024; #100;
A = 16'h002B; B = 16'h0025; #100;
A = 16'h002B; B = 16'h0026; #100;
A = 16'h002B; B = 16'h0027; #100;
A = 16'h002B; B = 16'h0028; #100;
A = 16'h002B; B = 16'h0029; #100;
A = 16'h002B; B = 16'h002A; #100;
A = 16'h002B; B = 16'h002B; #100;
A = 16'h002B; B = 16'h002C; #100;
A = 16'h002B; B = 16'h002D; #100;
A = 16'h002B; B = 16'h002E; #100;
A = 16'h002B; B = 16'h002F; #100;
A = 16'h002B; B = 16'h0030; #100;
A = 16'h002B; B = 16'h0031; #100;
A = 16'h002B; B = 16'h0032; #100;
A = 16'h002B; B = 16'h0033; #100;
A = 16'h002B; B = 16'h0034; #100;
A = 16'h002B; B = 16'h0035; #100;
A = 16'h002B; B = 16'h0036; #100;
A = 16'h002B; B = 16'h0037; #100;
A = 16'h002B; B = 16'h0038; #100;
A = 16'h002B; B = 16'h0039; #100;
A = 16'h002B; B = 16'h003A; #100;
A = 16'h002B; B = 16'h003B; #100;
A = 16'h002B; B = 16'h003C; #100;
A = 16'h002B; B = 16'h003D; #100;
A = 16'h002B; B = 16'h003E; #100;
A = 16'h002B; B = 16'h003F; #100;
A = 16'h002B; B = 16'h0040; #100;
A = 16'h002B; B = 16'h0041; #100;
A = 16'h002B; B = 16'h0042; #100;
A = 16'h002B; B = 16'h0043; #100;
A = 16'h002B; B = 16'h0044; #100;
A = 16'h002B; B = 16'h0045; #100;
A = 16'h002B; B = 16'h0046; #100;
A = 16'h002B; B = 16'h0047; #100;
A = 16'h002B; B = 16'h0048; #100;
A = 16'h002B; B = 16'h0049; #100;
A = 16'h002B; B = 16'h004A; #100;
A = 16'h002B; B = 16'h004B; #100;
A = 16'h002B; B = 16'h004C; #100;
A = 16'h002B; B = 16'h004D; #100;
A = 16'h002B; B = 16'h004E; #100;
A = 16'h002B; B = 16'h004F; #100;
A = 16'h002B; B = 16'h0050; #100;
A = 16'h002B; B = 16'h0051; #100;
A = 16'h002B; B = 16'h0052; #100;
A = 16'h002B; B = 16'h0053; #100;
A = 16'h002B; B = 16'h0054; #100;
A = 16'h002B; B = 16'h0055; #100;
A = 16'h002B; B = 16'h0056; #100;
A = 16'h002B; B = 16'h0057; #100;
A = 16'h002B; B = 16'h0058; #100;
A = 16'h002B; B = 16'h0059; #100;
A = 16'h002B; B = 16'h005A; #100;
A = 16'h002B; B = 16'h005B; #100;
A = 16'h002B; B = 16'h005C; #100;
A = 16'h002B; B = 16'h005D; #100;
A = 16'h002B; B = 16'h005E; #100;
A = 16'h002B; B = 16'h005F; #100;
A = 16'h002B; B = 16'h0060; #100;
A = 16'h002B; B = 16'h0061; #100;
A = 16'h002B; B = 16'h0062; #100;
A = 16'h002B; B = 16'h0063; #100;
A = 16'h002B; B = 16'h0064; #100;
A = 16'h002B; B = 16'h0065; #100;
A = 16'h002B; B = 16'h0066; #100;
A = 16'h002B; B = 16'h0067; #100;
A = 16'h002B; B = 16'h0068; #100;
A = 16'h002B; B = 16'h0069; #100;
A = 16'h002B; B = 16'h006A; #100;
A = 16'h002B; B = 16'h006B; #100;
A = 16'h002B; B = 16'h006C; #100;
A = 16'h002B; B = 16'h006D; #100;
A = 16'h002B; B = 16'h006E; #100;
A = 16'h002B; B = 16'h006F; #100;
A = 16'h002B; B = 16'h0070; #100;
A = 16'h002B; B = 16'h0071; #100;
A = 16'h002B; B = 16'h0072; #100;
A = 16'h002B; B = 16'h0073; #100;
A = 16'h002B; B = 16'h0074; #100;
A = 16'h002B; B = 16'h0075; #100;
A = 16'h002B; B = 16'h0076; #100;
A = 16'h002B; B = 16'h0077; #100;
A = 16'h002B; B = 16'h0078; #100;
A = 16'h002B; B = 16'h0079; #100;
A = 16'h002B; B = 16'h007A; #100;
A = 16'h002B; B = 16'h007B; #100;
A = 16'h002B; B = 16'h007C; #100;
A = 16'h002B; B = 16'h007D; #100;
A = 16'h002B; B = 16'h007E; #100;
A = 16'h002B; B = 16'h007F; #100;
A = 16'h002B; B = 16'h0080; #100;
A = 16'h002B; B = 16'h0081; #100;
A = 16'h002B; B = 16'h0082; #100;
A = 16'h002B; B = 16'h0083; #100;
A = 16'h002B; B = 16'h0084; #100;
A = 16'h002B; B = 16'h0085; #100;
A = 16'h002B; B = 16'h0086; #100;
A = 16'h002B; B = 16'h0087; #100;
A = 16'h002B; B = 16'h0088; #100;
A = 16'h002B; B = 16'h0089; #100;
A = 16'h002B; B = 16'h008A; #100;
A = 16'h002B; B = 16'h008B; #100;
A = 16'h002B; B = 16'h008C; #100;
A = 16'h002B; B = 16'h008D; #100;
A = 16'h002B; B = 16'h008E; #100;
A = 16'h002B; B = 16'h008F; #100;
A = 16'h002B; B = 16'h0090; #100;
A = 16'h002B; B = 16'h0091; #100;
A = 16'h002B; B = 16'h0092; #100;
A = 16'h002B; B = 16'h0093; #100;
A = 16'h002B; B = 16'h0094; #100;
A = 16'h002B; B = 16'h0095; #100;
A = 16'h002B; B = 16'h0096; #100;
A = 16'h002B; B = 16'h0097; #100;
A = 16'h002B; B = 16'h0098; #100;
A = 16'h002B; B = 16'h0099; #100;
A = 16'h002B; B = 16'h009A; #100;
A = 16'h002B; B = 16'h009B; #100;
A = 16'h002B; B = 16'h009C; #100;
A = 16'h002B; B = 16'h009D; #100;
A = 16'h002B; B = 16'h009E; #100;
A = 16'h002B; B = 16'h009F; #100;
A = 16'h002B; B = 16'h00A0; #100;
A = 16'h002B; B = 16'h00A1; #100;
A = 16'h002B; B = 16'h00A2; #100;
A = 16'h002B; B = 16'h00A3; #100;
A = 16'h002B; B = 16'h00A4; #100;
A = 16'h002B; B = 16'h00A5; #100;
A = 16'h002B; B = 16'h00A6; #100;
A = 16'h002B; B = 16'h00A7; #100;
A = 16'h002B; B = 16'h00A8; #100;
A = 16'h002B; B = 16'h00A9; #100;
A = 16'h002B; B = 16'h00AA; #100;
A = 16'h002B; B = 16'h00AB; #100;
A = 16'h002B; B = 16'h00AC; #100;
A = 16'h002B; B = 16'h00AD; #100;
A = 16'h002B; B = 16'h00AE; #100;
A = 16'h002B; B = 16'h00AF; #100;
A = 16'h002B; B = 16'h00B0; #100;
A = 16'h002B; B = 16'h00B1; #100;
A = 16'h002B; B = 16'h00B2; #100;
A = 16'h002B; B = 16'h00B3; #100;
A = 16'h002B; B = 16'h00B4; #100;
A = 16'h002B; B = 16'h00B5; #100;
A = 16'h002B; B = 16'h00B6; #100;
A = 16'h002B; B = 16'h00B7; #100;
A = 16'h002B; B = 16'h00B8; #100;
A = 16'h002B; B = 16'h00B9; #100;
A = 16'h002B; B = 16'h00BA; #100;
A = 16'h002B; B = 16'h00BB; #100;
A = 16'h002B; B = 16'h00BC; #100;
A = 16'h002B; B = 16'h00BD; #100;
A = 16'h002B; B = 16'h00BE; #100;
A = 16'h002B; B = 16'h00BF; #100;
A = 16'h002B; B = 16'h00C0; #100;
A = 16'h002B; B = 16'h00C1; #100;
A = 16'h002B; B = 16'h00C2; #100;
A = 16'h002B; B = 16'h00C3; #100;
A = 16'h002B; B = 16'h00C4; #100;
A = 16'h002B; B = 16'h00C5; #100;
A = 16'h002B; B = 16'h00C6; #100;
A = 16'h002B; B = 16'h00C7; #100;
A = 16'h002B; B = 16'h00C8; #100;
A = 16'h002B; B = 16'h00C9; #100;
A = 16'h002B; B = 16'h00CA; #100;
A = 16'h002B; B = 16'h00CB; #100;
A = 16'h002B; B = 16'h00CC; #100;
A = 16'h002B; B = 16'h00CD; #100;
A = 16'h002B; B = 16'h00CE; #100;
A = 16'h002B; B = 16'h00CF; #100;
A = 16'h002B; B = 16'h00D0; #100;
A = 16'h002B; B = 16'h00D1; #100;
A = 16'h002B; B = 16'h00D2; #100;
A = 16'h002B; B = 16'h00D3; #100;
A = 16'h002B; B = 16'h00D4; #100;
A = 16'h002B; B = 16'h00D5; #100;
A = 16'h002B; B = 16'h00D6; #100;
A = 16'h002B; B = 16'h00D7; #100;
A = 16'h002B; B = 16'h00D8; #100;
A = 16'h002B; B = 16'h00D9; #100;
A = 16'h002B; B = 16'h00DA; #100;
A = 16'h002B; B = 16'h00DB; #100;
A = 16'h002B; B = 16'h00DC; #100;
A = 16'h002B; B = 16'h00DD; #100;
A = 16'h002B; B = 16'h00DE; #100;
A = 16'h002B; B = 16'h00DF; #100;
A = 16'h002B; B = 16'h00E0; #100;
A = 16'h002B; B = 16'h00E1; #100;
A = 16'h002B; B = 16'h00E2; #100;
A = 16'h002B; B = 16'h00E3; #100;
A = 16'h002B; B = 16'h00E4; #100;
A = 16'h002B; B = 16'h00E5; #100;
A = 16'h002B; B = 16'h00E6; #100;
A = 16'h002B; B = 16'h00E7; #100;
A = 16'h002B; B = 16'h00E8; #100;
A = 16'h002B; B = 16'h00E9; #100;
A = 16'h002B; B = 16'h00EA; #100;
A = 16'h002B; B = 16'h00EB; #100;
A = 16'h002B; B = 16'h00EC; #100;
A = 16'h002B; B = 16'h00ED; #100;
A = 16'h002B; B = 16'h00EE; #100;
A = 16'h002B; B = 16'h00EF; #100;
A = 16'h002B; B = 16'h00F0; #100;
A = 16'h002B; B = 16'h00F1; #100;
A = 16'h002B; B = 16'h00F2; #100;
A = 16'h002B; B = 16'h00F3; #100;
A = 16'h002B; B = 16'h00F4; #100;
A = 16'h002B; B = 16'h00F5; #100;
A = 16'h002B; B = 16'h00F6; #100;
A = 16'h002B; B = 16'h00F7; #100;
A = 16'h002B; B = 16'h00F8; #100;
A = 16'h002B; B = 16'h00F9; #100;
A = 16'h002B; B = 16'h00FA; #100;
A = 16'h002B; B = 16'h00FB; #100;
A = 16'h002B; B = 16'h00FC; #100;
A = 16'h002B; B = 16'h00FD; #100;
A = 16'h002B; B = 16'h00FE; #100;
A = 16'h002B; B = 16'h00FF; #100;
A = 16'h002C; B = 16'h000; #100;
A = 16'h002C; B = 16'h001; #100;
A = 16'h002C; B = 16'h002; #100;
A = 16'h002C; B = 16'h003; #100;
A = 16'h002C; B = 16'h004; #100;
A = 16'h002C; B = 16'h005; #100;
A = 16'h002C; B = 16'h006; #100;
A = 16'h002C; B = 16'h007; #100;
A = 16'h002C; B = 16'h008; #100;
A = 16'h002C; B = 16'h009; #100;
A = 16'h002C; B = 16'h00A; #100;
A = 16'h002C; B = 16'h00B; #100;
A = 16'h002C; B = 16'h00C; #100;
A = 16'h002C; B = 16'h00D; #100;
A = 16'h002C; B = 16'h00E; #100;
A = 16'h002C; B = 16'h00F; #100;
A = 16'h002C; B = 16'h0010; #100;
A = 16'h002C; B = 16'h0011; #100;
A = 16'h002C; B = 16'h0012; #100;
A = 16'h002C; B = 16'h0013; #100;
A = 16'h002C; B = 16'h0014; #100;
A = 16'h002C; B = 16'h0015; #100;
A = 16'h002C; B = 16'h0016; #100;
A = 16'h002C; B = 16'h0017; #100;
A = 16'h002C; B = 16'h0018; #100;
A = 16'h002C; B = 16'h0019; #100;
A = 16'h002C; B = 16'h001A; #100;
A = 16'h002C; B = 16'h001B; #100;
A = 16'h002C; B = 16'h001C; #100;
A = 16'h002C; B = 16'h001D; #100;
A = 16'h002C; B = 16'h001E; #100;
A = 16'h002C; B = 16'h001F; #100;
A = 16'h002C; B = 16'h0020; #100;
A = 16'h002C; B = 16'h0021; #100;
A = 16'h002C; B = 16'h0022; #100;
A = 16'h002C; B = 16'h0023; #100;
A = 16'h002C; B = 16'h0024; #100;
A = 16'h002C; B = 16'h0025; #100;
A = 16'h002C; B = 16'h0026; #100;
A = 16'h002C; B = 16'h0027; #100;
A = 16'h002C; B = 16'h0028; #100;
A = 16'h002C; B = 16'h0029; #100;
A = 16'h002C; B = 16'h002A; #100;
A = 16'h002C; B = 16'h002B; #100;
A = 16'h002C; B = 16'h002C; #100;
A = 16'h002C; B = 16'h002D; #100;
A = 16'h002C; B = 16'h002E; #100;
A = 16'h002C; B = 16'h002F; #100;
A = 16'h002C; B = 16'h0030; #100;
A = 16'h002C; B = 16'h0031; #100;
A = 16'h002C; B = 16'h0032; #100;
A = 16'h002C; B = 16'h0033; #100;
A = 16'h002C; B = 16'h0034; #100;
A = 16'h002C; B = 16'h0035; #100;
A = 16'h002C; B = 16'h0036; #100;
A = 16'h002C; B = 16'h0037; #100;
A = 16'h002C; B = 16'h0038; #100;
A = 16'h002C; B = 16'h0039; #100;
A = 16'h002C; B = 16'h003A; #100;
A = 16'h002C; B = 16'h003B; #100;
A = 16'h002C; B = 16'h003C; #100;
A = 16'h002C; B = 16'h003D; #100;
A = 16'h002C; B = 16'h003E; #100;
A = 16'h002C; B = 16'h003F; #100;
A = 16'h002C; B = 16'h0040; #100;
A = 16'h002C; B = 16'h0041; #100;
A = 16'h002C; B = 16'h0042; #100;
A = 16'h002C; B = 16'h0043; #100;
A = 16'h002C; B = 16'h0044; #100;
A = 16'h002C; B = 16'h0045; #100;
A = 16'h002C; B = 16'h0046; #100;
A = 16'h002C; B = 16'h0047; #100;
A = 16'h002C; B = 16'h0048; #100;
A = 16'h002C; B = 16'h0049; #100;
A = 16'h002C; B = 16'h004A; #100;
A = 16'h002C; B = 16'h004B; #100;
A = 16'h002C; B = 16'h004C; #100;
A = 16'h002C; B = 16'h004D; #100;
A = 16'h002C; B = 16'h004E; #100;
A = 16'h002C; B = 16'h004F; #100;
A = 16'h002C; B = 16'h0050; #100;
A = 16'h002C; B = 16'h0051; #100;
A = 16'h002C; B = 16'h0052; #100;
A = 16'h002C; B = 16'h0053; #100;
A = 16'h002C; B = 16'h0054; #100;
A = 16'h002C; B = 16'h0055; #100;
A = 16'h002C; B = 16'h0056; #100;
A = 16'h002C; B = 16'h0057; #100;
A = 16'h002C; B = 16'h0058; #100;
A = 16'h002C; B = 16'h0059; #100;
A = 16'h002C; B = 16'h005A; #100;
A = 16'h002C; B = 16'h005B; #100;
A = 16'h002C; B = 16'h005C; #100;
A = 16'h002C; B = 16'h005D; #100;
A = 16'h002C; B = 16'h005E; #100;
A = 16'h002C; B = 16'h005F; #100;
A = 16'h002C; B = 16'h0060; #100;
A = 16'h002C; B = 16'h0061; #100;
A = 16'h002C; B = 16'h0062; #100;
A = 16'h002C; B = 16'h0063; #100;
A = 16'h002C; B = 16'h0064; #100;
A = 16'h002C; B = 16'h0065; #100;
A = 16'h002C; B = 16'h0066; #100;
A = 16'h002C; B = 16'h0067; #100;
A = 16'h002C; B = 16'h0068; #100;
A = 16'h002C; B = 16'h0069; #100;
A = 16'h002C; B = 16'h006A; #100;
A = 16'h002C; B = 16'h006B; #100;
A = 16'h002C; B = 16'h006C; #100;
A = 16'h002C; B = 16'h006D; #100;
A = 16'h002C; B = 16'h006E; #100;
A = 16'h002C; B = 16'h006F; #100;
A = 16'h002C; B = 16'h0070; #100;
A = 16'h002C; B = 16'h0071; #100;
A = 16'h002C; B = 16'h0072; #100;
A = 16'h002C; B = 16'h0073; #100;
A = 16'h002C; B = 16'h0074; #100;
A = 16'h002C; B = 16'h0075; #100;
A = 16'h002C; B = 16'h0076; #100;
A = 16'h002C; B = 16'h0077; #100;
A = 16'h002C; B = 16'h0078; #100;
A = 16'h002C; B = 16'h0079; #100;
A = 16'h002C; B = 16'h007A; #100;
A = 16'h002C; B = 16'h007B; #100;
A = 16'h002C; B = 16'h007C; #100;
A = 16'h002C; B = 16'h007D; #100;
A = 16'h002C; B = 16'h007E; #100;
A = 16'h002C; B = 16'h007F; #100;
A = 16'h002C; B = 16'h0080; #100;
A = 16'h002C; B = 16'h0081; #100;
A = 16'h002C; B = 16'h0082; #100;
A = 16'h002C; B = 16'h0083; #100;
A = 16'h002C; B = 16'h0084; #100;
A = 16'h002C; B = 16'h0085; #100;
A = 16'h002C; B = 16'h0086; #100;
A = 16'h002C; B = 16'h0087; #100;
A = 16'h002C; B = 16'h0088; #100;
A = 16'h002C; B = 16'h0089; #100;
A = 16'h002C; B = 16'h008A; #100;
A = 16'h002C; B = 16'h008B; #100;
A = 16'h002C; B = 16'h008C; #100;
A = 16'h002C; B = 16'h008D; #100;
A = 16'h002C; B = 16'h008E; #100;
A = 16'h002C; B = 16'h008F; #100;
A = 16'h002C; B = 16'h0090; #100;
A = 16'h002C; B = 16'h0091; #100;
A = 16'h002C; B = 16'h0092; #100;
A = 16'h002C; B = 16'h0093; #100;
A = 16'h002C; B = 16'h0094; #100;
A = 16'h002C; B = 16'h0095; #100;
A = 16'h002C; B = 16'h0096; #100;
A = 16'h002C; B = 16'h0097; #100;
A = 16'h002C; B = 16'h0098; #100;
A = 16'h002C; B = 16'h0099; #100;
A = 16'h002C; B = 16'h009A; #100;
A = 16'h002C; B = 16'h009B; #100;
A = 16'h002C; B = 16'h009C; #100;
A = 16'h002C; B = 16'h009D; #100;
A = 16'h002C; B = 16'h009E; #100;
A = 16'h002C; B = 16'h009F; #100;
A = 16'h002C; B = 16'h00A0; #100;
A = 16'h002C; B = 16'h00A1; #100;
A = 16'h002C; B = 16'h00A2; #100;
A = 16'h002C; B = 16'h00A3; #100;
A = 16'h002C; B = 16'h00A4; #100;
A = 16'h002C; B = 16'h00A5; #100;
A = 16'h002C; B = 16'h00A6; #100;
A = 16'h002C; B = 16'h00A7; #100;
A = 16'h002C; B = 16'h00A8; #100;
A = 16'h002C; B = 16'h00A9; #100;
A = 16'h002C; B = 16'h00AA; #100;
A = 16'h002C; B = 16'h00AB; #100;
A = 16'h002C; B = 16'h00AC; #100;
A = 16'h002C; B = 16'h00AD; #100;
A = 16'h002C; B = 16'h00AE; #100;
A = 16'h002C; B = 16'h00AF; #100;
A = 16'h002C; B = 16'h00B0; #100;
A = 16'h002C; B = 16'h00B1; #100;
A = 16'h002C; B = 16'h00B2; #100;
A = 16'h002C; B = 16'h00B3; #100;
A = 16'h002C; B = 16'h00B4; #100;
A = 16'h002C; B = 16'h00B5; #100;
A = 16'h002C; B = 16'h00B6; #100;
A = 16'h002C; B = 16'h00B7; #100;
A = 16'h002C; B = 16'h00B8; #100;
A = 16'h002C; B = 16'h00B9; #100;
A = 16'h002C; B = 16'h00BA; #100;
A = 16'h002C; B = 16'h00BB; #100;
A = 16'h002C; B = 16'h00BC; #100;
A = 16'h002C; B = 16'h00BD; #100;
A = 16'h002C; B = 16'h00BE; #100;
A = 16'h002C; B = 16'h00BF; #100;
A = 16'h002C; B = 16'h00C0; #100;
A = 16'h002C; B = 16'h00C1; #100;
A = 16'h002C; B = 16'h00C2; #100;
A = 16'h002C; B = 16'h00C3; #100;
A = 16'h002C; B = 16'h00C4; #100;
A = 16'h002C; B = 16'h00C5; #100;
A = 16'h002C; B = 16'h00C6; #100;
A = 16'h002C; B = 16'h00C7; #100;
A = 16'h002C; B = 16'h00C8; #100;
A = 16'h002C; B = 16'h00C9; #100;
A = 16'h002C; B = 16'h00CA; #100;
A = 16'h002C; B = 16'h00CB; #100;
A = 16'h002C; B = 16'h00CC; #100;
A = 16'h002C; B = 16'h00CD; #100;
A = 16'h002C; B = 16'h00CE; #100;
A = 16'h002C; B = 16'h00CF; #100;
A = 16'h002C; B = 16'h00D0; #100;
A = 16'h002C; B = 16'h00D1; #100;
A = 16'h002C; B = 16'h00D2; #100;
A = 16'h002C; B = 16'h00D3; #100;
A = 16'h002C; B = 16'h00D4; #100;
A = 16'h002C; B = 16'h00D5; #100;
A = 16'h002C; B = 16'h00D6; #100;
A = 16'h002C; B = 16'h00D7; #100;
A = 16'h002C; B = 16'h00D8; #100;
A = 16'h002C; B = 16'h00D9; #100;
A = 16'h002C; B = 16'h00DA; #100;
A = 16'h002C; B = 16'h00DB; #100;
A = 16'h002C; B = 16'h00DC; #100;
A = 16'h002C; B = 16'h00DD; #100;
A = 16'h002C; B = 16'h00DE; #100;
A = 16'h002C; B = 16'h00DF; #100;
A = 16'h002C; B = 16'h00E0; #100;
A = 16'h002C; B = 16'h00E1; #100;
A = 16'h002C; B = 16'h00E2; #100;
A = 16'h002C; B = 16'h00E3; #100;
A = 16'h002C; B = 16'h00E4; #100;
A = 16'h002C; B = 16'h00E5; #100;
A = 16'h002C; B = 16'h00E6; #100;
A = 16'h002C; B = 16'h00E7; #100;
A = 16'h002C; B = 16'h00E8; #100;
A = 16'h002C; B = 16'h00E9; #100;
A = 16'h002C; B = 16'h00EA; #100;
A = 16'h002C; B = 16'h00EB; #100;
A = 16'h002C; B = 16'h00EC; #100;
A = 16'h002C; B = 16'h00ED; #100;
A = 16'h002C; B = 16'h00EE; #100;
A = 16'h002C; B = 16'h00EF; #100;
A = 16'h002C; B = 16'h00F0; #100;
A = 16'h002C; B = 16'h00F1; #100;
A = 16'h002C; B = 16'h00F2; #100;
A = 16'h002C; B = 16'h00F3; #100;
A = 16'h002C; B = 16'h00F4; #100;
A = 16'h002C; B = 16'h00F5; #100;
A = 16'h002C; B = 16'h00F6; #100;
A = 16'h002C; B = 16'h00F7; #100;
A = 16'h002C; B = 16'h00F8; #100;
A = 16'h002C; B = 16'h00F9; #100;
A = 16'h002C; B = 16'h00FA; #100;
A = 16'h002C; B = 16'h00FB; #100;
A = 16'h002C; B = 16'h00FC; #100;
A = 16'h002C; B = 16'h00FD; #100;
A = 16'h002C; B = 16'h00FE; #100;
A = 16'h002C; B = 16'h00FF; #100;
A = 16'h002D; B = 16'h000; #100;
A = 16'h002D; B = 16'h001; #100;
A = 16'h002D; B = 16'h002; #100;
A = 16'h002D; B = 16'h003; #100;
A = 16'h002D; B = 16'h004; #100;
A = 16'h002D; B = 16'h005; #100;
A = 16'h002D; B = 16'h006; #100;
A = 16'h002D; B = 16'h007; #100;
A = 16'h002D; B = 16'h008; #100;
A = 16'h002D; B = 16'h009; #100;
A = 16'h002D; B = 16'h00A; #100;
A = 16'h002D; B = 16'h00B; #100;
A = 16'h002D; B = 16'h00C; #100;
A = 16'h002D; B = 16'h00D; #100;
A = 16'h002D; B = 16'h00E; #100;
A = 16'h002D; B = 16'h00F; #100;
A = 16'h002D; B = 16'h0010; #100;
A = 16'h002D; B = 16'h0011; #100;
A = 16'h002D; B = 16'h0012; #100;
A = 16'h002D; B = 16'h0013; #100;
A = 16'h002D; B = 16'h0014; #100;
A = 16'h002D; B = 16'h0015; #100;
A = 16'h002D; B = 16'h0016; #100;
A = 16'h002D; B = 16'h0017; #100;
A = 16'h002D; B = 16'h0018; #100;
A = 16'h002D; B = 16'h0019; #100;
A = 16'h002D; B = 16'h001A; #100;
A = 16'h002D; B = 16'h001B; #100;
A = 16'h002D; B = 16'h001C; #100;
A = 16'h002D; B = 16'h001D; #100;
A = 16'h002D; B = 16'h001E; #100;
A = 16'h002D; B = 16'h001F; #100;
A = 16'h002D; B = 16'h0020; #100;
A = 16'h002D; B = 16'h0021; #100;
A = 16'h002D; B = 16'h0022; #100;
A = 16'h002D; B = 16'h0023; #100;
A = 16'h002D; B = 16'h0024; #100;
A = 16'h002D; B = 16'h0025; #100;
A = 16'h002D; B = 16'h0026; #100;
A = 16'h002D; B = 16'h0027; #100;
A = 16'h002D; B = 16'h0028; #100;
A = 16'h002D; B = 16'h0029; #100;
A = 16'h002D; B = 16'h002A; #100;
A = 16'h002D; B = 16'h002B; #100;
A = 16'h002D; B = 16'h002C; #100;
A = 16'h002D; B = 16'h002D; #100;
A = 16'h002D; B = 16'h002E; #100;
A = 16'h002D; B = 16'h002F; #100;
A = 16'h002D; B = 16'h0030; #100;
A = 16'h002D; B = 16'h0031; #100;
A = 16'h002D; B = 16'h0032; #100;
A = 16'h002D; B = 16'h0033; #100;
A = 16'h002D; B = 16'h0034; #100;
A = 16'h002D; B = 16'h0035; #100;
A = 16'h002D; B = 16'h0036; #100;
A = 16'h002D; B = 16'h0037; #100;
A = 16'h002D; B = 16'h0038; #100;
A = 16'h002D; B = 16'h0039; #100;
A = 16'h002D; B = 16'h003A; #100;
A = 16'h002D; B = 16'h003B; #100;
A = 16'h002D; B = 16'h003C; #100;
A = 16'h002D; B = 16'h003D; #100;
A = 16'h002D; B = 16'h003E; #100;
A = 16'h002D; B = 16'h003F; #100;
A = 16'h002D; B = 16'h0040; #100;
A = 16'h002D; B = 16'h0041; #100;
A = 16'h002D; B = 16'h0042; #100;
A = 16'h002D; B = 16'h0043; #100;
A = 16'h002D; B = 16'h0044; #100;
A = 16'h002D; B = 16'h0045; #100;
A = 16'h002D; B = 16'h0046; #100;
A = 16'h002D; B = 16'h0047; #100;
A = 16'h002D; B = 16'h0048; #100;
A = 16'h002D; B = 16'h0049; #100;
A = 16'h002D; B = 16'h004A; #100;
A = 16'h002D; B = 16'h004B; #100;
A = 16'h002D; B = 16'h004C; #100;
A = 16'h002D; B = 16'h004D; #100;
A = 16'h002D; B = 16'h004E; #100;
A = 16'h002D; B = 16'h004F; #100;
A = 16'h002D; B = 16'h0050; #100;
A = 16'h002D; B = 16'h0051; #100;
A = 16'h002D; B = 16'h0052; #100;
A = 16'h002D; B = 16'h0053; #100;
A = 16'h002D; B = 16'h0054; #100;
A = 16'h002D; B = 16'h0055; #100;
A = 16'h002D; B = 16'h0056; #100;
A = 16'h002D; B = 16'h0057; #100;
A = 16'h002D; B = 16'h0058; #100;
A = 16'h002D; B = 16'h0059; #100;
A = 16'h002D; B = 16'h005A; #100;
A = 16'h002D; B = 16'h005B; #100;
A = 16'h002D; B = 16'h005C; #100;
A = 16'h002D; B = 16'h005D; #100;
A = 16'h002D; B = 16'h005E; #100;
A = 16'h002D; B = 16'h005F; #100;
A = 16'h002D; B = 16'h0060; #100;
A = 16'h002D; B = 16'h0061; #100;
A = 16'h002D; B = 16'h0062; #100;
A = 16'h002D; B = 16'h0063; #100;
A = 16'h002D; B = 16'h0064; #100;
A = 16'h002D; B = 16'h0065; #100;
A = 16'h002D; B = 16'h0066; #100;
A = 16'h002D; B = 16'h0067; #100;
A = 16'h002D; B = 16'h0068; #100;
A = 16'h002D; B = 16'h0069; #100;
A = 16'h002D; B = 16'h006A; #100;
A = 16'h002D; B = 16'h006B; #100;
A = 16'h002D; B = 16'h006C; #100;
A = 16'h002D; B = 16'h006D; #100;
A = 16'h002D; B = 16'h006E; #100;
A = 16'h002D; B = 16'h006F; #100;
A = 16'h002D; B = 16'h0070; #100;
A = 16'h002D; B = 16'h0071; #100;
A = 16'h002D; B = 16'h0072; #100;
A = 16'h002D; B = 16'h0073; #100;
A = 16'h002D; B = 16'h0074; #100;
A = 16'h002D; B = 16'h0075; #100;
A = 16'h002D; B = 16'h0076; #100;
A = 16'h002D; B = 16'h0077; #100;
A = 16'h002D; B = 16'h0078; #100;
A = 16'h002D; B = 16'h0079; #100;
A = 16'h002D; B = 16'h007A; #100;
A = 16'h002D; B = 16'h007B; #100;
A = 16'h002D; B = 16'h007C; #100;
A = 16'h002D; B = 16'h007D; #100;
A = 16'h002D; B = 16'h007E; #100;
A = 16'h002D; B = 16'h007F; #100;
A = 16'h002D; B = 16'h0080; #100;
A = 16'h002D; B = 16'h0081; #100;
A = 16'h002D; B = 16'h0082; #100;
A = 16'h002D; B = 16'h0083; #100;
A = 16'h002D; B = 16'h0084; #100;
A = 16'h002D; B = 16'h0085; #100;
A = 16'h002D; B = 16'h0086; #100;
A = 16'h002D; B = 16'h0087; #100;
A = 16'h002D; B = 16'h0088; #100;
A = 16'h002D; B = 16'h0089; #100;
A = 16'h002D; B = 16'h008A; #100;
A = 16'h002D; B = 16'h008B; #100;
A = 16'h002D; B = 16'h008C; #100;
A = 16'h002D; B = 16'h008D; #100;
A = 16'h002D; B = 16'h008E; #100;
A = 16'h002D; B = 16'h008F; #100;
A = 16'h002D; B = 16'h0090; #100;
A = 16'h002D; B = 16'h0091; #100;
A = 16'h002D; B = 16'h0092; #100;
A = 16'h002D; B = 16'h0093; #100;
A = 16'h002D; B = 16'h0094; #100;
A = 16'h002D; B = 16'h0095; #100;
A = 16'h002D; B = 16'h0096; #100;
A = 16'h002D; B = 16'h0097; #100;
A = 16'h002D; B = 16'h0098; #100;
A = 16'h002D; B = 16'h0099; #100;
A = 16'h002D; B = 16'h009A; #100;
A = 16'h002D; B = 16'h009B; #100;
A = 16'h002D; B = 16'h009C; #100;
A = 16'h002D; B = 16'h009D; #100;
A = 16'h002D; B = 16'h009E; #100;
A = 16'h002D; B = 16'h009F; #100;
A = 16'h002D; B = 16'h00A0; #100;
A = 16'h002D; B = 16'h00A1; #100;
A = 16'h002D; B = 16'h00A2; #100;
A = 16'h002D; B = 16'h00A3; #100;
A = 16'h002D; B = 16'h00A4; #100;
A = 16'h002D; B = 16'h00A5; #100;
A = 16'h002D; B = 16'h00A6; #100;
A = 16'h002D; B = 16'h00A7; #100;
A = 16'h002D; B = 16'h00A8; #100;
A = 16'h002D; B = 16'h00A9; #100;
A = 16'h002D; B = 16'h00AA; #100;
A = 16'h002D; B = 16'h00AB; #100;
A = 16'h002D; B = 16'h00AC; #100;
A = 16'h002D; B = 16'h00AD; #100;
A = 16'h002D; B = 16'h00AE; #100;
A = 16'h002D; B = 16'h00AF; #100;
A = 16'h002D; B = 16'h00B0; #100;
A = 16'h002D; B = 16'h00B1; #100;
A = 16'h002D; B = 16'h00B2; #100;
A = 16'h002D; B = 16'h00B3; #100;
A = 16'h002D; B = 16'h00B4; #100;
A = 16'h002D; B = 16'h00B5; #100;
A = 16'h002D; B = 16'h00B6; #100;
A = 16'h002D; B = 16'h00B7; #100;
A = 16'h002D; B = 16'h00B8; #100;
A = 16'h002D; B = 16'h00B9; #100;
A = 16'h002D; B = 16'h00BA; #100;
A = 16'h002D; B = 16'h00BB; #100;
A = 16'h002D; B = 16'h00BC; #100;
A = 16'h002D; B = 16'h00BD; #100;
A = 16'h002D; B = 16'h00BE; #100;
A = 16'h002D; B = 16'h00BF; #100;
A = 16'h002D; B = 16'h00C0; #100;
A = 16'h002D; B = 16'h00C1; #100;
A = 16'h002D; B = 16'h00C2; #100;
A = 16'h002D; B = 16'h00C3; #100;
A = 16'h002D; B = 16'h00C4; #100;
A = 16'h002D; B = 16'h00C5; #100;
A = 16'h002D; B = 16'h00C6; #100;
A = 16'h002D; B = 16'h00C7; #100;
A = 16'h002D; B = 16'h00C8; #100;
A = 16'h002D; B = 16'h00C9; #100;
A = 16'h002D; B = 16'h00CA; #100;
A = 16'h002D; B = 16'h00CB; #100;
A = 16'h002D; B = 16'h00CC; #100;
A = 16'h002D; B = 16'h00CD; #100;
A = 16'h002D; B = 16'h00CE; #100;
A = 16'h002D; B = 16'h00CF; #100;
A = 16'h002D; B = 16'h00D0; #100;
A = 16'h002D; B = 16'h00D1; #100;
A = 16'h002D; B = 16'h00D2; #100;
A = 16'h002D; B = 16'h00D3; #100;
A = 16'h002D; B = 16'h00D4; #100;
A = 16'h002D; B = 16'h00D5; #100;
A = 16'h002D; B = 16'h00D6; #100;
A = 16'h002D; B = 16'h00D7; #100;
A = 16'h002D; B = 16'h00D8; #100;
A = 16'h002D; B = 16'h00D9; #100;
A = 16'h002D; B = 16'h00DA; #100;
A = 16'h002D; B = 16'h00DB; #100;
A = 16'h002D; B = 16'h00DC; #100;
A = 16'h002D; B = 16'h00DD; #100;
A = 16'h002D; B = 16'h00DE; #100;
A = 16'h002D; B = 16'h00DF; #100;
A = 16'h002D; B = 16'h00E0; #100;
A = 16'h002D; B = 16'h00E1; #100;
A = 16'h002D; B = 16'h00E2; #100;
A = 16'h002D; B = 16'h00E3; #100;
A = 16'h002D; B = 16'h00E4; #100;
A = 16'h002D; B = 16'h00E5; #100;
A = 16'h002D; B = 16'h00E6; #100;
A = 16'h002D; B = 16'h00E7; #100;
A = 16'h002D; B = 16'h00E8; #100;
A = 16'h002D; B = 16'h00E9; #100;
A = 16'h002D; B = 16'h00EA; #100;
A = 16'h002D; B = 16'h00EB; #100;
A = 16'h002D; B = 16'h00EC; #100;
A = 16'h002D; B = 16'h00ED; #100;
A = 16'h002D; B = 16'h00EE; #100;
A = 16'h002D; B = 16'h00EF; #100;
A = 16'h002D; B = 16'h00F0; #100;
A = 16'h002D; B = 16'h00F1; #100;
A = 16'h002D; B = 16'h00F2; #100;
A = 16'h002D; B = 16'h00F3; #100;
A = 16'h002D; B = 16'h00F4; #100;
A = 16'h002D; B = 16'h00F5; #100;
A = 16'h002D; B = 16'h00F6; #100;
A = 16'h002D; B = 16'h00F7; #100;
A = 16'h002D; B = 16'h00F8; #100;
A = 16'h002D; B = 16'h00F9; #100;
A = 16'h002D; B = 16'h00FA; #100;
A = 16'h002D; B = 16'h00FB; #100;
A = 16'h002D; B = 16'h00FC; #100;
A = 16'h002D; B = 16'h00FD; #100;
A = 16'h002D; B = 16'h00FE; #100;
A = 16'h002D; B = 16'h00FF; #100;
A = 16'h002E; B = 16'h000; #100;
A = 16'h002E; B = 16'h001; #100;
A = 16'h002E; B = 16'h002; #100;
A = 16'h002E; B = 16'h003; #100;
A = 16'h002E; B = 16'h004; #100;
A = 16'h002E; B = 16'h005; #100;
A = 16'h002E; B = 16'h006; #100;
A = 16'h002E; B = 16'h007; #100;
A = 16'h002E; B = 16'h008; #100;
A = 16'h002E; B = 16'h009; #100;
A = 16'h002E; B = 16'h00A; #100;
A = 16'h002E; B = 16'h00B; #100;
A = 16'h002E; B = 16'h00C; #100;
A = 16'h002E; B = 16'h00D; #100;
A = 16'h002E; B = 16'h00E; #100;
A = 16'h002E; B = 16'h00F; #100;
A = 16'h002E; B = 16'h0010; #100;
A = 16'h002E; B = 16'h0011; #100;
A = 16'h002E; B = 16'h0012; #100;
A = 16'h002E; B = 16'h0013; #100;
A = 16'h002E; B = 16'h0014; #100;
A = 16'h002E; B = 16'h0015; #100;
A = 16'h002E; B = 16'h0016; #100;
A = 16'h002E; B = 16'h0017; #100;
A = 16'h002E; B = 16'h0018; #100;
A = 16'h002E; B = 16'h0019; #100;
A = 16'h002E; B = 16'h001A; #100;
A = 16'h002E; B = 16'h001B; #100;
A = 16'h002E; B = 16'h001C; #100;
A = 16'h002E; B = 16'h001D; #100;
A = 16'h002E; B = 16'h001E; #100;
A = 16'h002E; B = 16'h001F; #100;
A = 16'h002E; B = 16'h0020; #100;
A = 16'h002E; B = 16'h0021; #100;
A = 16'h002E; B = 16'h0022; #100;
A = 16'h002E; B = 16'h0023; #100;
A = 16'h002E; B = 16'h0024; #100;
A = 16'h002E; B = 16'h0025; #100;
A = 16'h002E; B = 16'h0026; #100;
A = 16'h002E; B = 16'h0027; #100;
A = 16'h002E; B = 16'h0028; #100;
A = 16'h002E; B = 16'h0029; #100;
A = 16'h002E; B = 16'h002A; #100;
A = 16'h002E; B = 16'h002B; #100;
A = 16'h002E; B = 16'h002C; #100;
A = 16'h002E; B = 16'h002D; #100;
A = 16'h002E; B = 16'h002E; #100;
A = 16'h002E; B = 16'h002F; #100;
A = 16'h002E; B = 16'h0030; #100;
A = 16'h002E; B = 16'h0031; #100;
A = 16'h002E; B = 16'h0032; #100;
A = 16'h002E; B = 16'h0033; #100;
A = 16'h002E; B = 16'h0034; #100;
A = 16'h002E; B = 16'h0035; #100;
A = 16'h002E; B = 16'h0036; #100;
A = 16'h002E; B = 16'h0037; #100;
A = 16'h002E; B = 16'h0038; #100;
A = 16'h002E; B = 16'h0039; #100;
A = 16'h002E; B = 16'h003A; #100;
A = 16'h002E; B = 16'h003B; #100;
A = 16'h002E; B = 16'h003C; #100;
A = 16'h002E; B = 16'h003D; #100;
A = 16'h002E; B = 16'h003E; #100;
A = 16'h002E; B = 16'h003F; #100;
A = 16'h002E; B = 16'h0040; #100;
A = 16'h002E; B = 16'h0041; #100;
A = 16'h002E; B = 16'h0042; #100;
A = 16'h002E; B = 16'h0043; #100;
A = 16'h002E; B = 16'h0044; #100;
A = 16'h002E; B = 16'h0045; #100;
A = 16'h002E; B = 16'h0046; #100;
A = 16'h002E; B = 16'h0047; #100;
A = 16'h002E; B = 16'h0048; #100;
A = 16'h002E; B = 16'h0049; #100;
A = 16'h002E; B = 16'h004A; #100;
A = 16'h002E; B = 16'h004B; #100;
A = 16'h002E; B = 16'h004C; #100;
A = 16'h002E; B = 16'h004D; #100;
A = 16'h002E; B = 16'h004E; #100;
A = 16'h002E; B = 16'h004F; #100;
A = 16'h002E; B = 16'h0050; #100;
A = 16'h002E; B = 16'h0051; #100;
A = 16'h002E; B = 16'h0052; #100;
A = 16'h002E; B = 16'h0053; #100;
A = 16'h002E; B = 16'h0054; #100;
A = 16'h002E; B = 16'h0055; #100;
A = 16'h002E; B = 16'h0056; #100;
A = 16'h002E; B = 16'h0057; #100;
A = 16'h002E; B = 16'h0058; #100;
A = 16'h002E; B = 16'h0059; #100;
A = 16'h002E; B = 16'h005A; #100;
A = 16'h002E; B = 16'h005B; #100;
A = 16'h002E; B = 16'h005C; #100;
A = 16'h002E; B = 16'h005D; #100;
A = 16'h002E; B = 16'h005E; #100;
A = 16'h002E; B = 16'h005F; #100;
A = 16'h002E; B = 16'h0060; #100;
A = 16'h002E; B = 16'h0061; #100;
A = 16'h002E; B = 16'h0062; #100;
A = 16'h002E; B = 16'h0063; #100;
A = 16'h002E; B = 16'h0064; #100;
A = 16'h002E; B = 16'h0065; #100;
A = 16'h002E; B = 16'h0066; #100;
A = 16'h002E; B = 16'h0067; #100;
A = 16'h002E; B = 16'h0068; #100;
A = 16'h002E; B = 16'h0069; #100;
A = 16'h002E; B = 16'h006A; #100;
A = 16'h002E; B = 16'h006B; #100;
A = 16'h002E; B = 16'h006C; #100;
A = 16'h002E; B = 16'h006D; #100;
A = 16'h002E; B = 16'h006E; #100;
A = 16'h002E; B = 16'h006F; #100;
A = 16'h002E; B = 16'h0070; #100;
A = 16'h002E; B = 16'h0071; #100;
A = 16'h002E; B = 16'h0072; #100;
A = 16'h002E; B = 16'h0073; #100;
A = 16'h002E; B = 16'h0074; #100;
A = 16'h002E; B = 16'h0075; #100;
A = 16'h002E; B = 16'h0076; #100;
A = 16'h002E; B = 16'h0077; #100;
A = 16'h002E; B = 16'h0078; #100;
A = 16'h002E; B = 16'h0079; #100;
A = 16'h002E; B = 16'h007A; #100;
A = 16'h002E; B = 16'h007B; #100;
A = 16'h002E; B = 16'h007C; #100;
A = 16'h002E; B = 16'h007D; #100;
A = 16'h002E; B = 16'h007E; #100;
A = 16'h002E; B = 16'h007F; #100;
A = 16'h002E; B = 16'h0080; #100;
A = 16'h002E; B = 16'h0081; #100;
A = 16'h002E; B = 16'h0082; #100;
A = 16'h002E; B = 16'h0083; #100;
A = 16'h002E; B = 16'h0084; #100;
A = 16'h002E; B = 16'h0085; #100;
A = 16'h002E; B = 16'h0086; #100;
A = 16'h002E; B = 16'h0087; #100;
A = 16'h002E; B = 16'h0088; #100;
A = 16'h002E; B = 16'h0089; #100;
A = 16'h002E; B = 16'h008A; #100;
A = 16'h002E; B = 16'h008B; #100;
A = 16'h002E; B = 16'h008C; #100;
A = 16'h002E; B = 16'h008D; #100;
A = 16'h002E; B = 16'h008E; #100;
A = 16'h002E; B = 16'h008F; #100;
A = 16'h002E; B = 16'h0090; #100;
A = 16'h002E; B = 16'h0091; #100;
A = 16'h002E; B = 16'h0092; #100;
A = 16'h002E; B = 16'h0093; #100;
A = 16'h002E; B = 16'h0094; #100;
A = 16'h002E; B = 16'h0095; #100;
A = 16'h002E; B = 16'h0096; #100;
A = 16'h002E; B = 16'h0097; #100;
A = 16'h002E; B = 16'h0098; #100;
A = 16'h002E; B = 16'h0099; #100;
A = 16'h002E; B = 16'h009A; #100;
A = 16'h002E; B = 16'h009B; #100;
A = 16'h002E; B = 16'h009C; #100;
A = 16'h002E; B = 16'h009D; #100;
A = 16'h002E; B = 16'h009E; #100;
A = 16'h002E; B = 16'h009F; #100;
A = 16'h002E; B = 16'h00A0; #100;
A = 16'h002E; B = 16'h00A1; #100;
A = 16'h002E; B = 16'h00A2; #100;
A = 16'h002E; B = 16'h00A3; #100;
A = 16'h002E; B = 16'h00A4; #100;
A = 16'h002E; B = 16'h00A5; #100;
A = 16'h002E; B = 16'h00A6; #100;
A = 16'h002E; B = 16'h00A7; #100;
A = 16'h002E; B = 16'h00A8; #100;
A = 16'h002E; B = 16'h00A9; #100;
A = 16'h002E; B = 16'h00AA; #100;
A = 16'h002E; B = 16'h00AB; #100;
A = 16'h002E; B = 16'h00AC; #100;
A = 16'h002E; B = 16'h00AD; #100;
A = 16'h002E; B = 16'h00AE; #100;
A = 16'h002E; B = 16'h00AF; #100;
A = 16'h002E; B = 16'h00B0; #100;
A = 16'h002E; B = 16'h00B1; #100;
A = 16'h002E; B = 16'h00B2; #100;
A = 16'h002E; B = 16'h00B3; #100;
A = 16'h002E; B = 16'h00B4; #100;
A = 16'h002E; B = 16'h00B5; #100;
A = 16'h002E; B = 16'h00B6; #100;
A = 16'h002E; B = 16'h00B7; #100;
A = 16'h002E; B = 16'h00B8; #100;
A = 16'h002E; B = 16'h00B9; #100;
A = 16'h002E; B = 16'h00BA; #100;
A = 16'h002E; B = 16'h00BB; #100;
A = 16'h002E; B = 16'h00BC; #100;
A = 16'h002E; B = 16'h00BD; #100;
A = 16'h002E; B = 16'h00BE; #100;
A = 16'h002E; B = 16'h00BF; #100;
A = 16'h002E; B = 16'h00C0; #100;
A = 16'h002E; B = 16'h00C1; #100;
A = 16'h002E; B = 16'h00C2; #100;
A = 16'h002E; B = 16'h00C3; #100;
A = 16'h002E; B = 16'h00C4; #100;
A = 16'h002E; B = 16'h00C5; #100;
A = 16'h002E; B = 16'h00C6; #100;
A = 16'h002E; B = 16'h00C7; #100;
A = 16'h002E; B = 16'h00C8; #100;
A = 16'h002E; B = 16'h00C9; #100;
A = 16'h002E; B = 16'h00CA; #100;
A = 16'h002E; B = 16'h00CB; #100;
A = 16'h002E; B = 16'h00CC; #100;
A = 16'h002E; B = 16'h00CD; #100;
A = 16'h002E; B = 16'h00CE; #100;
A = 16'h002E; B = 16'h00CF; #100;
A = 16'h002E; B = 16'h00D0; #100;
A = 16'h002E; B = 16'h00D1; #100;
A = 16'h002E; B = 16'h00D2; #100;
A = 16'h002E; B = 16'h00D3; #100;
A = 16'h002E; B = 16'h00D4; #100;
A = 16'h002E; B = 16'h00D5; #100;
A = 16'h002E; B = 16'h00D6; #100;
A = 16'h002E; B = 16'h00D7; #100;
A = 16'h002E; B = 16'h00D8; #100;
A = 16'h002E; B = 16'h00D9; #100;
A = 16'h002E; B = 16'h00DA; #100;
A = 16'h002E; B = 16'h00DB; #100;
A = 16'h002E; B = 16'h00DC; #100;
A = 16'h002E; B = 16'h00DD; #100;
A = 16'h002E; B = 16'h00DE; #100;
A = 16'h002E; B = 16'h00DF; #100;
A = 16'h002E; B = 16'h00E0; #100;
A = 16'h002E; B = 16'h00E1; #100;
A = 16'h002E; B = 16'h00E2; #100;
A = 16'h002E; B = 16'h00E3; #100;
A = 16'h002E; B = 16'h00E4; #100;
A = 16'h002E; B = 16'h00E5; #100;
A = 16'h002E; B = 16'h00E6; #100;
A = 16'h002E; B = 16'h00E7; #100;
A = 16'h002E; B = 16'h00E8; #100;
A = 16'h002E; B = 16'h00E9; #100;
A = 16'h002E; B = 16'h00EA; #100;
A = 16'h002E; B = 16'h00EB; #100;
A = 16'h002E; B = 16'h00EC; #100;
A = 16'h002E; B = 16'h00ED; #100;
A = 16'h002E; B = 16'h00EE; #100;
A = 16'h002E; B = 16'h00EF; #100;
A = 16'h002E; B = 16'h00F0; #100;
A = 16'h002E; B = 16'h00F1; #100;
A = 16'h002E; B = 16'h00F2; #100;
A = 16'h002E; B = 16'h00F3; #100;
A = 16'h002E; B = 16'h00F4; #100;
A = 16'h002E; B = 16'h00F5; #100;
A = 16'h002E; B = 16'h00F6; #100;
A = 16'h002E; B = 16'h00F7; #100;
A = 16'h002E; B = 16'h00F8; #100;
A = 16'h002E; B = 16'h00F9; #100;
A = 16'h002E; B = 16'h00FA; #100;
A = 16'h002E; B = 16'h00FB; #100;
A = 16'h002E; B = 16'h00FC; #100;
A = 16'h002E; B = 16'h00FD; #100;
A = 16'h002E; B = 16'h00FE; #100;
A = 16'h002E; B = 16'h00FF; #100;
A = 16'h002F; B = 16'h000; #100;
A = 16'h002F; B = 16'h001; #100;
A = 16'h002F; B = 16'h002; #100;
A = 16'h002F; B = 16'h003; #100;
A = 16'h002F; B = 16'h004; #100;
A = 16'h002F; B = 16'h005; #100;
A = 16'h002F; B = 16'h006; #100;
A = 16'h002F; B = 16'h007; #100;
A = 16'h002F; B = 16'h008; #100;
A = 16'h002F; B = 16'h009; #100;
A = 16'h002F; B = 16'h00A; #100;
A = 16'h002F; B = 16'h00B; #100;
A = 16'h002F; B = 16'h00C; #100;
A = 16'h002F; B = 16'h00D; #100;
A = 16'h002F; B = 16'h00E; #100;
A = 16'h002F; B = 16'h00F; #100;
A = 16'h002F; B = 16'h0010; #100;
A = 16'h002F; B = 16'h0011; #100;
A = 16'h002F; B = 16'h0012; #100;
A = 16'h002F; B = 16'h0013; #100;
A = 16'h002F; B = 16'h0014; #100;
A = 16'h002F; B = 16'h0015; #100;
A = 16'h002F; B = 16'h0016; #100;
A = 16'h002F; B = 16'h0017; #100;
A = 16'h002F; B = 16'h0018; #100;
A = 16'h002F; B = 16'h0019; #100;
A = 16'h002F; B = 16'h001A; #100;
A = 16'h002F; B = 16'h001B; #100;
A = 16'h002F; B = 16'h001C; #100;
A = 16'h002F; B = 16'h001D; #100;
A = 16'h002F; B = 16'h001E; #100;
A = 16'h002F; B = 16'h001F; #100;
A = 16'h002F; B = 16'h0020; #100;
A = 16'h002F; B = 16'h0021; #100;
A = 16'h002F; B = 16'h0022; #100;
A = 16'h002F; B = 16'h0023; #100;
A = 16'h002F; B = 16'h0024; #100;
A = 16'h002F; B = 16'h0025; #100;
A = 16'h002F; B = 16'h0026; #100;
A = 16'h002F; B = 16'h0027; #100;
A = 16'h002F; B = 16'h0028; #100;
A = 16'h002F; B = 16'h0029; #100;
A = 16'h002F; B = 16'h002A; #100;
A = 16'h002F; B = 16'h002B; #100;
A = 16'h002F; B = 16'h002C; #100;
A = 16'h002F; B = 16'h002D; #100;
A = 16'h002F; B = 16'h002E; #100;
A = 16'h002F; B = 16'h002F; #100;
A = 16'h002F; B = 16'h0030; #100;
A = 16'h002F; B = 16'h0031; #100;
A = 16'h002F; B = 16'h0032; #100;
A = 16'h002F; B = 16'h0033; #100;
A = 16'h002F; B = 16'h0034; #100;
A = 16'h002F; B = 16'h0035; #100;
A = 16'h002F; B = 16'h0036; #100;
A = 16'h002F; B = 16'h0037; #100;
A = 16'h002F; B = 16'h0038; #100;
A = 16'h002F; B = 16'h0039; #100;
A = 16'h002F; B = 16'h003A; #100;
A = 16'h002F; B = 16'h003B; #100;
A = 16'h002F; B = 16'h003C; #100;
A = 16'h002F; B = 16'h003D; #100;
A = 16'h002F; B = 16'h003E; #100;
A = 16'h002F; B = 16'h003F; #100;
A = 16'h002F; B = 16'h0040; #100;
A = 16'h002F; B = 16'h0041; #100;
A = 16'h002F; B = 16'h0042; #100;
A = 16'h002F; B = 16'h0043; #100;
A = 16'h002F; B = 16'h0044; #100;
A = 16'h002F; B = 16'h0045; #100;
A = 16'h002F; B = 16'h0046; #100;
A = 16'h002F; B = 16'h0047; #100;
A = 16'h002F; B = 16'h0048; #100;
A = 16'h002F; B = 16'h0049; #100;
A = 16'h002F; B = 16'h004A; #100;
A = 16'h002F; B = 16'h004B; #100;
A = 16'h002F; B = 16'h004C; #100;
A = 16'h002F; B = 16'h004D; #100;
A = 16'h002F; B = 16'h004E; #100;
A = 16'h002F; B = 16'h004F; #100;
A = 16'h002F; B = 16'h0050; #100;
A = 16'h002F; B = 16'h0051; #100;
A = 16'h002F; B = 16'h0052; #100;
A = 16'h002F; B = 16'h0053; #100;
A = 16'h002F; B = 16'h0054; #100;
A = 16'h002F; B = 16'h0055; #100;
A = 16'h002F; B = 16'h0056; #100;
A = 16'h002F; B = 16'h0057; #100;
A = 16'h002F; B = 16'h0058; #100;
A = 16'h002F; B = 16'h0059; #100;
A = 16'h002F; B = 16'h005A; #100;
A = 16'h002F; B = 16'h005B; #100;
A = 16'h002F; B = 16'h005C; #100;
A = 16'h002F; B = 16'h005D; #100;
A = 16'h002F; B = 16'h005E; #100;
A = 16'h002F; B = 16'h005F; #100;
A = 16'h002F; B = 16'h0060; #100;
A = 16'h002F; B = 16'h0061; #100;
A = 16'h002F; B = 16'h0062; #100;
A = 16'h002F; B = 16'h0063; #100;
A = 16'h002F; B = 16'h0064; #100;
A = 16'h002F; B = 16'h0065; #100;
A = 16'h002F; B = 16'h0066; #100;
A = 16'h002F; B = 16'h0067; #100;
A = 16'h002F; B = 16'h0068; #100;
A = 16'h002F; B = 16'h0069; #100;
A = 16'h002F; B = 16'h006A; #100;
A = 16'h002F; B = 16'h006B; #100;
A = 16'h002F; B = 16'h006C; #100;
A = 16'h002F; B = 16'h006D; #100;
A = 16'h002F; B = 16'h006E; #100;
A = 16'h002F; B = 16'h006F; #100;
A = 16'h002F; B = 16'h0070; #100;
A = 16'h002F; B = 16'h0071; #100;
A = 16'h002F; B = 16'h0072; #100;
A = 16'h002F; B = 16'h0073; #100;
A = 16'h002F; B = 16'h0074; #100;
A = 16'h002F; B = 16'h0075; #100;
A = 16'h002F; B = 16'h0076; #100;
A = 16'h002F; B = 16'h0077; #100;
A = 16'h002F; B = 16'h0078; #100;
A = 16'h002F; B = 16'h0079; #100;
A = 16'h002F; B = 16'h007A; #100;
A = 16'h002F; B = 16'h007B; #100;
A = 16'h002F; B = 16'h007C; #100;
A = 16'h002F; B = 16'h007D; #100;
A = 16'h002F; B = 16'h007E; #100;
A = 16'h002F; B = 16'h007F; #100;
A = 16'h002F; B = 16'h0080; #100;
A = 16'h002F; B = 16'h0081; #100;
A = 16'h002F; B = 16'h0082; #100;
A = 16'h002F; B = 16'h0083; #100;
A = 16'h002F; B = 16'h0084; #100;
A = 16'h002F; B = 16'h0085; #100;
A = 16'h002F; B = 16'h0086; #100;
A = 16'h002F; B = 16'h0087; #100;
A = 16'h002F; B = 16'h0088; #100;
A = 16'h002F; B = 16'h0089; #100;
A = 16'h002F; B = 16'h008A; #100;
A = 16'h002F; B = 16'h008B; #100;
A = 16'h002F; B = 16'h008C; #100;
A = 16'h002F; B = 16'h008D; #100;
A = 16'h002F; B = 16'h008E; #100;
A = 16'h002F; B = 16'h008F; #100;
A = 16'h002F; B = 16'h0090; #100;
A = 16'h002F; B = 16'h0091; #100;
A = 16'h002F; B = 16'h0092; #100;
A = 16'h002F; B = 16'h0093; #100;
A = 16'h002F; B = 16'h0094; #100;
A = 16'h002F; B = 16'h0095; #100;
A = 16'h002F; B = 16'h0096; #100;
A = 16'h002F; B = 16'h0097; #100;
A = 16'h002F; B = 16'h0098; #100;
A = 16'h002F; B = 16'h0099; #100;
A = 16'h002F; B = 16'h009A; #100;
A = 16'h002F; B = 16'h009B; #100;
A = 16'h002F; B = 16'h009C; #100;
A = 16'h002F; B = 16'h009D; #100;
A = 16'h002F; B = 16'h009E; #100;
A = 16'h002F; B = 16'h009F; #100;
A = 16'h002F; B = 16'h00A0; #100;
A = 16'h002F; B = 16'h00A1; #100;
A = 16'h002F; B = 16'h00A2; #100;
A = 16'h002F; B = 16'h00A3; #100;
A = 16'h002F; B = 16'h00A4; #100;
A = 16'h002F; B = 16'h00A5; #100;
A = 16'h002F; B = 16'h00A6; #100;
A = 16'h002F; B = 16'h00A7; #100;
A = 16'h002F; B = 16'h00A8; #100;
A = 16'h002F; B = 16'h00A9; #100;
A = 16'h002F; B = 16'h00AA; #100;
A = 16'h002F; B = 16'h00AB; #100;
A = 16'h002F; B = 16'h00AC; #100;
A = 16'h002F; B = 16'h00AD; #100;
A = 16'h002F; B = 16'h00AE; #100;
A = 16'h002F; B = 16'h00AF; #100;
A = 16'h002F; B = 16'h00B0; #100;
A = 16'h002F; B = 16'h00B1; #100;
A = 16'h002F; B = 16'h00B2; #100;
A = 16'h002F; B = 16'h00B3; #100;
A = 16'h002F; B = 16'h00B4; #100;
A = 16'h002F; B = 16'h00B5; #100;
A = 16'h002F; B = 16'h00B6; #100;
A = 16'h002F; B = 16'h00B7; #100;
A = 16'h002F; B = 16'h00B8; #100;
A = 16'h002F; B = 16'h00B9; #100;
A = 16'h002F; B = 16'h00BA; #100;
A = 16'h002F; B = 16'h00BB; #100;
A = 16'h002F; B = 16'h00BC; #100;
A = 16'h002F; B = 16'h00BD; #100;
A = 16'h002F; B = 16'h00BE; #100;
A = 16'h002F; B = 16'h00BF; #100;
A = 16'h002F; B = 16'h00C0; #100;
A = 16'h002F; B = 16'h00C1; #100;
A = 16'h002F; B = 16'h00C2; #100;
A = 16'h002F; B = 16'h00C3; #100;
A = 16'h002F; B = 16'h00C4; #100;
A = 16'h002F; B = 16'h00C5; #100;
A = 16'h002F; B = 16'h00C6; #100;
A = 16'h002F; B = 16'h00C7; #100;
A = 16'h002F; B = 16'h00C8; #100;
A = 16'h002F; B = 16'h00C9; #100;
A = 16'h002F; B = 16'h00CA; #100;
A = 16'h002F; B = 16'h00CB; #100;
A = 16'h002F; B = 16'h00CC; #100;
A = 16'h002F; B = 16'h00CD; #100;
A = 16'h002F; B = 16'h00CE; #100;
A = 16'h002F; B = 16'h00CF; #100;
A = 16'h002F; B = 16'h00D0; #100;
A = 16'h002F; B = 16'h00D1; #100;
A = 16'h002F; B = 16'h00D2; #100;
A = 16'h002F; B = 16'h00D3; #100;
A = 16'h002F; B = 16'h00D4; #100;
A = 16'h002F; B = 16'h00D5; #100;
A = 16'h002F; B = 16'h00D6; #100;
A = 16'h002F; B = 16'h00D7; #100;
A = 16'h002F; B = 16'h00D8; #100;
A = 16'h002F; B = 16'h00D9; #100;
A = 16'h002F; B = 16'h00DA; #100;
A = 16'h002F; B = 16'h00DB; #100;
A = 16'h002F; B = 16'h00DC; #100;
A = 16'h002F; B = 16'h00DD; #100;
A = 16'h002F; B = 16'h00DE; #100;
A = 16'h002F; B = 16'h00DF; #100;
A = 16'h002F; B = 16'h00E0; #100;
A = 16'h002F; B = 16'h00E1; #100;
A = 16'h002F; B = 16'h00E2; #100;
A = 16'h002F; B = 16'h00E3; #100;
A = 16'h002F; B = 16'h00E4; #100;
A = 16'h002F; B = 16'h00E5; #100;
A = 16'h002F; B = 16'h00E6; #100;
A = 16'h002F; B = 16'h00E7; #100;
A = 16'h002F; B = 16'h00E8; #100;
A = 16'h002F; B = 16'h00E9; #100;
A = 16'h002F; B = 16'h00EA; #100;
A = 16'h002F; B = 16'h00EB; #100;
A = 16'h002F; B = 16'h00EC; #100;
A = 16'h002F; B = 16'h00ED; #100;
A = 16'h002F; B = 16'h00EE; #100;
A = 16'h002F; B = 16'h00EF; #100;
A = 16'h002F; B = 16'h00F0; #100;
A = 16'h002F; B = 16'h00F1; #100;
A = 16'h002F; B = 16'h00F2; #100;
A = 16'h002F; B = 16'h00F3; #100;
A = 16'h002F; B = 16'h00F4; #100;
A = 16'h002F; B = 16'h00F5; #100;
A = 16'h002F; B = 16'h00F6; #100;
A = 16'h002F; B = 16'h00F7; #100;
A = 16'h002F; B = 16'h00F8; #100;
A = 16'h002F; B = 16'h00F9; #100;
A = 16'h002F; B = 16'h00FA; #100;
A = 16'h002F; B = 16'h00FB; #100;
A = 16'h002F; B = 16'h00FC; #100;
A = 16'h002F; B = 16'h00FD; #100;
A = 16'h002F; B = 16'h00FE; #100;
A = 16'h002F; B = 16'h00FF; #100;
A = 16'h0030; B = 16'h000; #100;
A = 16'h0030; B = 16'h001; #100;
A = 16'h0030; B = 16'h002; #100;
A = 16'h0030; B = 16'h003; #100;
A = 16'h0030; B = 16'h004; #100;
A = 16'h0030; B = 16'h005; #100;
A = 16'h0030; B = 16'h006; #100;
A = 16'h0030; B = 16'h007; #100;
A = 16'h0030; B = 16'h008; #100;
A = 16'h0030; B = 16'h009; #100;
A = 16'h0030; B = 16'h00A; #100;
A = 16'h0030; B = 16'h00B; #100;
A = 16'h0030; B = 16'h00C; #100;
A = 16'h0030; B = 16'h00D; #100;
A = 16'h0030; B = 16'h00E; #100;
A = 16'h0030; B = 16'h00F; #100;
A = 16'h0030; B = 16'h0010; #100;
A = 16'h0030; B = 16'h0011; #100;
A = 16'h0030; B = 16'h0012; #100;
A = 16'h0030; B = 16'h0013; #100;
A = 16'h0030; B = 16'h0014; #100;
A = 16'h0030; B = 16'h0015; #100;
A = 16'h0030; B = 16'h0016; #100;
A = 16'h0030; B = 16'h0017; #100;
A = 16'h0030; B = 16'h0018; #100;
A = 16'h0030; B = 16'h0019; #100;
A = 16'h0030; B = 16'h001A; #100;
A = 16'h0030; B = 16'h001B; #100;
A = 16'h0030; B = 16'h001C; #100;
A = 16'h0030; B = 16'h001D; #100;
A = 16'h0030; B = 16'h001E; #100;
A = 16'h0030; B = 16'h001F; #100;
A = 16'h0030; B = 16'h0020; #100;
A = 16'h0030; B = 16'h0021; #100;
A = 16'h0030; B = 16'h0022; #100;
A = 16'h0030; B = 16'h0023; #100;
A = 16'h0030; B = 16'h0024; #100;
A = 16'h0030; B = 16'h0025; #100;
A = 16'h0030; B = 16'h0026; #100;
A = 16'h0030; B = 16'h0027; #100;
A = 16'h0030; B = 16'h0028; #100;
A = 16'h0030; B = 16'h0029; #100;
A = 16'h0030; B = 16'h002A; #100;
A = 16'h0030; B = 16'h002B; #100;
A = 16'h0030; B = 16'h002C; #100;
A = 16'h0030; B = 16'h002D; #100;
A = 16'h0030; B = 16'h002E; #100;
A = 16'h0030; B = 16'h002F; #100;
A = 16'h0030; B = 16'h0030; #100;
A = 16'h0030; B = 16'h0031; #100;
A = 16'h0030; B = 16'h0032; #100;
A = 16'h0030; B = 16'h0033; #100;
A = 16'h0030; B = 16'h0034; #100;
A = 16'h0030; B = 16'h0035; #100;
A = 16'h0030; B = 16'h0036; #100;
A = 16'h0030; B = 16'h0037; #100;
A = 16'h0030; B = 16'h0038; #100;
A = 16'h0030; B = 16'h0039; #100;
A = 16'h0030; B = 16'h003A; #100;
A = 16'h0030; B = 16'h003B; #100;
A = 16'h0030; B = 16'h003C; #100;
A = 16'h0030; B = 16'h003D; #100;
A = 16'h0030; B = 16'h003E; #100;
A = 16'h0030; B = 16'h003F; #100;
A = 16'h0030; B = 16'h0040; #100;
A = 16'h0030; B = 16'h0041; #100;
A = 16'h0030; B = 16'h0042; #100;
A = 16'h0030; B = 16'h0043; #100;
A = 16'h0030; B = 16'h0044; #100;
A = 16'h0030; B = 16'h0045; #100;
A = 16'h0030; B = 16'h0046; #100;
A = 16'h0030; B = 16'h0047; #100;
A = 16'h0030; B = 16'h0048; #100;
A = 16'h0030; B = 16'h0049; #100;
A = 16'h0030; B = 16'h004A; #100;
A = 16'h0030; B = 16'h004B; #100;
A = 16'h0030; B = 16'h004C; #100;
A = 16'h0030; B = 16'h004D; #100;
A = 16'h0030; B = 16'h004E; #100;
A = 16'h0030; B = 16'h004F; #100;
A = 16'h0030; B = 16'h0050; #100;
A = 16'h0030; B = 16'h0051; #100;
A = 16'h0030; B = 16'h0052; #100;
A = 16'h0030; B = 16'h0053; #100;
A = 16'h0030; B = 16'h0054; #100;
A = 16'h0030; B = 16'h0055; #100;
A = 16'h0030; B = 16'h0056; #100;
A = 16'h0030; B = 16'h0057; #100;
A = 16'h0030; B = 16'h0058; #100;
A = 16'h0030; B = 16'h0059; #100;
A = 16'h0030; B = 16'h005A; #100;
A = 16'h0030; B = 16'h005B; #100;
A = 16'h0030; B = 16'h005C; #100;
A = 16'h0030; B = 16'h005D; #100;
A = 16'h0030; B = 16'h005E; #100;
A = 16'h0030; B = 16'h005F; #100;
A = 16'h0030; B = 16'h0060; #100;
A = 16'h0030; B = 16'h0061; #100;
A = 16'h0030; B = 16'h0062; #100;
A = 16'h0030; B = 16'h0063; #100;
A = 16'h0030; B = 16'h0064; #100;
A = 16'h0030; B = 16'h0065; #100;
A = 16'h0030; B = 16'h0066; #100;
A = 16'h0030; B = 16'h0067; #100;
A = 16'h0030; B = 16'h0068; #100;
A = 16'h0030; B = 16'h0069; #100;
A = 16'h0030; B = 16'h006A; #100;
A = 16'h0030; B = 16'h006B; #100;
A = 16'h0030; B = 16'h006C; #100;
A = 16'h0030; B = 16'h006D; #100;
A = 16'h0030; B = 16'h006E; #100;
A = 16'h0030; B = 16'h006F; #100;
A = 16'h0030; B = 16'h0070; #100;
A = 16'h0030; B = 16'h0071; #100;
A = 16'h0030; B = 16'h0072; #100;
A = 16'h0030; B = 16'h0073; #100;
A = 16'h0030; B = 16'h0074; #100;
A = 16'h0030; B = 16'h0075; #100;
A = 16'h0030; B = 16'h0076; #100;
A = 16'h0030; B = 16'h0077; #100;
A = 16'h0030; B = 16'h0078; #100;
A = 16'h0030; B = 16'h0079; #100;
A = 16'h0030; B = 16'h007A; #100;
A = 16'h0030; B = 16'h007B; #100;
A = 16'h0030; B = 16'h007C; #100;
A = 16'h0030; B = 16'h007D; #100;
A = 16'h0030; B = 16'h007E; #100;
A = 16'h0030; B = 16'h007F; #100;
A = 16'h0030; B = 16'h0080; #100;
A = 16'h0030; B = 16'h0081; #100;
A = 16'h0030; B = 16'h0082; #100;
A = 16'h0030; B = 16'h0083; #100;
A = 16'h0030; B = 16'h0084; #100;
A = 16'h0030; B = 16'h0085; #100;
A = 16'h0030; B = 16'h0086; #100;
A = 16'h0030; B = 16'h0087; #100;
A = 16'h0030; B = 16'h0088; #100;
A = 16'h0030; B = 16'h0089; #100;
A = 16'h0030; B = 16'h008A; #100;
A = 16'h0030; B = 16'h008B; #100;
A = 16'h0030; B = 16'h008C; #100;
A = 16'h0030; B = 16'h008D; #100;
A = 16'h0030; B = 16'h008E; #100;
A = 16'h0030; B = 16'h008F; #100;
A = 16'h0030; B = 16'h0090; #100;
A = 16'h0030; B = 16'h0091; #100;
A = 16'h0030; B = 16'h0092; #100;
A = 16'h0030; B = 16'h0093; #100;
A = 16'h0030; B = 16'h0094; #100;
A = 16'h0030; B = 16'h0095; #100;
A = 16'h0030; B = 16'h0096; #100;
A = 16'h0030; B = 16'h0097; #100;
A = 16'h0030; B = 16'h0098; #100;
A = 16'h0030; B = 16'h0099; #100;
A = 16'h0030; B = 16'h009A; #100;
A = 16'h0030; B = 16'h009B; #100;
A = 16'h0030; B = 16'h009C; #100;
A = 16'h0030; B = 16'h009D; #100;
A = 16'h0030; B = 16'h009E; #100;
A = 16'h0030; B = 16'h009F; #100;
A = 16'h0030; B = 16'h00A0; #100;
A = 16'h0030; B = 16'h00A1; #100;
A = 16'h0030; B = 16'h00A2; #100;
A = 16'h0030; B = 16'h00A3; #100;
A = 16'h0030; B = 16'h00A4; #100;
A = 16'h0030; B = 16'h00A5; #100;
A = 16'h0030; B = 16'h00A6; #100;
A = 16'h0030; B = 16'h00A7; #100;
A = 16'h0030; B = 16'h00A8; #100;
A = 16'h0030; B = 16'h00A9; #100;
A = 16'h0030; B = 16'h00AA; #100;
A = 16'h0030; B = 16'h00AB; #100;
A = 16'h0030; B = 16'h00AC; #100;
A = 16'h0030; B = 16'h00AD; #100;
A = 16'h0030; B = 16'h00AE; #100;
A = 16'h0030; B = 16'h00AF; #100;
A = 16'h0030; B = 16'h00B0; #100;
A = 16'h0030; B = 16'h00B1; #100;
A = 16'h0030; B = 16'h00B2; #100;
A = 16'h0030; B = 16'h00B3; #100;
A = 16'h0030; B = 16'h00B4; #100;
A = 16'h0030; B = 16'h00B5; #100;
A = 16'h0030; B = 16'h00B6; #100;
A = 16'h0030; B = 16'h00B7; #100;
A = 16'h0030; B = 16'h00B8; #100;
A = 16'h0030; B = 16'h00B9; #100;
A = 16'h0030; B = 16'h00BA; #100;
A = 16'h0030; B = 16'h00BB; #100;
A = 16'h0030; B = 16'h00BC; #100;
A = 16'h0030; B = 16'h00BD; #100;
A = 16'h0030; B = 16'h00BE; #100;
A = 16'h0030; B = 16'h00BF; #100;
A = 16'h0030; B = 16'h00C0; #100;
A = 16'h0030; B = 16'h00C1; #100;
A = 16'h0030; B = 16'h00C2; #100;
A = 16'h0030; B = 16'h00C3; #100;
A = 16'h0030; B = 16'h00C4; #100;
A = 16'h0030; B = 16'h00C5; #100;
A = 16'h0030; B = 16'h00C6; #100;
A = 16'h0030; B = 16'h00C7; #100;
A = 16'h0030; B = 16'h00C8; #100;
A = 16'h0030; B = 16'h00C9; #100;
A = 16'h0030; B = 16'h00CA; #100;
A = 16'h0030; B = 16'h00CB; #100;
A = 16'h0030; B = 16'h00CC; #100;
A = 16'h0030; B = 16'h00CD; #100;
A = 16'h0030; B = 16'h00CE; #100;
A = 16'h0030; B = 16'h00CF; #100;
A = 16'h0030; B = 16'h00D0; #100;
A = 16'h0030; B = 16'h00D1; #100;
A = 16'h0030; B = 16'h00D2; #100;
A = 16'h0030; B = 16'h00D3; #100;
A = 16'h0030; B = 16'h00D4; #100;
A = 16'h0030; B = 16'h00D5; #100;
A = 16'h0030; B = 16'h00D6; #100;
A = 16'h0030; B = 16'h00D7; #100;
A = 16'h0030; B = 16'h00D8; #100;
A = 16'h0030; B = 16'h00D9; #100;
A = 16'h0030; B = 16'h00DA; #100;
A = 16'h0030; B = 16'h00DB; #100;
A = 16'h0030; B = 16'h00DC; #100;
A = 16'h0030; B = 16'h00DD; #100;
A = 16'h0030; B = 16'h00DE; #100;
A = 16'h0030; B = 16'h00DF; #100;
A = 16'h0030; B = 16'h00E0; #100;
A = 16'h0030; B = 16'h00E1; #100;
A = 16'h0030; B = 16'h00E2; #100;
A = 16'h0030; B = 16'h00E3; #100;
A = 16'h0030; B = 16'h00E4; #100;
A = 16'h0030; B = 16'h00E5; #100;
A = 16'h0030; B = 16'h00E6; #100;
A = 16'h0030; B = 16'h00E7; #100;
A = 16'h0030; B = 16'h00E8; #100;
A = 16'h0030; B = 16'h00E9; #100;
A = 16'h0030; B = 16'h00EA; #100;
A = 16'h0030; B = 16'h00EB; #100;
A = 16'h0030; B = 16'h00EC; #100;
A = 16'h0030; B = 16'h00ED; #100;
A = 16'h0030; B = 16'h00EE; #100;
A = 16'h0030; B = 16'h00EF; #100;
A = 16'h0030; B = 16'h00F0; #100;
A = 16'h0030; B = 16'h00F1; #100;
A = 16'h0030; B = 16'h00F2; #100;
A = 16'h0030; B = 16'h00F3; #100;
A = 16'h0030; B = 16'h00F4; #100;
A = 16'h0030; B = 16'h00F5; #100;
A = 16'h0030; B = 16'h00F6; #100;
A = 16'h0030; B = 16'h00F7; #100;
A = 16'h0030; B = 16'h00F8; #100;
A = 16'h0030; B = 16'h00F9; #100;
A = 16'h0030; B = 16'h00FA; #100;
A = 16'h0030; B = 16'h00FB; #100;
A = 16'h0030; B = 16'h00FC; #100;
A = 16'h0030; B = 16'h00FD; #100;
A = 16'h0030; B = 16'h00FE; #100;
A = 16'h0030; B = 16'h00FF; #100;
A = 16'h0031; B = 16'h000; #100;
A = 16'h0031; B = 16'h001; #100;
A = 16'h0031; B = 16'h002; #100;
A = 16'h0031; B = 16'h003; #100;
A = 16'h0031; B = 16'h004; #100;
A = 16'h0031; B = 16'h005; #100;
A = 16'h0031; B = 16'h006; #100;
A = 16'h0031; B = 16'h007; #100;
A = 16'h0031; B = 16'h008; #100;
A = 16'h0031; B = 16'h009; #100;
A = 16'h0031; B = 16'h00A; #100;
A = 16'h0031; B = 16'h00B; #100;
A = 16'h0031; B = 16'h00C; #100;
A = 16'h0031; B = 16'h00D; #100;
A = 16'h0031; B = 16'h00E; #100;
A = 16'h0031; B = 16'h00F; #100;
A = 16'h0031; B = 16'h0010; #100;
A = 16'h0031; B = 16'h0011; #100;
A = 16'h0031; B = 16'h0012; #100;
A = 16'h0031; B = 16'h0013; #100;
A = 16'h0031; B = 16'h0014; #100;
A = 16'h0031; B = 16'h0015; #100;
A = 16'h0031; B = 16'h0016; #100;
A = 16'h0031; B = 16'h0017; #100;
A = 16'h0031; B = 16'h0018; #100;
A = 16'h0031; B = 16'h0019; #100;
A = 16'h0031; B = 16'h001A; #100;
A = 16'h0031; B = 16'h001B; #100;
A = 16'h0031; B = 16'h001C; #100;
A = 16'h0031; B = 16'h001D; #100;
A = 16'h0031; B = 16'h001E; #100;
A = 16'h0031; B = 16'h001F; #100;
A = 16'h0031; B = 16'h0020; #100;
A = 16'h0031; B = 16'h0021; #100;
A = 16'h0031; B = 16'h0022; #100;
A = 16'h0031; B = 16'h0023; #100;
A = 16'h0031; B = 16'h0024; #100;
A = 16'h0031; B = 16'h0025; #100;
A = 16'h0031; B = 16'h0026; #100;
A = 16'h0031; B = 16'h0027; #100;
A = 16'h0031; B = 16'h0028; #100;
A = 16'h0031; B = 16'h0029; #100;
A = 16'h0031; B = 16'h002A; #100;
A = 16'h0031; B = 16'h002B; #100;
A = 16'h0031; B = 16'h002C; #100;
A = 16'h0031; B = 16'h002D; #100;
A = 16'h0031; B = 16'h002E; #100;
A = 16'h0031; B = 16'h002F; #100;
A = 16'h0031; B = 16'h0030; #100;
A = 16'h0031; B = 16'h0031; #100;
A = 16'h0031; B = 16'h0032; #100;
A = 16'h0031; B = 16'h0033; #100;
A = 16'h0031; B = 16'h0034; #100;
A = 16'h0031; B = 16'h0035; #100;
A = 16'h0031; B = 16'h0036; #100;
A = 16'h0031; B = 16'h0037; #100;
A = 16'h0031; B = 16'h0038; #100;
A = 16'h0031; B = 16'h0039; #100;
A = 16'h0031; B = 16'h003A; #100;
A = 16'h0031; B = 16'h003B; #100;
A = 16'h0031; B = 16'h003C; #100;
A = 16'h0031; B = 16'h003D; #100;
A = 16'h0031; B = 16'h003E; #100;
A = 16'h0031; B = 16'h003F; #100;
A = 16'h0031; B = 16'h0040; #100;
A = 16'h0031; B = 16'h0041; #100;
A = 16'h0031; B = 16'h0042; #100;
A = 16'h0031; B = 16'h0043; #100;
A = 16'h0031; B = 16'h0044; #100;
A = 16'h0031; B = 16'h0045; #100;
A = 16'h0031; B = 16'h0046; #100;
A = 16'h0031; B = 16'h0047; #100;
A = 16'h0031; B = 16'h0048; #100;
A = 16'h0031; B = 16'h0049; #100;
A = 16'h0031; B = 16'h004A; #100;
A = 16'h0031; B = 16'h004B; #100;
A = 16'h0031; B = 16'h004C; #100;
A = 16'h0031; B = 16'h004D; #100;
A = 16'h0031; B = 16'h004E; #100;
A = 16'h0031; B = 16'h004F; #100;
A = 16'h0031; B = 16'h0050; #100;
A = 16'h0031; B = 16'h0051; #100;
A = 16'h0031; B = 16'h0052; #100;
A = 16'h0031; B = 16'h0053; #100;
A = 16'h0031; B = 16'h0054; #100;
A = 16'h0031; B = 16'h0055; #100;
A = 16'h0031; B = 16'h0056; #100;
A = 16'h0031; B = 16'h0057; #100;
A = 16'h0031; B = 16'h0058; #100;
A = 16'h0031; B = 16'h0059; #100;
A = 16'h0031; B = 16'h005A; #100;
A = 16'h0031; B = 16'h005B; #100;
A = 16'h0031; B = 16'h005C; #100;
A = 16'h0031; B = 16'h005D; #100;
A = 16'h0031; B = 16'h005E; #100;
A = 16'h0031; B = 16'h005F; #100;
A = 16'h0031; B = 16'h0060; #100;
A = 16'h0031; B = 16'h0061; #100;
A = 16'h0031; B = 16'h0062; #100;
A = 16'h0031; B = 16'h0063; #100;
A = 16'h0031; B = 16'h0064; #100;
A = 16'h0031; B = 16'h0065; #100;
A = 16'h0031; B = 16'h0066; #100;
A = 16'h0031; B = 16'h0067; #100;
A = 16'h0031; B = 16'h0068; #100;
A = 16'h0031; B = 16'h0069; #100;
A = 16'h0031; B = 16'h006A; #100;
A = 16'h0031; B = 16'h006B; #100;
A = 16'h0031; B = 16'h006C; #100;
A = 16'h0031; B = 16'h006D; #100;
A = 16'h0031; B = 16'h006E; #100;
A = 16'h0031; B = 16'h006F; #100;
A = 16'h0031; B = 16'h0070; #100;
A = 16'h0031; B = 16'h0071; #100;
A = 16'h0031; B = 16'h0072; #100;
A = 16'h0031; B = 16'h0073; #100;
A = 16'h0031; B = 16'h0074; #100;
A = 16'h0031; B = 16'h0075; #100;
A = 16'h0031; B = 16'h0076; #100;
A = 16'h0031; B = 16'h0077; #100;
A = 16'h0031; B = 16'h0078; #100;
A = 16'h0031; B = 16'h0079; #100;
A = 16'h0031; B = 16'h007A; #100;
A = 16'h0031; B = 16'h007B; #100;
A = 16'h0031; B = 16'h007C; #100;
A = 16'h0031; B = 16'h007D; #100;
A = 16'h0031; B = 16'h007E; #100;
A = 16'h0031; B = 16'h007F; #100;
A = 16'h0031; B = 16'h0080; #100;
A = 16'h0031; B = 16'h0081; #100;
A = 16'h0031; B = 16'h0082; #100;
A = 16'h0031; B = 16'h0083; #100;
A = 16'h0031; B = 16'h0084; #100;
A = 16'h0031; B = 16'h0085; #100;
A = 16'h0031; B = 16'h0086; #100;
A = 16'h0031; B = 16'h0087; #100;
A = 16'h0031; B = 16'h0088; #100;
A = 16'h0031; B = 16'h0089; #100;
A = 16'h0031; B = 16'h008A; #100;
A = 16'h0031; B = 16'h008B; #100;
A = 16'h0031; B = 16'h008C; #100;
A = 16'h0031; B = 16'h008D; #100;
A = 16'h0031; B = 16'h008E; #100;
A = 16'h0031; B = 16'h008F; #100;
A = 16'h0031; B = 16'h0090; #100;
A = 16'h0031; B = 16'h0091; #100;
A = 16'h0031; B = 16'h0092; #100;
A = 16'h0031; B = 16'h0093; #100;
A = 16'h0031; B = 16'h0094; #100;
A = 16'h0031; B = 16'h0095; #100;
A = 16'h0031; B = 16'h0096; #100;
A = 16'h0031; B = 16'h0097; #100;
A = 16'h0031; B = 16'h0098; #100;
A = 16'h0031; B = 16'h0099; #100;
A = 16'h0031; B = 16'h009A; #100;
A = 16'h0031; B = 16'h009B; #100;
A = 16'h0031; B = 16'h009C; #100;
A = 16'h0031; B = 16'h009D; #100;
A = 16'h0031; B = 16'h009E; #100;
A = 16'h0031; B = 16'h009F; #100;
A = 16'h0031; B = 16'h00A0; #100;
A = 16'h0031; B = 16'h00A1; #100;
A = 16'h0031; B = 16'h00A2; #100;
A = 16'h0031; B = 16'h00A3; #100;
A = 16'h0031; B = 16'h00A4; #100;
A = 16'h0031; B = 16'h00A5; #100;
A = 16'h0031; B = 16'h00A6; #100;
A = 16'h0031; B = 16'h00A7; #100;
A = 16'h0031; B = 16'h00A8; #100;
A = 16'h0031; B = 16'h00A9; #100;
A = 16'h0031; B = 16'h00AA; #100;
A = 16'h0031; B = 16'h00AB; #100;
A = 16'h0031; B = 16'h00AC; #100;
A = 16'h0031; B = 16'h00AD; #100;
A = 16'h0031; B = 16'h00AE; #100;
A = 16'h0031; B = 16'h00AF; #100;
A = 16'h0031; B = 16'h00B0; #100;
A = 16'h0031; B = 16'h00B1; #100;
A = 16'h0031; B = 16'h00B2; #100;
A = 16'h0031; B = 16'h00B3; #100;
A = 16'h0031; B = 16'h00B4; #100;
A = 16'h0031; B = 16'h00B5; #100;
A = 16'h0031; B = 16'h00B6; #100;
A = 16'h0031; B = 16'h00B7; #100;
A = 16'h0031; B = 16'h00B8; #100;
A = 16'h0031; B = 16'h00B9; #100;
A = 16'h0031; B = 16'h00BA; #100;
A = 16'h0031; B = 16'h00BB; #100;
A = 16'h0031; B = 16'h00BC; #100;
A = 16'h0031; B = 16'h00BD; #100;
A = 16'h0031; B = 16'h00BE; #100;
A = 16'h0031; B = 16'h00BF; #100;
A = 16'h0031; B = 16'h00C0; #100;
A = 16'h0031; B = 16'h00C1; #100;
A = 16'h0031; B = 16'h00C2; #100;
A = 16'h0031; B = 16'h00C3; #100;
A = 16'h0031; B = 16'h00C4; #100;
A = 16'h0031; B = 16'h00C5; #100;
A = 16'h0031; B = 16'h00C6; #100;
A = 16'h0031; B = 16'h00C7; #100;
A = 16'h0031; B = 16'h00C8; #100;
A = 16'h0031; B = 16'h00C9; #100;
A = 16'h0031; B = 16'h00CA; #100;
A = 16'h0031; B = 16'h00CB; #100;
A = 16'h0031; B = 16'h00CC; #100;
A = 16'h0031; B = 16'h00CD; #100;
A = 16'h0031; B = 16'h00CE; #100;
A = 16'h0031; B = 16'h00CF; #100;
A = 16'h0031; B = 16'h00D0; #100;
A = 16'h0031; B = 16'h00D1; #100;
A = 16'h0031; B = 16'h00D2; #100;
A = 16'h0031; B = 16'h00D3; #100;
A = 16'h0031; B = 16'h00D4; #100;
A = 16'h0031; B = 16'h00D5; #100;
A = 16'h0031; B = 16'h00D6; #100;
A = 16'h0031; B = 16'h00D7; #100;
A = 16'h0031; B = 16'h00D8; #100;
A = 16'h0031; B = 16'h00D9; #100;
A = 16'h0031; B = 16'h00DA; #100;
A = 16'h0031; B = 16'h00DB; #100;
A = 16'h0031; B = 16'h00DC; #100;
A = 16'h0031; B = 16'h00DD; #100;
A = 16'h0031; B = 16'h00DE; #100;
A = 16'h0031; B = 16'h00DF; #100;
A = 16'h0031; B = 16'h00E0; #100;
A = 16'h0031; B = 16'h00E1; #100;
A = 16'h0031; B = 16'h00E2; #100;
A = 16'h0031; B = 16'h00E3; #100;
A = 16'h0031; B = 16'h00E4; #100;
A = 16'h0031; B = 16'h00E5; #100;
A = 16'h0031; B = 16'h00E6; #100;
A = 16'h0031; B = 16'h00E7; #100;
A = 16'h0031; B = 16'h00E8; #100;
A = 16'h0031; B = 16'h00E9; #100;
A = 16'h0031; B = 16'h00EA; #100;
A = 16'h0031; B = 16'h00EB; #100;
A = 16'h0031; B = 16'h00EC; #100;
A = 16'h0031; B = 16'h00ED; #100;
A = 16'h0031; B = 16'h00EE; #100;
A = 16'h0031; B = 16'h00EF; #100;
A = 16'h0031; B = 16'h00F0; #100;
A = 16'h0031; B = 16'h00F1; #100;
A = 16'h0031; B = 16'h00F2; #100;
A = 16'h0031; B = 16'h00F3; #100;
A = 16'h0031; B = 16'h00F4; #100;
A = 16'h0031; B = 16'h00F5; #100;
A = 16'h0031; B = 16'h00F6; #100;
A = 16'h0031; B = 16'h00F7; #100;
A = 16'h0031; B = 16'h00F8; #100;
A = 16'h0031; B = 16'h00F9; #100;
A = 16'h0031; B = 16'h00FA; #100;
A = 16'h0031; B = 16'h00FB; #100;
A = 16'h0031; B = 16'h00FC; #100;
A = 16'h0031; B = 16'h00FD; #100;
A = 16'h0031; B = 16'h00FE; #100;
A = 16'h0031; B = 16'h00FF; #100;
A = 16'h0032; B = 16'h000; #100;
A = 16'h0032; B = 16'h001; #100;
A = 16'h0032; B = 16'h002; #100;
A = 16'h0032; B = 16'h003; #100;
A = 16'h0032; B = 16'h004; #100;
A = 16'h0032; B = 16'h005; #100;
A = 16'h0032; B = 16'h006; #100;
A = 16'h0032; B = 16'h007; #100;
A = 16'h0032; B = 16'h008; #100;
A = 16'h0032; B = 16'h009; #100;
A = 16'h0032; B = 16'h00A; #100;
A = 16'h0032; B = 16'h00B; #100;
A = 16'h0032; B = 16'h00C; #100;
A = 16'h0032; B = 16'h00D; #100;
A = 16'h0032; B = 16'h00E; #100;
A = 16'h0032; B = 16'h00F; #100;
A = 16'h0032; B = 16'h0010; #100;
A = 16'h0032; B = 16'h0011; #100;
A = 16'h0032; B = 16'h0012; #100;
A = 16'h0032; B = 16'h0013; #100;
A = 16'h0032; B = 16'h0014; #100;
A = 16'h0032; B = 16'h0015; #100;
A = 16'h0032; B = 16'h0016; #100;
A = 16'h0032; B = 16'h0017; #100;
A = 16'h0032; B = 16'h0018; #100;
A = 16'h0032; B = 16'h0019; #100;
A = 16'h0032; B = 16'h001A; #100;
A = 16'h0032; B = 16'h001B; #100;
A = 16'h0032; B = 16'h001C; #100;
A = 16'h0032; B = 16'h001D; #100;
A = 16'h0032; B = 16'h001E; #100;
A = 16'h0032; B = 16'h001F; #100;
A = 16'h0032; B = 16'h0020; #100;
A = 16'h0032; B = 16'h0021; #100;
A = 16'h0032; B = 16'h0022; #100;
A = 16'h0032; B = 16'h0023; #100;
A = 16'h0032; B = 16'h0024; #100;
A = 16'h0032; B = 16'h0025; #100;
A = 16'h0032; B = 16'h0026; #100;
A = 16'h0032; B = 16'h0027; #100;
A = 16'h0032; B = 16'h0028; #100;
A = 16'h0032; B = 16'h0029; #100;
A = 16'h0032; B = 16'h002A; #100;
A = 16'h0032; B = 16'h002B; #100;
A = 16'h0032; B = 16'h002C; #100;
A = 16'h0032; B = 16'h002D; #100;
A = 16'h0032; B = 16'h002E; #100;
A = 16'h0032; B = 16'h002F; #100;
A = 16'h0032; B = 16'h0030; #100;
A = 16'h0032; B = 16'h0031; #100;
A = 16'h0032; B = 16'h0032; #100;
A = 16'h0032; B = 16'h0033; #100;
A = 16'h0032; B = 16'h0034; #100;
A = 16'h0032; B = 16'h0035; #100;
A = 16'h0032; B = 16'h0036; #100;
A = 16'h0032; B = 16'h0037; #100;
A = 16'h0032; B = 16'h0038; #100;
A = 16'h0032; B = 16'h0039; #100;
A = 16'h0032; B = 16'h003A; #100;
A = 16'h0032; B = 16'h003B; #100;
A = 16'h0032; B = 16'h003C; #100;
A = 16'h0032; B = 16'h003D; #100;
A = 16'h0032; B = 16'h003E; #100;
A = 16'h0032; B = 16'h003F; #100;
A = 16'h0032; B = 16'h0040; #100;
A = 16'h0032; B = 16'h0041; #100;
A = 16'h0032; B = 16'h0042; #100;
A = 16'h0032; B = 16'h0043; #100;
A = 16'h0032; B = 16'h0044; #100;
A = 16'h0032; B = 16'h0045; #100;
A = 16'h0032; B = 16'h0046; #100;
A = 16'h0032; B = 16'h0047; #100;
A = 16'h0032; B = 16'h0048; #100;
A = 16'h0032; B = 16'h0049; #100;
A = 16'h0032; B = 16'h004A; #100;
A = 16'h0032; B = 16'h004B; #100;
A = 16'h0032; B = 16'h004C; #100;
A = 16'h0032; B = 16'h004D; #100;
A = 16'h0032; B = 16'h004E; #100;
A = 16'h0032; B = 16'h004F; #100;
A = 16'h0032; B = 16'h0050; #100;
A = 16'h0032; B = 16'h0051; #100;
A = 16'h0032; B = 16'h0052; #100;
A = 16'h0032; B = 16'h0053; #100;
A = 16'h0032; B = 16'h0054; #100;
A = 16'h0032; B = 16'h0055; #100;
A = 16'h0032; B = 16'h0056; #100;
A = 16'h0032; B = 16'h0057; #100;
A = 16'h0032; B = 16'h0058; #100;
A = 16'h0032; B = 16'h0059; #100;
A = 16'h0032; B = 16'h005A; #100;
A = 16'h0032; B = 16'h005B; #100;
A = 16'h0032; B = 16'h005C; #100;
A = 16'h0032; B = 16'h005D; #100;
A = 16'h0032; B = 16'h005E; #100;
A = 16'h0032; B = 16'h005F; #100;
A = 16'h0032; B = 16'h0060; #100;
A = 16'h0032; B = 16'h0061; #100;
A = 16'h0032; B = 16'h0062; #100;
A = 16'h0032; B = 16'h0063; #100;
A = 16'h0032; B = 16'h0064; #100;
A = 16'h0032; B = 16'h0065; #100;
A = 16'h0032; B = 16'h0066; #100;
A = 16'h0032; B = 16'h0067; #100;
A = 16'h0032; B = 16'h0068; #100;
A = 16'h0032; B = 16'h0069; #100;
A = 16'h0032; B = 16'h006A; #100;
A = 16'h0032; B = 16'h006B; #100;
A = 16'h0032; B = 16'h006C; #100;
A = 16'h0032; B = 16'h006D; #100;
A = 16'h0032; B = 16'h006E; #100;
A = 16'h0032; B = 16'h006F; #100;
A = 16'h0032; B = 16'h0070; #100;
A = 16'h0032; B = 16'h0071; #100;
A = 16'h0032; B = 16'h0072; #100;
A = 16'h0032; B = 16'h0073; #100;
A = 16'h0032; B = 16'h0074; #100;
A = 16'h0032; B = 16'h0075; #100;
A = 16'h0032; B = 16'h0076; #100;
A = 16'h0032; B = 16'h0077; #100;
A = 16'h0032; B = 16'h0078; #100;
A = 16'h0032; B = 16'h0079; #100;
A = 16'h0032; B = 16'h007A; #100;
A = 16'h0032; B = 16'h007B; #100;
A = 16'h0032; B = 16'h007C; #100;
A = 16'h0032; B = 16'h007D; #100;
A = 16'h0032; B = 16'h007E; #100;
A = 16'h0032; B = 16'h007F; #100;
A = 16'h0032; B = 16'h0080; #100;
A = 16'h0032; B = 16'h0081; #100;
A = 16'h0032; B = 16'h0082; #100;
A = 16'h0032; B = 16'h0083; #100;
A = 16'h0032; B = 16'h0084; #100;
A = 16'h0032; B = 16'h0085; #100;
A = 16'h0032; B = 16'h0086; #100;
A = 16'h0032; B = 16'h0087; #100;
A = 16'h0032; B = 16'h0088; #100;
A = 16'h0032; B = 16'h0089; #100;
A = 16'h0032; B = 16'h008A; #100;
A = 16'h0032; B = 16'h008B; #100;
A = 16'h0032; B = 16'h008C; #100;
A = 16'h0032; B = 16'h008D; #100;
A = 16'h0032; B = 16'h008E; #100;
A = 16'h0032; B = 16'h008F; #100;
A = 16'h0032; B = 16'h0090; #100;
A = 16'h0032; B = 16'h0091; #100;
A = 16'h0032; B = 16'h0092; #100;
A = 16'h0032; B = 16'h0093; #100;
A = 16'h0032; B = 16'h0094; #100;
A = 16'h0032; B = 16'h0095; #100;
A = 16'h0032; B = 16'h0096; #100;
A = 16'h0032; B = 16'h0097; #100;
A = 16'h0032; B = 16'h0098; #100;
A = 16'h0032; B = 16'h0099; #100;
A = 16'h0032; B = 16'h009A; #100;
A = 16'h0032; B = 16'h009B; #100;
A = 16'h0032; B = 16'h009C; #100;
A = 16'h0032; B = 16'h009D; #100;
A = 16'h0032; B = 16'h009E; #100;
A = 16'h0032; B = 16'h009F; #100;
A = 16'h0032; B = 16'h00A0; #100;
A = 16'h0032; B = 16'h00A1; #100;
A = 16'h0032; B = 16'h00A2; #100;
A = 16'h0032; B = 16'h00A3; #100;
A = 16'h0032; B = 16'h00A4; #100;
A = 16'h0032; B = 16'h00A5; #100;
A = 16'h0032; B = 16'h00A6; #100;
A = 16'h0032; B = 16'h00A7; #100;
A = 16'h0032; B = 16'h00A8; #100;
A = 16'h0032; B = 16'h00A9; #100;
A = 16'h0032; B = 16'h00AA; #100;
A = 16'h0032; B = 16'h00AB; #100;
A = 16'h0032; B = 16'h00AC; #100;
A = 16'h0032; B = 16'h00AD; #100;
A = 16'h0032; B = 16'h00AE; #100;
A = 16'h0032; B = 16'h00AF; #100;
A = 16'h0032; B = 16'h00B0; #100;
A = 16'h0032; B = 16'h00B1; #100;
A = 16'h0032; B = 16'h00B2; #100;
A = 16'h0032; B = 16'h00B3; #100;
A = 16'h0032; B = 16'h00B4; #100;
A = 16'h0032; B = 16'h00B5; #100;
A = 16'h0032; B = 16'h00B6; #100;
A = 16'h0032; B = 16'h00B7; #100;
A = 16'h0032; B = 16'h00B8; #100;
A = 16'h0032; B = 16'h00B9; #100;
A = 16'h0032; B = 16'h00BA; #100;
A = 16'h0032; B = 16'h00BB; #100;
A = 16'h0032; B = 16'h00BC; #100;
A = 16'h0032; B = 16'h00BD; #100;
A = 16'h0032; B = 16'h00BE; #100;
A = 16'h0032; B = 16'h00BF; #100;
A = 16'h0032; B = 16'h00C0; #100;
A = 16'h0032; B = 16'h00C1; #100;
A = 16'h0032; B = 16'h00C2; #100;
A = 16'h0032; B = 16'h00C3; #100;
A = 16'h0032; B = 16'h00C4; #100;
A = 16'h0032; B = 16'h00C5; #100;
A = 16'h0032; B = 16'h00C6; #100;
A = 16'h0032; B = 16'h00C7; #100;
A = 16'h0032; B = 16'h00C8; #100;
A = 16'h0032; B = 16'h00C9; #100;
A = 16'h0032; B = 16'h00CA; #100;
A = 16'h0032; B = 16'h00CB; #100;
A = 16'h0032; B = 16'h00CC; #100;
A = 16'h0032; B = 16'h00CD; #100;
A = 16'h0032; B = 16'h00CE; #100;
A = 16'h0032; B = 16'h00CF; #100;
A = 16'h0032; B = 16'h00D0; #100;
A = 16'h0032; B = 16'h00D1; #100;
A = 16'h0032; B = 16'h00D2; #100;
A = 16'h0032; B = 16'h00D3; #100;
A = 16'h0032; B = 16'h00D4; #100;
A = 16'h0032; B = 16'h00D5; #100;
A = 16'h0032; B = 16'h00D6; #100;
A = 16'h0032; B = 16'h00D7; #100;
A = 16'h0032; B = 16'h00D8; #100;
A = 16'h0032; B = 16'h00D9; #100;
A = 16'h0032; B = 16'h00DA; #100;
A = 16'h0032; B = 16'h00DB; #100;
A = 16'h0032; B = 16'h00DC; #100;
A = 16'h0032; B = 16'h00DD; #100;
A = 16'h0032; B = 16'h00DE; #100;
A = 16'h0032; B = 16'h00DF; #100;
A = 16'h0032; B = 16'h00E0; #100;
A = 16'h0032; B = 16'h00E1; #100;
A = 16'h0032; B = 16'h00E2; #100;
A = 16'h0032; B = 16'h00E3; #100;
A = 16'h0032; B = 16'h00E4; #100;
A = 16'h0032; B = 16'h00E5; #100;
A = 16'h0032; B = 16'h00E6; #100;
A = 16'h0032; B = 16'h00E7; #100;
A = 16'h0032; B = 16'h00E8; #100;
A = 16'h0032; B = 16'h00E9; #100;
A = 16'h0032; B = 16'h00EA; #100;
A = 16'h0032; B = 16'h00EB; #100;
A = 16'h0032; B = 16'h00EC; #100;
A = 16'h0032; B = 16'h00ED; #100;
A = 16'h0032; B = 16'h00EE; #100;
A = 16'h0032; B = 16'h00EF; #100;
A = 16'h0032; B = 16'h00F0; #100;
A = 16'h0032; B = 16'h00F1; #100;
A = 16'h0032; B = 16'h00F2; #100;
A = 16'h0032; B = 16'h00F3; #100;
A = 16'h0032; B = 16'h00F4; #100;
A = 16'h0032; B = 16'h00F5; #100;
A = 16'h0032; B = 16'h00F6; #100;
A = 16'h0032; B = 16'h00F7; #100;
A = 16'h0032; B = 16'h00F8; #100;
A = 16'h0032; B = 16'h00F9; #100;
A = 16'h0032; B = 16'h00FA; #100;
A = 16'h0032; B = 16'h00FB; #100;
A = 16'h0032; B = 16'h00FC; #100;
A = 16'h0032; B = 16'h00FD; #100;
A = 16'h0032; B = 16'h00FE; #100;
A = 16'h0032; B = 16'h00FF; #100;
A = 16'h0033; B = 16'h000; #100;
A = 16'h0033; B = 16'h001; #100;
A = 16'h0033; B = 16'h002; #100;
A = 16'h0033; B = 16'h003; #100;
A = 16'h0033; B = 16'h004; #100;
A = 16'h0033; B = 16'h005; #100;
A = 16'h0033; B = 16'h006; #100;
A = 16'h0033; B = 16'h007; #100;
A = 16'h0033; B = 16'h008; #100;
A = 16'h0033; B = 16'h009; #100;
A = 16'h0033; B = 16'h00A; #100;
A = 16'h0033; B = 16'h00B; #100;
A = 16'h0033; B = 16'h00C; #100;
A = 16'h0033; B = 16'h00D; #100;
A = 16'h0033; B = 16'h00E; #100;
A = 16'h0033; B = 16'h00F; #100;
A = 16'h0033; B = 16'h0010; #100;
A = 16'h0033; B = 16'h0011; #100;
A = 16'h0033; B = 16'h0012; #100;
A = 16'h0033; B = 16'h0013; #100;
A = 16'h0033; B = 16'h0014; #100;
A = 16'h0033; B = 16'h0015; #100;
A = 16'h0033; B = 16'h0016; #100;
A = 16'h0033; B = 16'h0017; #100;
A = 16'h0033; B = 16'h0018; #100;
A = 16'h0033; B = 16'h0019; #100;
A = 16'h0033; B = 16'h001A; #100;
A = 16'h0033; B = 16'h001B; #100;
A = 16'h0033; B = 16'h001C; #100;
A = 16'h0033; B = 16'h001D; #100;
A = 16'h0033; B = 16'h001E; #100;
A = 16'h0033; B = 16'h001F; #100;
A = 16'h0033; B = 16'h0020; #100;
A = 16'h0033; B = 16'h0021; #100;
A = 16'h0033; B = 16'h0022; #100;
A = 16'h0033; B = 16'h0023; #100;
A = 16'h0033; B = 16'h0024; #100;
A = 16'h0033; B = 16'h0025; #100;
A = 16'h0033; B = 16'h0026; #100;
A = 16'h0033; B = 16'h0027; #100;
A = 16'h0033; B = 16'h0028; #100;
A = 16'h0033; B = 16'h0029; #100;
A = 16'h0033; B = 16'h002A; #100;
A = 16'h0033; B = 16'h002B; #100;
A = 16'h0033; B = 16'h002C; #100;
A = 16'h0033; B = 16'h002D; #100;
A = 16'h0033; B = 16'h002E; #100;
A = 16'h0033; B = 16'h002F; #100;
A = 16'h0033; B = 16'h0030; #100;
A = 16'h0033; B = 16'h0031; #100;
A = 16'h0033; B = 16'h0032; #100;
A = 16'h0033; B = 16'h0033; #100;
A = 16'h0033; B = 16'h0034; #100;
A = 16'h0033; B = 16'h0035; #100;
A = 16'h0033; B = 16'h0036; #100;
A = 16'h0033; B = 16'h0037; #100;
A = 16'h0033; B = 16'h0038; #100;
A = 16'h0033; B = 16'h0039; #100;
A = 16'h0033; B = 16'h003A; #100;
A = 16'h0033; B = 16'h003B; #100;
A = 16'h0033; B = 16'h003C; #100;
A = 16'h0033; B = 16'h003D; #100;
A = 16'h0033; B = 16'h003E; #100;
A = 16'h0033; B = 16'h003F; #100;
A = 16'h0033; B = 16'h0040; #100;
A = 16'h0033; B = 16'h0041; #100;
A = 16'h0033; B = 16'h0042; #100;
A = 16'h0033; B = 16'h0043; #100;
A = 16'h0033; B = 16'h0044; #100;
A = 16'h0033; B = 16'h0045; #100;
A = 16'h0033; B = 16'h0046; #100;
A = 16'h0033; B = 16'h0047; #100;
A = 16'h0033; B = 16'h0048; #100;
A = 16'h0033; B = 16'h0049; #100;
A = 16'h0033; B = 16'h004A; #100;
A = 16'h0033; B = 16'h004B; #100;
A = 16'h0033; B = 16'h004C; #100;
A = 16'h0033; B = 16'h004D; #100;
A = 16'h0033; B = 16'h004E; #100;
A = 16'h0033; B = 16'h004F; #100;
A = 16'h0033; B = 16'h0050; #100;
A = 16'h0033; B = 16'h0051; #100;
A = 16'h0033; B = 16'h0052; #100;
A = 16'h0033; B = 16'h0053; #100;
A = 16'h0033; B = 16'h0054; #100;
A = 16'h0033; B = 16'h0055; #100;
A = 16'h0033; B = 16'h0056; #100;
A = 16'h0033; B = 16'h0057; #100;
A = 16'h0033; B = 16'h0058; #100;
A = 16'h0033; B = 16'h0059; #100;
A = 16'h0033; B = 16'h005A; #100;
A = 16'h0033; B = 16'h005B; #100;
A = 16'h0033; B = 16'h005C; #100;
A = 16'h0033; B = 16'h005D; #100;
A = 16'h0033; B = 16'h005E; #100;
A = 16'h0033; B = 16'h005F; #100;
A = 16'h0033; B = 16'h0060; #100;
A = 16'h0033; B = 16'h0061; #100;
A = 16'h0033; B = 16'h0062; #100;
A = 16'h0033; B = 16'h0063; #100;
A = 16'h0033; B = 16'h0064; #100;
A = 16'h0033; B = 16'h0065; #100;
A = 16'h0033; B = 16'h0066; #100;
A = 16'h0033; B = 16'h0067; #100;
A = 16'h0033; B = 16'h0068; #100;
A = 16'h0033; B = 16'h0069; #100;
A = 16'h0033; B = 16'h006A; #100;
A = 16'h0033; B = 16'h006B; #100;
A = 16'h0033; B = 16'h006C; #100;
A = 16'h0033; B = 16'h006D; #100;
A = 16'h0033; B = 16'h006E; #100;
A = 16'h0033; B = 16'h006F; #100;
A = 16'h0033; B = 16'h0070; #100;
A = 16'h0033; B = 16'h0071; #100;
A = 16'h0033; B = 16'h0072; #100;
A = 16'h0033; B = 16'h0073; #100;
A = 16'h0033; B = 16'h0074; #100;
A = 16'h0033; B = 16'h0075; #100;
A = 16'h0033; B = 16'h0076; #100;
A = 16'h0033; B = 16'h0077; #100;
A = 16'h0033; B = 16'h0078; #100;
A = 16'h0033; B = 16'h0079; #100;
A = 16'h0033; B = 16'h007A; #100;
A = 16'h0033; B = 16'h007B; #100;
A = 16'h0033; B = 16'h007C; #100;
A = 16'h0033; B = 16'h007D; #100;
A = 16'h0033; B = 16'h007E; #100;
A = 16'h0033; B = 16'h007F; #100;
A = 16'h0033; B = 16'h0080; #100;
A = 16'h0033; B = 16'h0081; #100;
A = 16'h0033; B = 16'h0082; #100;
A = 16'h0033; B = 16'h0083; #100;
A = 16'h0033; B = 16'h0084; #100;
A = 16'h0033; B = 16'h0085; #100;
A = 16'h0033; B = 16'h0086; #100;
A = 16'h0033; B = 16'h0087; #100;
A = 16'h0033; B = 16'h0088; #100;
A = 16'h0033; B = 16'h0089; #100;
A = 16'h0033; B = 16'h008A; #100;
A = 16'h0033; B = 16'h008B; #100;
A = 16'h0033; B = 16'h008C; #100;
A = 16'h0033; B = 16'h008D; #100;
A = 16'h0033; B = 16'h008E; #100;
A = 16'h0033; B = 16'h008F; #100;
A = 16'h0033; B = 16'h0090; #100;
A = 16'h0033; B = 16'h0091; #100;
A = 16'h0033; B = 16'h0092; #100;
A = 16'h0033; B = 16'h0093; #100;
A = 16'h0033; B = 16'h0094; #100;
A = 16'h0033; B = 16'h0095; #100;
A = 16'h0033; B = 16'h0096; #100;
A = 16'h0033; B = 16'h0097; #100;
A = 16'h0033; B = 16'h0098; #100;
A = 16'h0033; B = 16'h0099; #100;
A = 16'h0033; B = 16'h009A; #100;
A = 16'h0033; B = 16'h009B; #100;
A = 16'h0033; B = 16'h009C; #100;
A = 16'h0033; B = 16'h009D; #100;
A = 16'h0033; B = 16'h009E; #100;
A = 16'h0033; B = 16'h009F; #100;
A = 16'h0033; B = 16'h00A0; #100;
A = 16'h0033; B = 16'h00A1; #100;
A = 16'h0033; B = 16'h00A2; #100;
A = 16'h0033; B = 16'h00A3; #100;
A = 16'h0033; B = 16'h00A4; #100;
A = 16'h0033; B = 16'h00A5; #100;
A = 16'h0033; B = 16'h00A6; #100;
A = 16'h0033; B = 16'h00A7; #100;
A = 16'h0033; B = 16'h00A8; #100;
A = 16'h0033; B = 16'h00A9; #100;
A = 16'h0033; B = 16'h00AA; #100;
A = 16'h0033; B = 16'h00AB; #100;
A = 16'h0033; B = 16'h00AC; #100;
A = 16'h0033; B = 16'h00AD; #100;
A = 16'h0033; B = 16'h00AE; #100;
A = 16'h0033; B = 16'h00AF; #100;
A = 16'h0033; B = 16'h00B0; #100;
A = 16'h0033; B = 16'h00B1; #100;
A = 16'h0033; B = 16'h00B2; #100;
A = 16'h0033; B = 16'h00B3; #100;
A = 16'h0033; B = 16'h00B4; #100;
A = 16'h0033; B = 16'h00B5; #100;
A = 16'h0033; B = 16'h00B6; #100;
A = 16'h0033; B = 16'h00B7; #100;
A = 16'h0033; B = 16'h00B8; #100;
A = 16'h0033; B = 16'h00B9; #100;
A = 16'h0033; B = 16'h00BA; #100;
A = 16'h0033; B = 16'h00BB; #100;
A = 16'h0033; B = 16'h00BC; #100;
A = 16'h0033; B = 16'h00BD; #100;
A = 16'h0033; B = 16'h00BE; #100;
A = 16'h0033; B = 16'h00BF; #100;
A = 16'h0033; B = 16'h00C0; #100;
A = 16'h0033; B = 16'h00C1; #100;
A = 16'h0033; B = 16'h00C2; #100;
A = 16'h0033; B = 16'h00C3; #100;
A = 16'h0033; B = 16'h00C4; #100;
A = 16'h0033; B = 16'h00C5; #100;
A = 16'h0033; B = 16'h00C6; #100;
A = 16'h0033; B = 16'h00C7; #100;
A = 16'h0033; B = 16'h00C8; #100;
A = 16'h0033; B = 16'h00C9; #100;
A = 16'h0033; B = 16'h00CA; #100;
A = 16'h0033; B = 16'h00CB; #100;
A = 16'h0033; B = 16'h00CC; #100;
A = 16'h0033; B = 16'h00CD; #100;
A = 16'h0033; B = 16'h00CE; #100;
A = 16'h0033; B = 16'h00CF; #100;
A = 16'h0033; B = 16'h00D0; #100;
A = 16'h0033; B = 16'h00D1; #100;
A = 16'h0033; B = 16'h00D2; #100;
A = 16'h0033; B = 16'h00D3; #100;
A = 16'h0033; B = 16'h00D4; #100;
A = 16'h0033; B = 16'h00D5; #100;
A = 16'h0033; B = 16'h00D6; #100;
A = 16'h0033; B = 16'h00D7; #100;
A = 16'h0033; B = 16'h00D8; #100;
A = 16'h0033; B = 16'h00D9; #100;
A = 16'h0033; B = 16'h00DA; #100;
A = 16'h0033; B = 16'h00DB; #100;
A = 16'h0033; B = 16'h00DC; #100;
A = 16'h0033; B = 16'h00DD; #100;
A = 16'h0033; B = 16'h00DE; #100;
A = 16'h0033; B = 16'h00DF; #100;
A = 16'h0033; B = 16'h00E0; #100;
A = 16'h0033; B = 16'h00E1; #100;
A = 16'h0033; B = 16'h00E2; #100;
A = 16'h0033; B = 16'h00E3; #100;
A = 16'h0033; B = 16'h00E4; #100;
A = 16'h0033; B = 16'h00E5; #100;
A = 16'h0033; B = 16'h00E6; #100;
A = 16'h0033; B = 16'h00E7; #100;
A = 16'h0033; B = 16'h00E8; #100;
A = 16'h0033; B = 16'h00E9; #100;
A = 16'h0033; B = 16'h00EA; #100;
A = 16'h0033; B = 16'h00EB; #100;
A = 16'h0033; B = 16'h00EC; #100;
A = 16'h0033; B = 16'h00ED; #100;
A = 16'h0033; B = 16'h00EE; #100;
A = 16'h0033; B = 16'h00EF; #100;
A = 16'h0033; B = 16'h00F0; #100;
A = 16'h0033; B = 16'h00F1; #100;
A = 16'h0033; B = 16'h00F2; #100;
A = 16'h0033; B = 16'h00F3; #100;
A = 16'h0033; B = 16'h00F4; #100;
A = 16'h0033; B = 16'h00F5; #100;
A = 16'h0033; B = 16'h00F6; #100;
A = 16'h0033; B = 16'h00F7; #100;
A = 16'h0033; B = 16'h00F8; #100;
A = 16'h0033; B = 16'h00F9; #100;
A = 16'h0033; B = 16'h00FA; #100;
A = 16'h0033; B = 16'h00FB; #100;
A = 16'h0033; B = 16'h00FC; #100;
A = 16'h0033; B = 16'h00FD; #100;
A = 16'h0033; B = 16'h00FE; #100;
A = 16'h0033; B = 16'h00FF; #100;
A = 16'h0034; B = 16'h000; #100;
A = 16'h0034; B = 16'h001; #100;
A = 16'h0034; B = 16'h002; #100;
A = 16'h0034; B = 16'h003; #100;
A = 16'h0034; B = 16'h004; #100;
A = 16'h0034; B = 16'h005; #100;
A = 16'h0034; B = 16'h006; #100;
A = 16'h0034; B = 16'h007; #100;
A = 16'h0034; B = 16'h008; #100;
A = 16'h0034; B = 16'h009; #100;
A = 16'h0034; B = 16'h00A; #100;
A = 16'h0034; B = 16'h00B; #100;
A = 16'h0034; B = 16'h00C; #100;
A = 16'h0034; B = 16'h00D; #100;
A = 16'h0034; B = 16'h00E; #100;
A = 16'h0034; B = 16'h00F; #100;
A = 16'h0034; B = 16'h0010; #100;
A = 16'h0034; B = 16'h0011; #100;
A = 16'h0034; B = 16'h0012; #100;
A = 16'h0034; B = 16'h0013; #100;
A = 16'h0034; B = 16'h0014; #100;
A = 16'h0034; B = 16'h0015; #100;
A = 16'h0034; B = 16'h0016; #100;
A = 16'h0034; B = 16'h0017; #100;
A = 16'h0034; B = 16'h0018; #100;
A = 16'h0034; B = 16'h0019; #100;
A = 16'h0034; B = 16'h001A; #100;
A = 16'h0034; B = 16'h001B; #100;
A = 16'h0034; B = 16'h001C; #100;
A = 16'h0034; B = 16'h001D; #100;
A = 16'h0034; B = 16'h001E; #100;
A = 16'h0034; B = 16'h001F; #100;
A = 16'h0034; B = 16'h0020; #100;
A = 16'h0034; B = 16'h0021; #100;
A = 16'h0034; B = 16'h0022; #100;
A = 16'h0034; B = 16'h0023; #100;
A = 16'h0034; B = 16'h0024; #100;
A = 16'h0034; B = 16'h0025; #100;
A = 16'h0034; B = 16'h0026; #100;
A = 16'h0034; B = 16'h0027; #100;
A = 16'h0034; B = 16'h0028; #100;
A = 16'h0034; B = 16'h0029; #100;
A = 16'h0034; B = 16'h002A; #100;
A = 16'h0034; B = 16'h002B; #100;
A = 16'h0034; B = 16'h002C; #100;
A = 16'h0034; B = 16'h002D; #100;
A = 16'h0034; B = 16'h002E; #100;
A = 16'h0034; B = 16'h002F; #100;
A = 16'h0034; B = 16'h0030; #100;
A = 16'h0034; B = 16'h0031; #100;
A = 16'h0034; B = 16'h0032; #100;
A = 16'h0034; B = 16'h0033; #100;
A = 16'h0034; B = 16'h0034; #100;
A = 16'h0034; B = 16'h0035; #100;
A = 16'h0034; B = 16'h0036; #100;
A = 16'h0034; B = 16'h0037; #100;
A = 16'h0034; B = 16'h0038; #100;
A = 16'h0034; B = 16'h0039; #100;
A = 16'h0034; B = 16'h003A; #100;
A = 16'h0034; B = 16'h003B; #100;
A = 16'h0034; B = 16'h003C; #100;
A = 16'h0034; B = 16'h003D; #100;
A = 16'h0034; B = 16'h003E; #100;
A = 16'h0034; B = 16'h003F; #100;
A = 16'h0034; B = 16'h0040; #100;
A = 16'h0034; B = 16'h0041; #100;
A = 16'h0034; B = 16'h0042; #100;
A = 16'h0034; B = 16'h0043; #100;
A = 16'h0034; B = 16'h0044; #100;
A = 16'h0034; B = 16'h0045; #100;
A = 16'h0034; B = 16'h0046; #100;
A = 16'h0034; B = 16'h0047; #100;
A = 16'h0034; B = 16'h0048; #100;
A = 16'h0034; B = 16'h0049; #100;
A = 16'h0034; B = 16'h004A; #100;
A = 16'h0034; B = 16'h004B; #100;
A = 16'h0034; B = 16'h004C; #100;
A = 16'h0034; B = 16'h004D; #100;
A = 16'h0034; B = 16'h004E; #100;
A = 16'h0034; B = 16'h004F; #100;
A = 16'h0034; B = 16'h0050; #100;
A = 16'h0034; B = 16'h0051; #100;
A = 16'h0034; B = 16'h0052; #100;
A = 16'h0034; B = 16'h0053; #100;
A = 16'h0034; B = 16'h0054; #100;
A = 16'h0034; B = 16'h0055; #100;
A = 16'h0034; B = 16'h0056; #100;
A = 16'h0034; B = 16'h0057; #100;
A = 16'h0034; B = 16'h0058; #100;
A = 16'h0034; B = 16'h0059; #100;
A = 16'h0034; B = 16'h005A; #100;
A = 16'h0034; B = 16'h005B; #100;
A = 16'h0034; B = 16'h005C; #100;
A = 16'h0034; B = 16'h005D; #100;
A = 16'h0034; B = 16'h005E; #100;
A = 16'h0034; B = 16'h005F; #100;
A = 16'h0034; B = 16'h0060; #100;
A = 16'h0034; B = 16'h0061; #100;
A = 16'h0034; B = 16'h0062; #100;
A = 16'h0034; B = 16'h0063; #100;
A = 16'h0034; B = 16'h0064; #100;
A = 16'h0034; B = 16'h0065; #100;
A = 16'h0034; B = 16'h0066; #100;
A = 16'h0034; B = 16'h0067; #100;
A = 16'h0034; B = 16'h0068; #100;
A = 16'h0034; B = 16'h0069; #100;
A = 16'h0034; B = 16'h006A; #100;
A = 16'h0034; B = 16'h006B; #100;
A = 16'h0034; B = 16'h006C; #100;
A = 16'h0034; B = 16'h006D; #100;
A = 16'h0034; B = 16'h006E; #100;
A = 16'h0034; B = 16'h006F; #100;
A = 16'h0034; B = 16'h0070; #100;
A = 16'h0034; B = 16'h0071; #100;
A = 16'h0034; B = 16'h0072; #100;
A = 16'h0034; B = 16'h0073; #100;
A = 16'h0034; B = 16'h0074; #100;
A = 16'h0034; B = 16'h0075; #100;
A = 16'h0034; B = 16'h0076; #100;
A = 16'h0034; B = 16'h0077; #100;
A = 16'h0034; B = 16'h0078; #100;
A = 16'h0034; B = 16'h0079; #100;
A = 16'h0034; B = 16'h007A; #100;
A = 16'h0034; B = 16'h007B; #100;
A = 16'h0034; B = 16'h007C; #100;
A = 16'h0034; B = 16'h007D; #100;
A = 16'h0034; B = 16'h007E; #100;
A = 16'h0034; B = 16'h007F; #100;
A = 16'h0034; B = 16'h0080; #100;
A = 16'h0034; B = 16'h0081; #100;
A = 16'h0034; B = 16'h0082; #100;
A = 16'h0034; B = 16'h0083; #100;
A = 16'h0034; B = 16'h0084; #100;
A = 16'h0034; B = 16'h0085; #100;
A = 16'h0034; B = 16'h0086; #100;
A = 16'h0034; B = 16'h0087; #100;
A = 16'h0034; B = 16'h0088; #100;
A = 16'h0034; B = 16'h0089; #100;
A = 16'h0034; B = 16'h008A; #100;
A = 16'h0034; B = 16'h008B; #100;
A = 16'h0034; B = 16'h008C; #100;
A = 16'h0034; B = 16'h008D; #100;
A = 16'h0034; B = 16'h008E; #100;
A = 16'h0034; B = 16'h008F; #100;
A = 16'h0034; B = 16'h0090; #100;
A = 16'h0034; B = 16'h0091; #100;
A = 16'h0034; B = 16'h0092; #100;
A = 16'h0034; B = 16'h0093; #100;
A = 16'h0034; B = 16'h0094; #100;
A = 16'h0034; B = 16'h0095; #100;
A = 16'h0034; B = 16'h0096; #100;
A = 16'h0034; B = 16'h0097; #100;
A = 16'h0034; B = 16'h0098; #100;
A = 16'h0034; B = 16'h0099; #100;
A = 16'h0034; B = 16'h009A; #100;
A = 16'h0034; B = 16'h009B; #100;
A = 16'h0034; B = 16'h009C; #100;
A = 16'h0034; B = 16'h009D; #100;
A = 16'h0034; B = 16'h009E; #100;
A = 16'h0034; B = 16'h009F; #100;
A = 16'h0034; B = 16'h00A0; #100;
A = 16'h0034; B = 16'h00A1; #100;
A = 16'h0034; B = 16'h00A2; #100;
A = 16'h0034; B = 16'h00A3; #100;
A = 16'h0034; B = 16'h00A4; #100;
A = 16'h0034; B = 16'h00A5; #100;
A = 16'h0034; B = 16'h00A6; #100;
A = 16'h0034; B = 16'h00A7; #100;
A = 16'h0034; B = 16'h00A8; #100;
A = 16'h0034; B = 16'h00A9; #100;
A = 16'h0034; B = 16'h00AA; #100;
A = 16'h0034; B = 16'h00AB; #100;
A = 16'h0034; B = 16'h00AC; #100;
A = 16'h0034; B = 16'h00AD; #100;
A = 16'h0034; B = 16'h00AE; #100;
A = 16'h0034; B = 16'h00AF; #100;
A = 16'h0034; B = 16'h00B0; #100;
A = 16'h0034; B = 16'h00B1; #100;
A = 16'h0034; B = 16'h00B2; #100;
A = 16'h0034; B = 16'h00B3; #100;
A = 16'h0034; B = 16'h00B4; #100;
A = 16'h0034; B = 16'h00B5; #100;
A = 16'h0034; B = 16'h00B6; #100;
A = 16'h0034; B = 16'h00B7; #100;
A = 16'h0034; B = 16'h00B8; #100;
A = 16'h0034; B = 16'h00B9; #100;
A = 16'h0034; B = 16'h00BA; #100;
A = 16'h0034; B = 16'h00BB; #100;
A = 16'h0034; B = 16'h00BC; #100;
A = 16'h0034; B = 16'h00BD; #100;
A = 16'h0034; B = 16'h00BE; #100;
A = 16'h0034; B = 16'h00BF; #100;
A = 16'h0034; B = 16'h00C0; #100;
A = 16'h0034; B = 16'h00C1; #100;
A = 16'h0034; B = 16'h00C2; #100;
A = 16'h0034; B = 16'h00C3; #100;
A = 16'h0034; B = 16'h00C4; #100;
A = 16'h0034; B = 16'h00C5; #100;
A = 16'h0034; B = 16'h00C6; #100;
A = 16'h0034; B = 16'h00C7; #100;
A = 16'h0034; B = 16'h00C8; #100;
A = 16'h0034; B = 16'h00C9; #100;
A = 16'h0034; B = 16'h00CA; #100;
A = 16'h0034; B = 16'h00CB; #100;
A = 16'h0034; B = 16'h00CC; #100;
A = 16'h0034; B = 16'h00CD; #100;
A = 16'h0034; B = 16'h00CE; #100;
A = 16'h0034; B = 16'h00CF; #100;
A = 16'h0034; B = 16'h00D0; #100;
A = 16'h0034; B = 16'h00D1; #100;
A = 16'h0034; B = 16'h00D2; #100;
A = 16'h0034; B = 16'h00D3; #100;
A = 16'h0034; B = 16'h00D4; #100;
A = 16'h0034; B = 16'h00D5; #100;
A = 16'h0034; B = 16'h00D6; #100;
A = 16'h0034; B = 16'h00D7; #100;
A = 16'h0034; B = 16'h00D8; #100;
A = 16'h0034; B = 16'h00D9; #100;
A = 16'h0034; B = 16'h00DA; #100;
A = 16'h0034; B = 16'h00DB; #100;
A = 16'h0034; B = 16'h00DC; #100;
A = 16'h0034; B = 16'h00DD; #100;
A = 16'h0034; B = 16'h00DE; #100;
A = 16'h0034; B = 16'h00DF; #100;
A = 16'h0034; B = 16'h00E0; #100;
A = 16'h0034; B = 16'h00E1; #100;
A = 16'h0034; B = 16'h00E2; #100;
A = 16'h0034; B = 16'h00E3; #100;
A = 16'h0034; B = 16'h00E4; #100;
A = 16'h0034; B = 16'h00E5; #100;
A = 16'h0034; B = 16'h00E6; #100;
A = 16'h0034; B = 16'h00E7; #100;
A = 16'h0034; B = 16'h00E8; #100;
A = 16'h0034; B = 16'h00E9; #100;
A = 16'h0034; B = 16'h00EA; #100;
A = 16'h0034; B = 16'h00EB; #100;
A = 16'h0034; B = 16'h00EC; #100;
A = 16'h0034; B = 16'h00ED; #100;
A = 16'h0034; B = 16'h00EE; #100;
A = 16'h0034; B = 16'h00EF; #100;
A = 16'h0034; B = 16'h00F0; #100;
A = 16'h0034; B = 16'h00F1; #100;
A = 16'h0034; B = 16'h00F2; #100;
A = 16'h0034; B = 16'h00F3; #100;
A = 16'h0034; B = 16'h00F4; #100;
A = 16'h0034; B = 16'h00F5; #100;
A = 16'h0034; B = 16'h00F6; #100;
A = 16'h0034; B = 16'h00F7; #100;
A = 16'h0034; B = 16'h00F8; #100;
A = 16'h0034; B = 16'h00F9; #100;
A = 16'h0034; B = 16'h00FA; #100;
A = 16'h0034; B = 16'h00FB; #100;
A = 16'h0034; B = 16'h00FC; #100;
A = 16'h0034; B = 16'h00FD; #100;
A = 16'h0034; B = 16'h00FE; #100;
A = 16'h0034; B = 16'h00FF; #100;
A = 16'h0035; B = 16'h000; #100;
A = 16'h0035; B = 16'h001; #100;
A = 16'h0035; B = 16'h002; #100;
A = 16'h0035; B = 16'h003; #100;
A = 16'h0035; B = 16'h004; #100;
A = 16'h0035; B = 16'h005; #100;
A = 16'h0035; B = 16'h006; #100;
A = 16'h0035; B = 16'h007; #100;
A = 16'h0035; B = 16'h008; #100;
A = 16'h0035; B = 16'h009; #100;
A = 16'h0035; B = 16'h00A; #100;
A = 16'h0035; B = 16'h00B; #100;
A = 16'h0035; B = 16'h00C; #100;
A = 16'h0035; B = 16'h00D; #100;
A = 16'h0035; B = 16'h00E; #100;
A = 16'h0035; B = 16'h00F; #100;
A = 16'h0035; B = 16'h0010; #100;
A = 16'h0035; B = 16'h0011; #100;
A = 16'h0035; B = 16'h0012; #100;
A = 16'h0035; B = 16'h0013; #100;
A = 16'h0035; B = 16'h0014; #100;
A = 16'h0035; B = 16'h0015; #100;
A = 16'h0035; B = 16'h0016; #100;
A = 16'h0035; B = 16'h0017; #100;
A = 16'h0035; B = 16'h0018; #100;
A = 16'h0035; B = 16'h0019; #100;
A = 16'h0035; B = 16'h001A; #100;
A = 16'h0035; B = 16'h001B; #100;
A = 16'h0035; B = 16'h001C; #100;
A = 16'h0035; B = 16'h001D; #100;
A = 16'h0035; B = 16'h001E; #100;
A = 16'h0035; B = 16'h001F; #100;
A = 16'h0035; B = 16'h0020; #100;
A = 16'h0035; B = 16'h0021; #100;
A = 16'h0035; B = 16'h0022; #100;
A = 16'h0035; B = 16'h0023; #100;
A = 16'h0035; B = 16'h0024; #100;
A = 16'h0035; B = 16'h0025; #100;
A = 16'h0035; B = 16'h0026; #100;
A = 16'h0035; B = 16'h0027; #100;
A = 16'h0035; B = 16'h0028; #100;
A = 16'h0035; B = 16'h0029; #100;
A = 16'h0035; B = 16'h002A; #100;
A = 16'h0035; B = 16'h002B; #100;
A = 16'h0035; B = 16'h002C; #100;
A = 16'h0035; B = 16'h002D; #100;
A = 16'h0035; B = 16'h002E; #100;
A = 16'h0035; B = 16'h002F; #100;
A = 16'h0035; B = 16'h0030; #100;
A = 16'h0035; B = 16'h0031; #100;
A = 16'h0035; B = 16'h0032; #100;
A = 16'h0035; B = 16'h0033; #100;
A = 16'h0035; B = 16'h0034; #100;
A = 16'h0035; B = 16'h0035; #100;
A = 16'h0035; B = 16'h0036; #100;
A = 16'h0035; B = 16'h0037; #100;
A = 16'h0035; B = 16'h0038; #100;
A = 16'h0035; B = 16'h0039; #100;
A = 16'h0035; B = 16'h003A; #100;
A = 16'h0035; B = 16'h003B; #100;
A = 16'h0035; B = 16'h003C; #100;
A = 16'h0035; B = 16'h003D; #100;
A = 16'h0035; B = 16'h003E; #100;
A = 16'h0035; B = 16'h003F; #100;
A = 16'h0035; B = 16'h0040; #100;
A = 16'h0035; B = 16'h0041; #100;
A = 16'h0035; B = 16'h0042; #100;
A = 16'h0035; B = 16'h0043; #100;
A = 16'h0035; B = 16'h0044; #100;
A = 16'h0035; B = 16'h0045; #100;
A = 16'h0035; B = 16'h0046; #100;
A = 16'h0035; B = 16'h0047; #100;
A = 16'h0035; B = 16'h0048; #100;
A = 16'h0035; B = 16'h0049; #100;
A = 16'h0035; B = 16'h004A; #100;
A = 16'h0035; B = 16'h004B; #100;
A = 16'h0035; B = 16'h004C; #100;
A = 16'h0035; B = 16'h004D; #100;
A = 16'h0035; B = 16'h004E; #100;
A = 16'h0035; B = 16'h004F; #100;
A = 16'h0035; B = 16'h0050; #100;
A = 16'h0035; B = 16'h0051; #100;
A = 16'h0035; B = 16'h0052; #100;
A = 16'h0035; B = 16'h0053; #100;
A = 16'h0035; B = 16'h0054; #100;
A = 16'h0035; B = 16'h0055; #100;
A = 16'h0035; B = 16'h0056; #100;
A = 16'h0035; B = 16'h0057; #100;
A = 16'h0035; B = 16'h0058; #100;
A = 16'h0035; B = 16'h0059; #100;
A = 16'h0035; B = 16'h005A; #100;
A = 16'h0035; B = 16'h005B; #100;
A = 16'h0035; B = 16'h005C; #100;
A = 16'h0035; B = 16'h005D; #100;
A = 16'h0035; B = 16'h005E; #100;
A = 16'h0035; B = 16'h005F; #100;
A = 16'h0035; B = 16'h0060; #100;
A = 16'h0035; B = 16'h0061; #100;
A = 16'h0035; B = 16'h0062; #100;
A = 16'h0035; B = 16'h0063; #100;
A = 16'h0035; B = 16'h0064; #100;
A = 16'h0035; B = 16'h0065; #100;
A = 16'h0035; B = 16'h0066; #100;
A = 16'h0035; B = 16'h0067; #100;
A = 16'h0035; B = 16'h0068; #100;
A = 16'h0035; B = 16'h0069; #100;
A = 16'h0035; B = 16'h006A; #100;
A = 16'h0035; B = 16'h006B; #100;
A = 16'h0035; B = 16'h006C; #100;
A = 16'h0035; B = 16'h006D; #100;
A = 16'h0035; B = 16'h006E; #100;
A = 16'h0035; B = 16'h006F; #100;
A = 16'h0035; B = 16'h0070; #100;
A = 16'h0035; B = 16'h0071; #100;
A = 16'h0035; B = 16'h0072; #100;
A = 16'h0035; B = 16'h0073; #100;
A = 16'h0035; B = 16'h0074; #100;
A = 16'h0035; B = 16'h0075; #100;
A = 16'h0035; B = 16'h0076; #100;
A = 16'h0035; B = 16'h0077; #100;
A = 16'h0035; B = 16'h0078; #100;
A = 16'h0035; B = 16'h0079; #100;
A = 16'h0035; B = 16'h007A; #100;
A = 16'h0035; B = 16'h007B; #100;
A = 16'h0035; B = 16'h007C; #100;
A = 16'h0035; B = 16'h007D; #100;
A = 16'h0035; B = 16'h007E; #100;
A = 16'h0035; B = 16'h007F; #100;
A = 16'h0035; B = 16'h0080; #100;
A = 16'h0035; B = 16'h0081; #100;
A = 16'h0035; B = 16'h0082; #100;
A = 16'h0035; B = 16'h0083; #100;
A = 16'h0035; B = 16'h0084; #100;
A = 16'h0035; B = 16'h0085; #100;
A = 16'h0035; B = 16'h0086; #100;
A = 16'h0035; B = 16'h0087; #100;
A = 16'h0035; B = 16'h0088; #100;
A = 16'h0035; B = 16'h0089; #100;
A = 16'h0035; B = 16'h008A; #100;
A = 16'h0035; B = 16'h008B; #100;
A = 16'h0035; B = 16'h008C; #100;
A = 16'h0035; B = 16'h008D; #100;
A = 16'h0035; B = 16'h008E; #100;
A = 16'h0035; B = 16'h008F; #100;
A = 16'h0035; B = 16'h0090; #100;
A = 16'h0035; B = 16'h0091; #100;
A = 16'h0035; B = 16'h0092; #100;
A = 16'h0035; B = 16'h0093; #100;
A = 16'h0035; B = 16'h0094; #100;
A = 16'h0035; B = 16'h0095; #100;
A = 16'h0035; B = 16'h0096; #100;
A = 16'h0035; B = 16'h0097; #100;
A = 16'h0035; B = 16'h0098; #100;
A = 16'h0035; B = 16'h0099; #100;
A = 16'h0035; B = 16'h009A; #100;
A = 16'h0035; B = 16'h009B; #100;
A = 16'h0035; B = 16'h009C; #100;
A = 16'h0035; B = 16'h009D; #100;
A = 16'h0035; B = 16'h009E; #100;
A = 16'h0035; B = 16'h009F; #100;
A = 16'h0035; B = 16'h00A0; #100;
A = 16'h0035; B = 16'h00A1; #100;
A = 16'h0035; B = 16'h00A2; #100;
A = 16'h0035; B = 16'h00A3; #100;
A = 16'h0035; B = 16'h00A4; #100;
A = 16'h0035; B = 16'h00A5; #100;
A = 16'h0035; B = 16'h00A6; #100;
A = 16'h0035; B = 16'h00A7; #100;
A = 16'h0035; B = 16'h00A8; #100;
A = 16'h0035; B = 16'h00A9; #100;
A = 16'h0035; B = 16'h00AA; #100;
A = 16'h0035; B = 16'h00AB; #100;
A = 16'h0035; B = 16'h00AC; #100;
A = 16'h0035; B = 16'h00AD; #100;
A = 16'h0035; B = 16'h00AE; #100;
A = 16'h0035; B = 16'h00AF; #100;
A = 16'h0035; B = 16'h00B0; #100;
A = 16'h0035; B = 16'h00B1; #100;
A = 16'h0035; B = 16'h00B2; #100;
A = 16'h0035; B = 16'h00B3; #100;
A = 16'h0035; B = 16'h00B4; #100;
A = 16'h0035; B = 16'h00B5; #100;
A = 16'h0035; B = 16'h00B6; #100;
A = 16'h0035; B = 16'h00B7; #100;
A = 16'h0035; B = 16'h00B8; #100;
A = 16'h0035; B = 16'h00B9; #100;
A = 16'h0035; B = 16'h00BA; #100;
A = 16'h0035; B = 16'h00BB; #100;
A = 16'h0035; B = 16'h00BC; #100;
A = 16'h0035; B = 16'h00BD; #100;
A = 16'h0035; B = 16'h00BE; #100;
A = 16'h0035; B = 16'h00BF; #100;
A = 16'h0035; B = 16'h00C0; #100;
A = 16'h0035; B = 16'h00C1; #100;
A = 16'h0035; B = 16'h00C2; #100;
A = 16'h0035; B = 16'h00C3; #100;
A = 16'h0035; B = 16'h00C4; #100;
A = 16'h0035; B = 16'h00C5; #100;
A = 16'h0035; B = 16'h00C6; #100;
A = 16'h0035; B = 16'h00C7; #100;
A = 16'h0035; B = 16'h00C8; #100;
A = 16'h0035; B = 16'h00C9; #100;
A = 16'h0035; B = 16'h00CA; #100;
A = 16'h0035; B = 16'h00CB; #100;
A = 16'h0035; B = 16'h00CC; #100;
A = 16'h0035; B = 16'h00CD; #100;
A = 16'h0035; B = 16'h00CE; #100;
A = 16'h0035; B = 16'h00CF; #100;
A = 16'h0035; B = 16'h00D0; #100;
A = 16'h0035; B = 16'h00D1; #100;
A = 16'h0035; B = 16'h00D2; #100;
A = 16'h0035; B = 16'h00D3; #100;
A = 16'h0035; B = 16'h00D4; #100;
A = 16'h0035; B = 16'h00D5; #100;
A = 16'h0035; B = 16'h00D6; #100;
A = 16'h0035; B = 16'h00D7; #100;
A = 16'h0035; B = 16'h00D8; #100;
A = 16'h0035; B = 16'h00D9; #100;
A = 16'h0035; B = 16'h00DA; #100;
A = 16'h0035; B = 16'h00DB; #100;
A = 16'h0035; B = 16'h00DC; #100;
A = 16'h0035; B = 16'h00DD; #100;
A = 16'h0035; B = 16'h00DE; #100;
A = 16'h0035; B = 16'h00DF; #100;
A = 16'h0035; B = 16'h00E0; #100;
A = 16'h0035; B = 16'h00E1; #100;
A = 16'h0035; B = 16'h00E2; #100;
A = 16'h0035; B = 16'h00E3; #100;
A = 16'h0035; B = 16'h00E4; #100;
A = 16'h0035; B = 16'h00E5; #100;
A = 16'h0035; B = 16'h00E6; #100;
A = 16'h0035; B = 16'h00E7; #100;
A = 16'h0035; B = 16'h00E8; #100;
A = 16'h0035; B = 16'h00E9; #100;
A = 16'h0035; B = 16'h00EA; #100;
A = 16'h0035; B = 16'h00EB; #100;
A = 16'h0035; B = 16'h00EC; #100;
A = 16'h0035; B = 16'h00ED; #100;
A = 16'h0035; B = 16'h00EE; #100;
A = 16'h0035; B = 16'h00EF; #100;
A = 16'h0035; B = 16'h00F0; #100;
A = 16'h0035; B = 16'h00F1; #100;
A = 16'h0035; B = 16'h00F2; #100;
A = 16'h0035; B = 16'h00F3; #100;
A = 16'h0035; B = 16'h00F4; #100;
A = 16'h0035; B = 16'h00F5; #100;
A = 16'h0035; B = 16'h00F6; #100;
A = 16'h0035; B = 16'h00F7; #100;
A = 16'h0035; B = 16'h00F8; #100;
A = 16'h0035; B = 16'h00F9; #100;
A = 16'h0035; B = 16'h00FA; #100;
A = 16'h0035; B = 16'h00FB; #100;
A = 16'h0035; B = 16'h00FC; #100;
A = 16'h0035; B = 16'h00FD; #100;
A = 16'h0035; B = 16'h00FE; #100;
A = 16'h0035; B = 16'h00FF; #100;
A = 16'h0036; B = 16'h000; #100;
A = 16'h0036; B = 16'h001; #100;
A = 16'h0036; B = 16'h002; #100;
A = 16'h0036; B = 16'h003; #100;
A = 16'h0036; B = 16'h004; #100;
A = 16'h0036; B = 16'h005; #100;
A = 16'h0036; B = 16'h006; #100;
A = 16'h0036; B = 16'h007; #100;
A = 16'h0036; B = 16'h008; #100;
A = 16'h0036; B = 16'h009; #100;
A = 16'h0036; B = 16'h00A; #100;
A = 16'h0036; B = 16'h00B; #100;
A = 16'h0036; B = 16'h00C; #100;
A = 16'h0036; B = 16'h00D; #100;
A = 16'h0036; B = 16'h00E; #100;
A = 16'h0036; B = 16'h00F; #100;
A = 16'h0036; B = 16'h0010; #100;
A = 16'h0036; B = 16'h0011; #100;
A = 16'h0036; B = 16'h0012; #100;
A = 16'h0036; B = 16'h0013; #100;
A = 16'h0036; B = 16'h0014; #100;
A = 16'h0036; B = 16'h0015; #100;
A = 16'h0036; B = 16'h0016; #100;
A = 16'h0036; B = 16'h0017; #100;
A = 16'h0036; B = 16'h0018; #100;
A = 16'h0036; B = 16'h0019; #100;
A = 16'h0036; B = 16'h001A; #100;
A = 16'h0036; B = 16'h001B; #100;
A = 16'h0036; B = 16'h001C; #100;
A = 16'h0036; B = 16'h001D; #100;
A = 16'h0036; B = 16'h001E; #100;
A = 16'h0036; B = 16'h001F; #100;
A = 16'h0036; B = 16'h0020; #100;
A = 16'h0036; B = 16'h0021; #100;
A = 16'h0036; B = 16'h0022; #100;
A = 16'h0036; B = 16'h0023; #100;
A = 16'h0036; B = 16'h0024; #100;
A = 16'h0036; B = 16'h0025; #100;
A = 16'h0036; B = 16'h0026; #100;
A = 16'h0036; B = 16'h0027; #100;
A = 16'h0036; B = 16'h0028; #100;
A = 16'h0036; B = 16'h0029; #100;
A = 16'h0036; B = 16'h002A; #100;
A = 16'h0036; B = 16'h002B; #100;
A = 16'h0036; B = 16'h002C; #100;
A = 16'h0036; B = 16'h002D; #100;
A = 16'h0036; B = 16'h002E; #100;
A = 16'h0036; B = 16'h002F; #100;
A = 16'h0036; B = 16'h0030; #100;
A = 16'h0036; B = 16'h0031; #100;
A = 16'h0036; B = 16'h0032; #100;
A = 16'h0036; B = 16'h0033; #100;
A = 16'h0036; B = 16'h0034; #100;
A = 16'h0036; B = 16'h0035; #100;
A = 16'h0036; B = 16'h0036; #100;
A = 16'h0036; B = 16'h0037; #100;
A = 16'h0036; B = 16'h0038; #100;
A = 16'h0036; B = 16'h0039; #100;
A = 16'h0036; B = 16'h003A; #100;
A = 16'h0036; B = 16'h003B; #100;
A = 16'h0036; B = 16'h003C; #100;
A = 16'h0036; B = 16'h003D; #100;
A = 16'h0036; B = 16'h003E; #100;
A = 16'h0036; B = 16'h003F; #100;
A = 16'h0036; B = 16'h0040; #100;
A = 16'h0036; B = 16'h0041; #100;
A = 16'h0036; B = 16'h0042; #100;
A = 16'h0036; B = 16'h0043; #100;
A = 16'h0036; B = 16'h0044; #100;
A = 16'h0036; B = 16'h0045; #100;
A = 16'h0036; B = 16'h0046; #100;
A = 16'h0036; B = 16'h0047; #100;
A = 16'h0036; B = 16'h0048; #100;
A = 16'h0036; B = 16'h0049; #100;
A = 16'h0036; B = 16'h004A; #100;
A = 16'h0036; B = 16'h004B; #100;
A = 16'h0036; B = 16'h004C; #100;
A = 16'h0036; B = 16'h004D; #100;
A = 16'h0036; B = 16'h004E; #100;
A = 16'h0036; B = 16'h004F; #100;
A = 16'h0036; B = 16'h0050; #100;
A = 16'h0036; B = 16'h0051; #100;
A = 16'h0036; B = 16'h0052; #100;
A = 16'h0036; B = 16'h0053; #100;
A = 16'h0036; B = 16'h0054; #100;
A = 16'h0036; B = 16'h0055; #100;
A = 16'h0036; B = 16'h0056; #100;
A = 16'h0036; B = 16'h0057; #100;
A = 16'h0036; B = 16'h0058; #100;
A = 16'h0036; B = 16'h0059; #100;
A = 16'h0036; B = 16'h005A; #100;
A = 16'h0036; B = 16'h005B; #100;
A = 16'h0036; B = 16'h005C; #100;
A = 16'h0036; B = 16'h005D; #100;
A = 16'h0036; B = 16'h005E; #100;
A = 16'h0036; B = 16'h005F; #100;
A = 16'h0036; B = 16'h0060; #100;
A = 16'h0036; B = 16'h0061; #100;
A = 16'h0036; B = 16'h0062; #100;
A = 16'h0036; B = 16'h0063; #100;
A = 16'h0036; B = 16'h0064; #100;
A = 16'h0036; B = 16'h0065; #100;
A = 16'h0036; B = 16'h0066; #100;
A = 16'h0036; B = 16'h0067; #100;
A = 16'h0036; B = 16'h0068; #100;
A = 16'h0036; B = 16'h0069; #100;
A = 16'h0036; B = 16'h006A; #100;
A = 16'h0036; B = 16'h006B; #100;
A = 16'h0036; B = 16'h006C; #100;
A = 16'h0036; B = 16'h006D; #100;
A = 16'h0036; B = 16'h006E; #100;
A = 16'h0036; B = 16'h006F; #100;
A = 16'h0036; B = 16'h0070; #100;
A = 16'h0036; B = 16'h0071; #100;
A = 16'h0036; B = 16'h0072; #100;
A = 16'h0036; B = 16'h0073; #100;
A = 16'h0036; B = 16'h0074; #100;
A = 16'h0036; B = 16'h0075; #100;
A = 16'h0036; B = 16'h0076; #100;
A = 16'h0036; B = 16'h0077; #100;
A = 16'h0036; B = 16'h0078; #100;
A = 16'h0036; B = 16'h0079; #100;
A = 16'h0036; B = 16'h007A; #100;
A = 16'h0036; B = 16'h007B; #100;
A = 16'h0036; B = 16'h007C; #100;
A = 16'h0036; B = 16'h007D; #100;
A = 16'h0036; B = 16'h007E; #100;
A = 16'h0036; B = 16'h007F; #100;
A = 16'h0036; B = 16'h0080; #100;
A = 16'h0036; B = 16'h0081; #100;
A = 16'h0036; B = 16'h0082; #100;
A = 16'h0036; B = 16'h0083; #100;
A = 16'h0036; B = 16'h0084; #100;
A = 16'h0036; B = 16'h0085; #100;
A = 16'h0036; B = 16'h0086; #100;
A = 16'h0036; B = 16'h0087; #100;
A = 16'h0036; B = 16'h0088; #100;
A = 16'h0036; B = 16'h0089; #100;
A = 16'h0036; B = 16'h008A; #100;
A = 16'h0036; B = 16'h008B; #100;
A = 16'h0036; B = 16'h008C; #100;
A = 16'h0036; B = 16'h008D; #100;
A = 16'h0036; B = 16'h008E; #100;
A = 16'h0036; B = 16'h008F; #100;
A = 16'h0036; B = 16'h0090; #100;
A = 16'h0036; B = 16'h0091; #100;
A = 16'h0036; B = 16'h0092; #100;
A = 16'h0036; B = 16'h0093; #100;
A = 16'h0036; B = 16'h0094; #100;
A = 16'h0036; B = 16'h0095; #100;
A = 16'h0036; B = 16'h0096; #100;
A = 16'h0036; B = 16'h0097; #100;
A = 16'h0036; B = 16'h0098; #100;
A = 16'h0036; B = 16'h0099; #100;
A = 16'h0036; B = 16'h009A; #100;
A = 16'h0036; B = 16'h009B; #100;
A = 16'h0036; B = 16'h009C; #100;
A = 16'h0036; B = 16'h009D; #100;
A = 16'h0036; B = 16'h009E; #100;
A = 16'h0036; B = 16'h009F; #100;
A = 16'h0036; B = 16'h00A0; #100;
A = 16'h0036; B = 16'h00A1; #100;
A = 16'h0036; B = 16'h00A2; #100;
A = 16'h0036; B = 16'h00A3; #100;
A = 16'h0036; B = 16'h00A4; #100;
A = 16'h0036; B = 16'h00A5; #100;
A = 16'h0036; B = 16'h00A6; #100;
A = 16'h0036; B = 16'h00A7; #100;
A = 16'h0036; B = 16'h00A8; #100;
A = 16'h0036; B = 16'h00A9; #100;
A = 16'h0036; B = 16'h00AA; #100;
A = 16'h0036; B = 16'h00AB; #100;
A = 16'h0036; B = 16'h00AC; #100;
A = 16'h0036; B = 16'h00AD; #100;
A = 16'h0036; B = 16'h00AE; #100;
A = 16'h0036; B = 16'h00AF; #100;
A = 16'h0036; B = 16'h00B0; #100;
A = 16'h0036; B = 16'h00B1; #100;
A = 16'h0036; B = 16'h00B2; #100;
A = 16'h0036; B = 16'h00B3; #100;
A = 16'h0036; B = 16'h00B4; #100;
A = 16'h0036; B = 16'h00B5; #100;
A = 16'h0036; B = 16'h00B6; #100;
A = 16'h0036; B = 16'h00B7; #100;
A = 16'h0036; B = 16'h00B8; #100;
A = 16'h0036; B = 16'h00B9; #100;
A = 16'h0036; B = 16'h00BA; #100;
A = 16'h0036; B = 16'h00BB; #100;
A = 16'h0036; B = 16'h00BC; #100;
A = 16'h0036; B = 16'h00BD; #100;
A = 16'h0036; B = 16'h00BE; #100;
A = 16'h0036; B = 16'h00BF; #100;
A = 16'h0036; B = 16'h00C0; #100;
A = 16'h0036; B = 16'h00C1; #100;
A = 16'h0036; B = 16'h00C2; #100;
A = 16'h0036; B = 16'h00C3; #100;
A = 16'h0036; B = 16'h00C4; #100;
A = 16'h0036; B = 16'h00C5; #100;
A = 16'h0036; B = 16'h00C6; #100;
A = 16'h0036; B = 16'h00C7; #100;
A = 16'h0036; B = 16'h00C8; #100;
A = 16'h0036; B = 16'h00C9; #100;
A = 16'h0036; B = 16'h00CA; #100;
A = 16'h0036; B = 16'h00CB; #100;
A = 16'h0036; B = 16'h00CC; #100;
A = 16'h0036; B = 16'h00CD; #100;
A = 16'h0036; B = 16'h00CE; #100;
A = 16'h0036; B = 16'h00CF; #100;
A = 16'h0036; B = 16'h00D0; #100;
A = 16'h0036; B = 16'h00D1; #100;
A = 16'h0036; B = 16'h00D2; #100;
A = 16'h0036; B = 16'h00D3; #100;
A = 16'h0036; B = 16'h00D4; #100;
A = 16'h0036; B = 16'h00D5; #100;
A = 16'h0036; B = 16'h00D6; #100;
A = 16'h0036; B = 16'h00D7; #100;
A = 16'h0036; B = 16'h00D8; #100;
A = 16'h0036; B = 16'h00D9; #100;
A = 16'h0036; B = 16'h00DA; #100;
A = 16'h0036; B = 16'h00DB; #100;
A = 16'h0036; B = 16'h00DC; #100;
A = 16'h0036; B = 16'h00DD; #100;
A = 16'h0036; B = 16'h00DE; #100;
A = 16'h0036; B = 16'h00DF; #100;
A = 16'h0036; B = 16'h00E0; #100;
A = 16'h0036; B = 16'h00E1; #100;
A = 16'h0036; B = 16'h00E2; #100;
A = 16'h0036; B = 16'h00E3; #100;
A = 16'h0036; B = 16'h00E4; #100;
A = 16'h0036; B = 16'h00E5; #100;
A = 16'h0036; B = 16'h00E6; #100;
A = 16'h0036; B = 16'h00E7; #100;
A = 16'h0036; B = 16'h00E8; #100;
A = 16'h0036; B = 16'h00E9; #100;
A = 16'h0036; B = 16'h00EA; #100;
A = 16'h0036; B = 16'h00EB; #100;
A = 16'h0036; B = 16'h00EC; #100;
A = 16'h0036; B = 16'h00ED; #100;
A = 16'h0036; B = 16'h00EE; #100;
A = 16'h0036; B = 16'h00EF; #100;
A = 16'h0036; B = 16'h00F0; #100;
A = 16'h0036; B = 16'h00F1; #100;
A = 16'h0036; B = 16'h00F2; #100;
A = 16'h0036; B = 16'h00F3; #100;
A = 16'h0036; B = 16'h00F4; #100;
A = 16'h0036; B = 16'h00F5; #100;
A = 16'h0036; B = 16'h00F6; #100;
A = 16'h0036; B = 16'h00F7; #100;
A = 16'h0036; B = 16'h00F8; #100;
A = 16'h0036; B = 16'h00F9; #100;
A = 16'h0036; B = 16'h00FA; #100;
A = 16'h0036; B = 16'h00FB; #100;
A = 16'h0036; B = 16'h00FC; #100;
A = 16'h0036; B = 16'h00FD; #100;
A = 16'h0036; B = 16'h00FE; #100;
A = 16'h0036; B = 16'h00FF; #100;
A = 16'h0037; B = 16'h000; #100;
A = 16'h0037; B = 16'h001; #100;
A = 16'h0037; B = 16'h002; #100;
A = 16'h0037; B = 16'h003; #100;
A = 16'h0037; B = 16'h004; #100;
A = 16'h0037; B = 16'h005; #100;
A = 16'h0037; B = 16'h006; #100;
A = 16'h0037; B = 16'h007; #100;
A = 16'h0037; B = 16'h008; #100;
A = 16'h0037; B = 16'h009; #100;
A = 16'h0037; B = 16'h00A; #100;
A = 16'h0037; B = 16'h00B; #100;
A = 16'h0037; B = 16'h00C; #100;
A = 16'h0037; B = 16'h00D; #100;
A = 16'h0037; B = 16'h00E; #100;
A = 16'h0037; B = 16'h00F; #100;
A = 16'h0037; B = 16'h0010; #100;
A = 16'h0037; B = 16'h0011; #100;
A = 16'h0037; B = 16'h0012; #100;
A = 16'h0037; B = 16'h0013; #100;
A = 16'h0037; B = 16'h0014; #100;
A = 16'h0037; B = 16'h0015; #100;
A = 16'h0037; B = 16'h0016; #100;
A = 16'h0037; B = 16'h0017; #100;
A = 16'h0037; B = 16'h0018; #100;
A = 16'h0037; B = 16'h0019; #100;
A = 16'h0037; B = 16'h001A; #100;
A = 16'h0037; B = 16'h001B; #100;
A = 16'h0037; B = 16'h001C; #100;
A = 16'h0037; B = 16'h001D; #100;
A = 16'h0037; B = 16'h001E; #100;
A = 16'h0037; B = 16'h001F; #100;
A = 16'h0037; B = 16'h0020; #100;
A = 16'h0037; B = 16'h0021; #100;
A = 16'h0037; B = 16'h0022; #100;
A = 16'h0037; B = 16'h0023; #100;
A = 16'h0037; B = 16'h0024; #100;
A = 16'h0037; B = 16'h0025; #100;
A = 16'h0037; B = 16'h0026; #100;
A = 16'h0037; B = 16'h0027; #100;
A = 16'h0037; B = 16'h0028; #100;
A = 16'h0037; B = 16'h0029; #100;
A = 16'h0037; B = 16'h002A; #100;
A = 16'h0037; B = 16'h002B; #100;
A = 16'h0037; B = 16'h002C; #100;
A = 16'h0037; B = 16'h002D; #100;
A = 16'h0037; B = 16'h002E; #100;
A = 16'h0037; B = 16'h002F; #100;
A = 16'h0037; B = 16'h0030; #100;
A = 16'h0037; B = 16'h0031; #100;
A = 16'h0037; B = 16'h0032; #100;
A = 16'h0037; B = 16'h0033; #100;
A = 16'h0037; B = 16'h0034; #100;
A = 16'h0037; B = 16'h0035; #100;
A = 16'h0037; B = 16'h0036; #100;
A = 16'h0037; B = 16'h0037; #100;
A = 16'h0037; B = 16'h0038; #100;
A = 16'h0037; B = 16'h0039; #100;
A = 16'h0037; B = 16'h003A; #100;
A = 16'h0037; B = 16'h003B; #100;
A = 16'h0037; B = 16'h003C; #100;
A = 16'h0037; B = 16'h003D; #100;
A = 16'h0037; B = 16'h003E; #100;
A = 16'h0037; B = 16'h003F; #100;
A = 16'h0037; B = 16'h0040; #100;
A = 16'h0037; B = 16'h0041; #100;
A = 16'h0037; B = 16'h0042; #100;
A = 16'h0037; B = 16'h0043; #100;
A = 16'h0037; B = 16'h0044; #100;
A = 16'h0037; B = 16'h0045; #100;
A = 16'h0037; B = 16'h0046; #100;
A = 16'h0037; B = 16'h0047; #100;
A = 16'h0037; B = 16'h0048; #100;
A = 16'h0037; B = 16'h0049; #100;
A = 16'h0037; B = 16'h004A; #100;
A = 16'h0037; B = 16'h004B; #100;
A = 16'h0037; B = 16'h004C; #100;
A = 16'h0037; B = 16'h004D; #100;
A = 16'h0037; B = 16'h004E; #100;
A = 16'h0037; B = 16'h004F; #100;
A = 16'h0037; B = 16'h0050; #100;
A = 16'h0037; B = 16'h0051; #100;
A = 16'h0037; B = 16'h0052; #100;
A = 16'h0037; B = 16'h0053; #100;
A = 16'h0037; B = 16'h0054; #100;
A = 16'h0037; B = 16'h0055; #100;
A = 16'h0037; B = 16'h0056; #100;
A = 16'h0037; B = 16'h0057; #100;
A = 16'h0037; B = 16'h0058; #100;
A = 16'h0037; B = 16'h0059; #100;
A = 16'h0037; B = 16'h005A; #100;
A = 16'h0037; B = 16'h005B; #100;
A = 16'h0037; B = 16'h005C; #100;
A = 16'h0037; B = 16'h005D; #100;
A = 16'h0037; B = 16'h005E; #100;
A = 16'h0037; B = 16'h005F; #100;
A = 16'h0037; B = 16'h0060; #100;
A = 16'h0037; B = 16'h0061; #100;
A = 16'h0037; B = 16'h0062; #100;
A = 16'h0037; B = 16'h0063; #100;
A = 16'h0037; B = 16'h0064; #100;
A = 16'h0037; B = 16'h0065; #100;
A = 16'h0037; B = 16'h0066; #100;
A = 16'h0037; B = 16'h0067; #100;
A = 16'h0037; B = 16'h0068; #100;
A = 16'h0037; B = 16'h0069; #100;
A = 16'h0037; B = 16'h006A; #100;
A = 16'h0037; B = 16'h006B; #100;
A = 16'h0037; B = 16'h006C; #100;
A = 16'h0037; B = 16'h006D; #100;
A = 16'h0037; B = 16'h006E; #100;
A = 16'h0037; B = 16'h006F; #100;
A = 16'h0037; B = 16'h0070; #100;
A = 16'h0037; B = 16'h0071; #100;
A = 16'h0037; B = 16'h0072; #100;
A = 16'h0037; B = 16'h0073; #100;
A = 16'h0037; B = 16'h0074; #100;
A = 16'h0037; B = 16'h0075; #100;
A = 16'h0037; B = 16'h0076; #100;
A = 16'h0037; B = 16'h0077; #100;
A = 16'h0037; B = 16'h0078; #100;
A = 16'h0037; B = 16'h0079; #100;
A = 16'h0037; B = 16'h007A; #100;
A = 16'h0037; B = 16'h007B; #100;
A = 16'h0037; B = 16'h007C; #100;
A = 16'h0037; B = 16'h007D; #100;
A = 16'h0037; B = 16'h007E; #100;
A = 16'h0037; B = 16'h007F; #100;
A = 16'h0037; B = 16'h0080; #100;
A = 16'h0037; B = 16'h0081; #100;
A = 16'h0037; B = 16'h0082; #100;
A = 16'h0037; B = 16'h0083; #100;
A = 16'h0037; B = 16'h0084; #100;
A = 16'h0037; B = 16'h0085; #100;
A = 16'h0037; B = 16'h0086; #100;
A = 16'h0037; B = 16'h0087; #100;
A = 16'h0037; B = 16'h0088; #100;
A = 16'h0037; B = 16'h0089; #100;
A = 16'h0037; B = 16'h008A; #100;
A = 16'h0037; B = 16'h008B; #100;
A = 16'h0037; B = 16'h008C; #100;
A = 16'h0037; B = 16'h008D; #100;
A = 16'h0037; B = 16'h008E; #100;
A = 16'h0037; B = 16'h008F; #100;
A = 16'h0037; B = 16'h0090; #100;
A = 16'h0037; B = 16'h0091; #100;
A = 16'h0037; B = 16'h0092; #100;
A = 16'h0037; B = 16'h0093; #100;
A = 16'h0037; B = 16'h0094; #100;
A = 16'h0037; B = 16'h0095; #100;
A = 16'h0037; B = 16'h0096; #100;
A = 16'h0037; B = 16'h0097; #100;
A = 16'h0037; B = 16'h0098; #100;
A = 16'h0037; B = 16'h0099; #100;
A = 16'h0037; B = 16'h009A; #100;
A = 16'h0037; B = 16'h009B; #100;
A = 16'h0037; B = 16'h009C; #100;
A = 16'h0037; B = 16'h009D; #100;
A = 16'h0037; B = 16'h009E; #100;
A = 16'h0037; B = 16'h009F; #100;
A = 16'h0037; B = 16'h00A0; #100;
A = 16'h0037; B = 16'h00A1; #100;
A = 16'h0037; B = 16'h00A2; #100;
A = 16'h0037; B = 16'h00A3; #100;
A = 16'h0037; B = 16'h00A4; #100;
A = 16'h0037; B = 16'h00A5; #100;
A = 16'h0037; B = 16'h00A6; #100;
A = 16'h0037; B = 16'h00A7; #100;
A = 16'h0037; B = 16'h00A8; #100;
A = 16'h0037; B = 16'h00A9; #100;
A = 16'h0037; B = 16'h00AA; #100;
A = 16'h0037; B = 16'h00AB; #100;
A = 16'h0037; B = 16'h00AC; #100;
A = 16'h0037; B = 16'h00AD; #100;
A = 16'h0037; B = 16'h00AE; #100;
A = 16'h0037; B = 16'h00AF; #100;
A = 16'h0037; B = 16'h00B0; #100;
A = 16'h0037; B = 16'h00B1; #100;
A = 16'h0037; B = 16'h00B2; #100;
A = 16'h0037; B = 16'h00B3; #100;
A = 16'h0037; B = 16'h00B4; #100;
A = 16'h0037; B = 16'h00B5; #100;
A = 16'h0037; B = 16'h00B6; #100;
A = 16'h0037; B = 16'h00B7; #100;
A = 16'h0037; B = 16'h00B8; #100;
A = 16'h0037; B = 16'h00B9; #100;
A = 16'h0037; B = 16'h00BA; #100;
A = 16'h0037; B = 16'h00BB; #100;
A = 16'h0037; B = 16'h00BC; #100;
A = 16'h0037; B = 16'h00BD; #100;
A = 16'h0037; B = 16'h00BE; #100;
A = 16'h0037; B = 16'h00BF; #100;
A = 16'h0037; B = 16'h00C0; #100;
A = 16'h0037; B = 16'h00C1; #100;
A = 16'h0037; B = 16'h00C2; #100;
A = 16'h0037; B = 16'h00C3; #100;
A = 16'h0037; B = 16'h00C4; #100;
A = 16'h0037; B = 16'h00C5; #100;
A = 16'h0037; B = 16'h00C6; #100;
A = 16'h0037; B = 16'h00C7; #100;
A = 16'h0037; B = 16'h00C8; #100;
A = 16'h0037; B = 16'h00C9; #100;
A = 16'h0037; B = 16'h00CA; #100;
A = 16'h0037; B = 16'h00CB; #100;
A = 16'h0037; B = 16'h00CC; #100;
A = 16'h0037; B = 16'h00CD; #100;
A = 16'h0037; B = 16'h00CE; #100;
A = 16'h0037; B = 16'h00CF; #100;
A = 16'h0037; B = 16'h00D0; #100;
A = 16'h0037; B = 16'h00D1; #100;
A = 16'h0037; B = 16'h00D2; #100;
A = 16'h0037; B = 16'h00D3; #100;
A = 16'h0037; B = 16'h00D4; #100;
A = 16'h0037; B = 16'h00D5; #100;
A = 16'h0037; B = 16'h00D6; #100;
A = 16'h0037; B = 16'h00D7; #100;
A = 16'h0037; B = 16'h00D8; #100;
A = 16'h0037; B = 16'h00D9; #100;
A = 16'h0037; B = 16'h00DA; #100;
A = 16'h0037; B = 16'h00DB; #100;
A = 16'h0037; B = 16'h00DC; #100;
A = 16'h0037; B = 16'h00DD; #100;
A = 16'h0037; B = 16'h00DE; #100;
A = 16'h0037; B = 16'h00DF; #100;
A = 16'h0037; B = 16'h00E0; #100;
A = 16'h0037; B = 16'h00E1; #100;
A = 16'h0037; B = 16'h00E2; #100;
A = 16'h0037; B = 16'h00E3; #100;
A = 16'h0037; B = 16'h00E4; #100;
A = 16'h0037; B = 16'h00E5; #100;
A = 16'h0037; B = 16'h00E6; #100;
A = 16'h0037; B = 16'h00E7; #100;
A = 16'h0037; B = 16'h00E8; #100;
A = 16'h0037; B = 16'h00E9; #100;
A = 16'h0037; B = 16'h00EA; #100;
A = 16'h0037; B = 16'h00EB; #100;
A = 16'h0037; B = 16'h00EC; #100;
A = 16'h0037; B = 16'h00ED; #100;
A = 16'h0037; B = 16'h00EE; #100;
A = 16'h0037; B = 16'h00EF; #100;
A = 16'h0037; B = 16'h00F0; #100;
A = 16'h0037; B = 16'h00F1; #100;
A = 16'h0037; B = 16'h00F2; #100;
A = 16'h0037; B = 16'h00F3; #100;
A = 16'h0037; B = 16'h00F4; #100;
A = 16'h0037; B = 16'h00F5; #100;
A = 16'h0037; B = 16'h00F6; #100;
A = 16'h0037; B = 16'h00F7; #100;
A = 16'h0037; B = 16'h00F8; #100;
A = 16'h0037; B = 16'h00F9; #100;
A = 16'h0037; B = 16'h00FA; #100;
A = 16'h0037; B = 16'h00FB; #100;
A = 16'h0037; B = 16'h00FC; #100;
A = 16'h0037; B = 16'h00FD; #100;
A = 16'h0037; B = 16'h00FE; #100;
A = 16'h0037; B = 16'h00FF; #100;
A = 16'h0038; B = 16'h000; #100;
A = 16'h0038; B = 16'h001; #100;
A = 16'h0038; B = 16'h002; #100;
A = 16'h0038; B = 16'h003; #100;
A = 16'h0038; B = 16'h004; #100;
A = 16'h0038; B = 16'h005; #100;
A = 16'h0038; B = 16'h006; #100;
A = 16'h0038; B = 16'h007; #100;
A = 16'h0038; B = 16'h008; #100;
A = 16'h0038; B = 16'h009; #100;
A = 16'h0038; B = 16'h00A; #100;
A = 16'h0038; B = 16'h00B; #100;
A = 16'h0038; B = 16'h00C; #100;
A = 16'h0038; B = 16'h00D; #100;
A = 16'h0038; B = 16'h00E; #100;
A = 16'h0038; B = 16'h00F; #100;
A = 16'h0038; B = 16'h0010; #100;
A = 16'h0038; B = 16'h0011; #100;
A = 16'h0038; B = 16'h0012; #100;
A = 16'h0038; B = 16'h0013; #100;
A = 16'h0038; B = 16'h0014; #100;
A = 16'h0038; B = 16'h0015; #100;
A = 16'h0038; B = 16'h0016; #100;
A = 16'h0038; B = 16'h0017; #100;
A = 16'h0038; B = 16'h0018; #100;
A = 16'h0038; B = 16'h0019; #100;
A = 16'h0038; B = 16'h001A; #100;
A = 16'h0038; B = 16'h001B; #100;
A = 16'h0038; B = 16'h001C; #100;
A = 16'h0038; B = 16'h001D; #100;
A = 16'h0038; B = 16'h001E; #100;
A = 16'h0038; B = 16'h001F; #100;
A = 16'h0038; B = 16'h0020; #100;
A = 16'h0038; B = 16'h0021; #100;
A = 16'h0038; B = 16'h0022; #100;
A = 16'h0038; B = 16'h0023; #100;
A = 16'h0038; B = 16'h0024; #100;
A = 16'h0038; B = 16'h0025; #100;
A = 16'h0038; B = 16'h0026; #100;
A = 16'h0038; B = 16'h0027; #100;
A = 16'h0038; B = 16'h0028; #100;
A = 16'h0038; B = 16'h0029; #100;
A = 16'h0038; B = 16'h002A; #100;
A = 16'h0038; B = 16'h002B; #100;
A = 16'h0038; B = 16'h002C; #100;
A = 16'h0038; B = 16'h002D; #100;
A = 16'h0038; B = 16'h002E; #100;
A = 16'h0038; B = 16'h002F; #100;
A = 16'h0038; B = 16'h0030; #100;
A = 16'h0038; B = 16'h0031; #100;
A = 16'h0038; B = 16'h0032; #100;
A = 16'h0038; B = 16'h0033; #100;
A = 16'h0038; B = 16'h0034; #100;
A = 16'h0038; B = 16'h0035; #100;
A = 16'h0038; B = 16'h0036; #100;
A = 16'h0038; B = 16'h0037; #100;
A = 16'h0038; B = 16'h0038; #100;
A = 16'h0038; B = 16'h0039; #100;
A = 16'h0038; B = 16'h003A; #100;
A = 16'h0038; B = 16'h003B; #100;
A = 16'h0038; B = 16'h003C; #100;
A = 16'h0038; B = 16'h003D; #100;
A = 16'h0038; B = 16'h003E; #100;
A = 16'h0038; B = 16'h003F; #100;
A = 16'h0038; B = 16'h0040; #100;
A = 16'h0038; B = 16'h0041; #100;
A = 16'h0038; B = 16'h0042; #100;
A = 16'h0038; B = 16'h0043; #100;
A = 16'h0038; B = 16'h0044; #100;
A = 16'h0038; B = 16'h0045; #100;
A = 16'h0038; B = 16'h0046; #100;
A = 16'h0038; B = 16'h0047; #100;
A = 16'h0038; B = 16'h0048; #100;
A = 16'h0038; B = 16'h0049; #100;
A = 16'h0038; B = 16'h004A; #100;
A = 16'h0038; B = 16'h004B; #100;
A = 16'h0038; B = 16'h004C; #100;
A = 16'h0038; B = 16'h004D; #100;
A = 16'h0038; B = 16'h004E; #100;
A = 16'h0038; B = 16'h004F; #100;
A = 16'h0038; B = 16'h0050; #100;
A = 16'h0038; B = 16'h0051; #100;
A = 16'h0038; B = 16'h0052; #100;
A = 16'h0038; B = 16'h0053; #100;
A = 16'h0038; B = 16'h0054; #100;
A = 16'h0038; B = 16'h0055; #100;
A = 16'h0038; B = 16'h0056; #100;
A = 16'h0038; B = 16'h0057; #100;
A = 16'h0038; B = 16'h0058; #100;
A = 16'h0038; B = 16'h0059; #100;
A = 16'h0038; B = 16'h005A; #100;
A = 16'h0038; B = 16'h005B; #100;
A = 16'h0038; B = 16'h005C; #100;
A = 16'h0038; B = 16'h005D; #100;
A = 16'h0038; B = 16'h005E; #100;
A = 16'h0038; B = 16'h005F; #100;
A = 16'h0038; B = 16'h0060; #100;
A = 16'h0038; B = 16'h0061; #100;
A = 16'h0038; B = 16'h0062; #100;
A = 16'h0038; B = 16'h0063; #100;
A = 16'h0038; B = 16'h0064; #100;
A = 16'h0038; B = 16'h0065; #100;
A = 16'h0038; B = 16'h0066; #100;
A = 16'h0038; B = 16'h0067; #100;
A = 16'h0038; B = 16'h0068; #100;
A = 16'h0038; B = 16'h0069; #100;
A = 16'h0038; B = 16'h006A; #100;
A = 16'h0038; B = 16'h006B; #100;
A = 16'h0038; B = 16'h006C; #100;
A = 16'h0038; B = 16'h006D; #100;
A = 16'h0038; B = 16'h006E; #100;
A = 16'h0038; B = 16'h006F; #100;
A = 16'h0038; B = 16'h0070; #100;
A = 16'h0038; B = 16'h0071; #100;
A = 16'h0038; B = 16'h0072; #100;
A = 16'h0038; B = 16'h0073; #100;
A = 16'h0038; B = 16'h0074; #100;
A = 16'h0038; B = 16'h0075; #100;
A = 16'h0038; B = 16'h0076; #100;
A = 16'h0038; B = 16'h0077; #100;
A = 16'h0038; B = 16'h0078; #100;
A = 16'h0038; B = 16'h0079; #100;
A = 16'h0038; B = 16'h007A; #100;
A = 16'h0038; B = 16'h007B; #100;
A = 16'h0038; B = 16'h007C; #100;
A = 16'h0038; B = 16'h007D; #100;
A = 16'h0038; B = 16'h007E; #100;
A = 16'h0038; B = 16'h007F; #100;
A = 16'h0038; B = 16'h0080; #100;
A = 16'h0038; B = 16'h0081; #100;
A = 16'h0038; B = 16'h0082; #100;
A = 16'h0038; B = 16'h0083; #100;
A = 16'h0038; B = 16'h0084; #100;
A = 16'h0038; B = 16'h0085; #100;
A = 16'h0038; B = 16'h0086; #100;
A = 16'h0038; B = 16'h0087; #100;
A = 16'h0038; B = 16'h0088; #100;
A = 16'h0038; B = 16'h0089; #100;
A = 16'h0038; B = 16'h008A; #100;
A = 16'h0038; B = 16'h008B; #100;
A = 16'h0038; B = 16'h008C; #100;
A = 16'h0038; B = 16'h008D; #100;
A = 16'h0038; B = 16'h008E; #100;
A = 16'h0038; B = 16'h008F; #100;
A = 16'h0038; B = 16'h0090; #100;
A = 16'h0038; B = 16'h0091; #100;
A = 16'h0038; B = 16'h0092; #100;
A = 16'h0038; B = 16'h0093; #100;
A = 16'h0038; B = 16'h0094; #100;
A = 16'h0038; B = 16'h0095; #100;
A = 16'h0038; B = 16'h0096; #100;
A = 16'h0038; B = 16'h0097; #100;
A = 16'h0038; B = 16'h0098; #100;
A = 16'h0038; B = 16'h0099; #100;
A = 16'h0038; B = 16'h009A; #100;
A = 16'h0038; B = 16'h009B; #100;
A = 16'h0038; B = 16'h009C; #100;
A = 16'h0038; B = 16'h009D; #100;
A = 16'h0038; B = 16'h009E; #100;
A = 16'h0038; B = 16'h009F; #100;
A = 16'h0038; B = 16'h00A0; #100;
A = 16'h0038; B = 16'h00A1; #100;
A = 16'h0038; B = 16'h00A2; #100;
A = 16'h0038; B = 16'h00A3; #100;
A = 16'h0038; B = 16'h00A4; #100;
A = 16'h0038; B = 16'h00A5; #100;
A = 16'h0038; B = 16'h00A6; #100;
A = 16'h0038; B = 16'h00A7; #100;
A = 16'h0038; B = 16'h00A8; #100;
A = 16'h0038; B = 16'h00A9; #100;
A = 16'h0038; B = 16'h00AA; #100;
A = 16'h0038; B = 16'h00AB; #100;
A = 16'h0038; B = 16'h00AC; #100;
A = 16'h0038; B = 16'h00AD; #100;
A = 16'h0038; B = 16'h00AE; #100;
A = 16'h0038; B = 16'h00AF; #100;
A = 16'h0038; B = 16'h00B0; #100;
A = 16'h0038; B = 16'h00B1; #100;
A = 16'h0038; B = 16'h00B2; #100;
A = 16'h0038; B = 16'h00B3; #100;
A = 16'h0038; B = 16'h00B4; #100;
A = 16'h0038; B = 16'h00B5; #100;
A = 16'h0038; B = 16'h00B6; #100;
A = 16'h0038; B = 16'h00B7; #100;
A = 16'h0038; B = 16'h00B8; #100;
A = 16'h0038; B = 16'h00B9; #100;
A = 16'h0038; B = 16'h00BA; #100;
A = 16'h0038; B = 16'h00BB; #100;
A = 16'h0038; B = 16'h00BC; #100;
A = 16'h0038; B = 16'h00BD; #100;
A = 16'h0038; B = 16'h00BE; #100;
A = 16'h0038; B = 16'h00BF; #100;
A = 16'h0038; B = 16'h00C0; #100;
A = 16'h0038; B = 16'h00C1; #100;
A = 16'h0038; B = 16'h00C2; #100;
A = 16'h0038; B = 16'h00C3; #100;
A = 16'h0038; B = 16'h00C4; #100;
A = 16'h0038; B = 16'h00C5; #100;
A = 16'h0038; B = 16'h00C6; #100;
A = 16'h0038; B = 16'h00C7; #100;
A = 16'h0038; B = 16'h00C8; #100;
A = 16'h0038; B = 16'h00C9; #100;
A = 16'h0038; B = 16'h00CA; #100;
A = 16'h0038; B = 16'h00CB; #100;
A = 16'h0038; B = 16'h00CC; #100;
A = 16'h0038; B = 16'h00CD; #100;
A = 16'h0038; B = 16'h00CE; #100;
A = 16'h0038; B = 16'h00CF; #100;
A = 16'h0038; B = 16'h00D0; #100;
A = 16'h0038; B = 16'h00D1; #100;
A = 16'h0038; B = 16'h00D2; #100;
A = 16'h0038; B = 16'h00D3; #100;
A = 16'h0038; B = 16'h00D4; #100;
A = 16'h0038; B = 16'h00D5; #100;
A = 16'h0038; B = 16'h00D6; #100;
A = 16'h0038; B = 16'h00D7; #100;
A = 16'h0038; B = 16'h00D8; #100;
A = 16'h0038; B = 16'h00D9; #100;
A = 16'h0038; B = 16'h00DA; #100;
A = 16'h0038; B = 16'h00DB; #100;
A = 16'h0038; B = 16'h00DC; #100;
A = 16'h0038; B = 16'h00DD; #100;
A = 16'h0038; B = 16'h00DE; #100;
A = 16'h0038; B = 16'h00DF; #100;
A = 16'h0038; B = 16'h00E0; #100;
A = 16'h0038; B = 16'h00E1; #100;
A = 16'h0038; B = 16'h00E2; #100;
A = 16'h0038; B = 16'h00E3; #100;
A = 16'h0038; B = 16'h00E4; #100;
A = 16'h0038; B = 16'h00E5; #100;
A = 16'h0038; B = 16'h00E6; #100;
A = 16'h0038; B = 16'h00E7; #100;
A = 16'h0038; B = 16'h00E8; #100;
A = 16'h0038; B = 16'h00E9; #100;
A = 16'h0038; B = 16'h00EA; #100;
A = 16'h0038; B = 16'h00EB; #100;
A = 16'h0038; B = 16'h00EC; #100;
A = 16'h0038; B = 16'h00ED; #100;
A = 16'h0038; B = 16'h00EE; #100;
A = 16'h0038; B = 16'h00EF; #100;
A = 16'h0038; B = 16'h00F0; #100;
A = 16'h0038; B = 16'h00F1; #100;
A = 16'h0038; B = 16'h00F2; #100;
A = 16'h0038; B = 16'h00F3; #100;
A = 16'h0038; B = 16'h00F4; #100;
A = 16'h0038; B = 16'h00F5; #100;
A = 16'h0038; B = 16'h00F6; #100;
A = 16'h0038; B = 16'h00F7; #100;
A = 16'h0038; B = 16'h00F8; #100;
A = 16'h0038; B = 16'h00F9; #100;
A = 16'h0038; B = 16'h00FA; #100;
A = 16'h0038; B = 16'h00FB; #100;
A = 16'h0038; B = 16'h00FC; #100;
A = 16'h0038; B = 16'h00FD; #100;
A = 16'h0038; B = 16'h00FE; #100;
A = 16'h0038; B = 16'h00FF; #100;
A = 16'h0039; B = 16'h000; #100;
A = 16'h0039; B = 16'h001; #100;
A = 16'h0039; B = 16'h002; #100;
A = 16'h0039; B = 16'h003; #100;
A = 16'h0039; B = 16'h004; #100;
A = 16'h0039; B = 16'h005; #100;
A = 16'h0039; B = 16'h006; #100;
A = 16'h0039; B = 16'h007; #100;
A = 16'h0039; B = 16'h008; #100;
A = 16'h0039; B = 16'h009; #100;
A = 16'h0039; B = 16'h00A; #100;
A = 16'h0039; B = 16'h00B; #100;
A = 16'h0039; B = 16'h00C; #100;
A = 16'h0039; B = 16'h00D; #100;
A = 16'h0039; B = 16'h00E; #100;
A = 16'h0039; B = 16'h00F; #100;
A = 16'h0039; B = 16'h0010; #100;
A = 16'h0039; B = 16'h0011; #100;
A = 16'h0039; B = 16'h0012; #100;
A = 16'h0039; B = 16'h0013; #100;
A = 16'h0039; B = 16'h0014; #100;
A = 16'h0039; B = 16'h0015; #100;
A = 16'h0039; B = 16'h0016; #100;
A = 16'h0039; B = 16'h0017; #100;
A = 16'h0039; B = 16'h0018; #100;
A = 16'h0039; B = 16'h0019; #100;
A = 16'h0039; B = 16'h001A; #100;
A = 16'h0039; B = 16'h001B; #100;
A = 16'h0039; B = 16'h001C; #100;
A = 16'h0039; B = 16'h001D; #100;
A = 16'h0039; B = 16'h001E; #100;
A = 16'h0039; B = 16'h001F; #100;
A = 16'h0039; B = 16'h0020; #100;
A = 16'h0039; B = 16'h0021; #100;
A = 16'h0039; B = 16'h0022; #100;
A = 16'h0039; B = 16'h0023; #100;
A = 16'h0039; B = 16'h0024; #100;
A = 16'h0039; B = 16'h0025; #100;
A = 16'h0039; B = 16'h0026; #100;
A = 16'h0039; B = 16'h0027; #100;
A = 16'h0039; B = 16'h0028; #100;
A = 16'h0039; B = 16'h0029; #100;
A = 16'h0039; B = 16'h002A; #100;
A = 16'h0039; B = 16'h002B; #100;
A = 16'h0039; B = 16'h002C; #100;
A = 16'h0039; B = 16'h002D; #100;
A = 16'h0039; B = 16'h002E; #100;
A = 16'h0039; B = 16'h002F; #100;
A = 16'h0039; B = 16'h0030; #100;
A = 16'h0039; B = 16'h0031; #100;
A = 16'h0039; B = 16'h0032; #100;
A = 16'h0039; B = 16'h0033; #100;
A = 16'h0039; B = 16'h0034; #100;
A = 16'h0039; B = 16'h0035; #100;
A = 16'h0039; B = 16'h0036; #100;
A = 16'h0039; B = 16'h0037; #100;
A = 16'h0039; B = 16'h0038; #100;
A = 16'h0039; B = 16'h0039; #100;
A = 16'h0039; B = 16'h003A; #100;
A = 16'h0039; B = 16'h003B; #100;
A = 16'h0039; B = 16'h003C; #100;
A = 16'h0039; B = 16'h003D; #100;
A = 16'h0039; B = 16'h003E; #100;
A = 16'h0039; B = 16'h003F; #100;
A = 16'h0039; B = 16'h0040; #100;
A = 16'h0039; B = 16'h0041; #100;
A = 16'h0039; B = 16'h0042; #100;
A = 16'h0039; B = 16'h0043; #100;
A = 16'h0039; B = 16'h0044; #100;
A = 16'h0039; B = 16'h0045; #100;
A = 16'h0039; B = 16'h0046; #100;
A = 16'h0039; B = 16'h0047; #100;
A = 16'h0039; B = 16'h0048; #100;
A = 16'h0039; B = 16'h0049; #100;
A = 16'h0039; B = 16'h004A; #100;
A = 16'h0039; B = 16'h004B; #100;
A = 16'h0039; B = 16'h004C; #100;
A = 16'h0039; B = 16'h004D; #100;
A = 16'h0039; B = 16'h004E; #100;
A = 16'h0039; B = 16'h004F; #100;
A = 16'h0039; B = 16'h0050; #100;
A = 16'h0039; B = 16'h0051; #100;
A = 16'h0039; B = 16'h0052; #100;
A = 16'h0039; B = 16'h0053; #100;
A = 16'h0039; B = 16'h0054; #100;
A = 16'h0039; B = 16'h0055; #100;
A = 16'h0039; B = 16'h0056; #100;
A = 16'h0039; B = 16'h0057; #100;
A = 16'h0039; B = 16'h0058; #100;
A = 16'h0039; B = 16'h0059; #100;
A = 16'h0039; B = 16'h005A; #100;
A = 16'h0039; B = 16'h005B; #100;
A = 16'h0039; B = 16'h005C; #100;
A = 16'h0039; B = 16'h005D; #100;
A = 16'h0039; B = 16'h005E; #100;
A = 16'h0039; B = 16'h005F; #100;
A = 16'h0039; B = 16'h0060; #100;
A = 16'h0039; B = 16'h0061; #100;
A = 16'h0039; B = 16'h0062; #100;
A = 16'h0039; B = 16'h0063; #100;
A = 16'h0039; B = 16'h0064; #100;
A = 16'h0039; B = 16'h0065; #100;
A = 16'h0039; B = 16'h0066; #100;
A = 16'h0039; B = 16'h0067; #100;
A = 16'h0039; B = 16'h0068; #100;
A = 16'h0039; B = 16'h0069; #100;
A = 16'h0039; B = 16'h006A; #100;
A = 16'h0039; B = 16'h006B; #100;
A = 16'h0039; B = 16'h006C; #100;
A = 16'h0039; B = 16'h006D; #100;
A = 16'h0039; B = 16'h006E; #100;
A = 16'h0039; B = 16'h006F; #100;
A = 16'h0039; B = 16'h0070; #100;
A = 16'h0039; B = 16'h0071; #100;
A = 16'h0039; B = 16'h0072; #100;
A = 16'h0039; B = 16'h0073; #100;
A = 16'h0039; B = 16'h0074; #100;
A = 16'h0039; B = 16'h0075; #100;
A = 16'h0039; B = 16'h0076; #100;
A = 16'h0039; B = 16'h0077; #100;
A = 16'h0039; B = 16'h0078; #100;
A = 16'h0039; B = 16'h0079; #100;
A = 16'h0039; B = 16'h007A; #100;
A = 16'h0039; B = 16'h007B; #100;
A = 16'h0039; B = 16'h007C; #100;
A = 16'h0039; B = 16'h007D; #100;
A = 16'h0039; B = 16'h007E; #100;
A = 16'h0039; B = 16'h007F; #100;
A = 16'h0039; B = 16'h0080; #100;
A = 16'h0039; B = 16'h0081; #100;
A = 16'h0039; B = 16'h0082; #100;
A = 16'h0039; B = 16'h0083; #100;
A = 16'h0039; B = 16'h0084; #100;
A = 16'h0039; B = 16'h0085; #100;
A = 16'h0039; B = 16'h0086; #100;
A = 16'h0039; B = 16'h0087; #100;
A = 16'h0039; B = 16'h0088; #100;
A = 16'h0039; B = 16'h0089; #100;
A = 16'h0039; B = 16'h008A; #100;
A = 16'h0039; B = 16'h008B; #100;
A = 16'h0039; B = 16'h008C; #100;
A = 16'h0039; B = 16'h008D; #100;
A = 16'h0039; B = 16'h008E; #100;
A = 16'h0039; B = 16'h008F; #100;
A = 16'h0039; B = 16'h0090; #100;
A = 16'h0039; B = 16'h0091; #100;
A = 16'h0039; B = 16'h0092; #100;
A = 16'h0039; B = 16'h0093; #100;
A = 16'h0039; B = 16'h0094; #100;
A = 16'h0039; B = 16'h0095; #100;
A = 16'h0039; B = 16'h0096; #100;
A = 16'h0039; B = 16'h0097; #100;
A = 16'h0039; B = 16'h0098; #100;
A = 16'h0039; B = 16'h0099; #100;
A = 16'h0039; B = 16'h009A; #100;
A = 16'h0039; B = 16'h009B; #100;
A = 16'h0039; B = 16'h009C; #100;
A = 16'h0039; B = 16'h009D; #100;
A = 16'h0039; B = 16'h009E; #100;
A = 16'h0039; B = 16'h009F; #100;
A = 16'h0039; B = 16'h00A0; #100;
A = 16'h0039; B = 16'h00A1; #100;
A = 16'h0039; B = 16'h00A2; #100;
A = 16'h0039; B = 16'h00A3; #100;
A = 16'h0039; B = 16'h00A4; #100;
A = 16'h0039; B = 16'h00A5; #100;
A = 16'h0039; B = 16'h00A6; #100;
A = 16'h0039; B = 16'h00A7; #100;
A = 16'h0039; B = 16'h00A8; #100;
A = 16'h0039; B = 16'h00A9; #100;
A = 16'h0039; B = 16'h00AA; #100;
A = 16'h0039; B = 16'h00AB; #100;
A = 16'h0039; B = 16'h00AC; #100;
A = 16'h0039; B = 16'h00AD; #100;
A = 16'h0039; B = 16'h00AE; #100;
A = 16'h0039; B = 16'h00AF; #100;
A = 16'h0039; B = 16'h00B0; #100;
A = 16'h0039; B = 16'h00B1; #100;
A = 16'h0039; B = 16'h00B2; #100;
A = 16'h0039; B = 16'h00B3; #100;
A = 16'h0039; B = 16'h00B4; #100;
A = 16'h0039; B = 16'h00B5; #100;
A = 16'h0039; B = 16'h00B6; #100;
A = 16'h0039; B = 16'h00B7; #100;
A = 16'h0039; B = 16'h00B8; #100;
A = 16'h0039; B = 16'h00B9; #100;
A = 16'h0039; B = 16'h00BA; #100;
A = 16'h0039; B = 16'h00BB; #100;
A = 16'h0039; B = 16'h00BC; #100;
A = 16'h0039; B = 16'h00BD; #100;
A = 16'h0039; B = 16'h00BE; #100;
A = 16'h0039; B = 16'h00BF; #100;
A = 16'h0039; B = 16'h00C0; #100;
A = 16'h0039; B = 16'h00C1; #100;
A = 16'h0039; B = 16'h00C2; #100;
A = 16'h0039; B = 16'h00C3; #100;
A = 16'h0039; B = 16'h00C4; #100;
A = 16'h0039; B = 16'h00C5; #100;
A = 16'h0039; B = 16'h00C6; #100;
A = 16'h0039; B = 16'h00C7; #100;
A = 16'h0039; B = 16'h00C8; #100;
A = 16'h0039; B = 16'h00C9; #100;
A = 16'h0039; B = 16'h00CA; #100;
A = 16'h0039; B = 16'h00CB; #100;
A = 16'h0039; B = 16'h00CC; #100;
A = 16'h0039; B = 16'h00CD; #100;
A = 16'h0039; B = 16'h00CE; #100;
A = 16'h0039; B = 16'h00CF; #100;
A = 16'h0039; B = 16'h00D0; #100;
A = 16'h0039; B = 16'h00D1; #100;
A = 16'h0039; B = 16'h00D2; #100;
A = 16'h0039; B = 16'h00D3; #100;
A = 16'h0039; B = 16'h00D4; #100;
A = 16'h0039; B = 16'h00D5; #100;
A = 16'h0039; B = 16'h00D6; #100;
A = 16'h0039; B = 16'h00D7; #100;
A = 16'h0039; B = 16'h00D8; #100;
A = 16'h0039; B = 16'h00D9; #100;
A = 16'h0039; B = 16'h00DA; #100;
A = 16'h0039; B = 16'h00DB; #100;
A = 16'h0039; B = 16'h00DC; #100;
A = 16'h0039; B = 16'h00DD; #100;
A = 16'h0039; B = 16'h00DE; #100;
A = 16'h0039; B = 16'h00DF; #100;
A = 16'h0039; B = 16'h00E0; #100;
A = 16'h0039; B = 16'h00E1; #100;
A = 16'h0039; B = 16'h00E2; #100;
A = 16'h0039; B = 16'h00E3; #100;
A = 16'h0039; B = 16'h00E4; #100;
A = 16'h0039; B = 16'h00E5; #100;
A = 16'h0039; B = 16'h00E6; #100;
A = 16'h0039; B = 16'h00E7; #100;
A = 16'h0039; B = 16'h00E8; #100;
A = 16'h0039; B = 16'h00E9; #100;
A = 16'h0039; B = 16'h00EA; #100;
A = 16'h0039; B = 16'h00EB; #100;
A = 16'h0039; B = 16'h00EC; #100;
A = 16'h0039; B = 16'h00ED; #100;
A = 16'h0039; B = 16'h00EE; #100;
A = 16'h0039; B = 16'h00EF; #100;
A = 16'h0039; B = 16'h00F0; #100;
A = 16'h0039; B = 16'h00F1; #100;
A = 16'h0039; B = 16'h00F2; #100;
A = 16'h0039; B = 16'h00F3; #100;
A = 16'h0039; B = 16'h00F4; #100;
A = 16'h0039; B = 16'h00F5; #100;
A = 16'h0039; B = 16'h00F6; #100;
A = 16'h0039; B = 16'h00F7; #100;
A = 16'h0039; B = 16'h00F8; #100;
A = 16'h0039; B = 16'h00F9; #100;
A = 16'h0039; B = 16'h00FA; #100;
A = 16'h0039; B = 16'h00FB; #100;
A = 16'h0039; B = 16'h00FC; #100;
A = 16'h0039; B = 16'h00FD; #100;
A = 16'h0039; B = 16'h00FE; #100;
A = 16'h0039; B = 16'h00FF; #100;
A = 16'h003A; B = 16'h000; #100;
A = 16'h003A; B = 16'h001; #100;
A = 16'h003A; B = 16'h002; #100;
A = 16'h003A; B = 16'h003; #100;
A = 16'h003A; B = 16'h004; #100;
A = 16'h003A; B = 16'h005; #100;
A = 16'h003A; B = 16'h006; #100;
A = 16'h003A; B = 16'h007; #100;
A = 16'h003A; B = 16'h008; #100;
A = 16'h003A; B = 16'h009; #100;
A = 16'h003A; B = 16'h00A; #100;
A = 16'h003A; B = 16'h00B; #100;
A = 16'h003A; B = 16'h00C; #100;
A = 16'h003A; B = 16'h00D; #100;
A = 16'h003A; B = 16'h00E; #100;
A = 16'h003A; B = 16'h00F; #100;
A = 16'h003A; B = 16'h0010; #100;
A = 16'h003A; B = 16'h0011; #100;
A = 16'h003A; B = 16'h0012; #100;
A = 16'h003A; B = 16'h0013; #100;
A = 16'h003A; B = 16'h0014; #100;
A = 16'h003A; B = 16'h0015; #100;
A = 16'h003A; B = 16'h0016; #100;
A = 16'h003A; B = 16'h0017; #100;
A = 16'h003A; B = 16'h0018; #100;
A = 16'h003A; B = 16'h0019; #100;
A = 16'h003A; B = 16'h001A; #100;
A = 16'h003A; B = 16'h001B; #100;
A = 16'h003A; B = 16'h001C; #100;
A = 16'h003A; B = 16'h001D; #100;
A = 16'h003A; B = 16'h001E; #100;
A = 16'h003A; B = 16'h001F; #100;
A = 16'h003A; B = 16'h0020; #100;
A = 16'h003A; B = 16'h0021; #100;
A = 16'h003A; B = 16'h0022; #100;
A = 16'h003A; B = 16'h0023; #100;
A = 16'h003A; B = 16'h0024; #100;
A = 16'h003A; B = 16'h0025; #100;
A = 16'h003A; B = 16'h0026; #100;
A = 16'h003A; B = 16'h0027; #100;
A = 16'h003A; B = 16'h0028; #100;
A = 16'h003A; B = 16'h0029; #100;
A = 16'h003A; B = 16'h002A; #100;
A = 16'h003A; B = 16'h002B; #100;
A = 16'h003A; B = 16'h002C; #100;
A = 16'h003A; B = 16'h002D; #100;
A = 16'h003A; B = 16'h002E; #100;
A = 16'h003A; B = 16'h002F; #100;
A = 16'h003A; B = 16'h0030; #100;
A = 16'h003A; B = 16'h0031; #100;
A = 16'h003A; B = 16'h0032; #100;
A = 16'h003A; B = 16'h0033; #100;
A = 16'h003A; B = 16'h0034; #100;
A = 16'h003A; B = 16'h0035; #100;
A = 16'h003A; B = 16'h0036; #100;
A = 16'h003A; B = 16'h0037; #100;
A = 16'h003A; B = 16'h0038; #100;
A = 16'h003A; B = 16'h0039; #100;
A = 16'h003A; B = 16'h003A; #100;
A = 16'h003A; B = 16'h003B; #100;
A = 16'h003A; B = 16'h003C; #100;
A = 16'h003A; B = 16'h003D; #100;
A = 16'h003A; B = 16'h003E; #100;
A = 16'h003A; B = 16'h003F; #100;
A = 16'h003A; B = 16'h0040; #100;
A = 16'h003A; B = 16'h0041; #100;
A = 16'h003A; B = 16'h0042; #100;
A = 16'h003A; B = 16'h0043; #100;
A = 16'h003A; B = 16'h0044; #100;
A = 16'h003A; B = 16'h0045; #100;
A = 16'h003A; B = 16'h0046; #100;
A = 16'h003A; B = 16'h0047; #100;
A = 16'h003A; B = 16'h0048; #100;
A = 16'h003A; B = 16'h0049; #100;
A = 16'h003A; B = 16'h004A; #100;
A = 16'h003A; B = 16'h004B; #100;
A = 16'h003A; B = 16'h004C; #100;
A = 16'h003A; B = 16'h004D; #100;
A = 16'h003A; B = 16'h004E; #100;
A = 16'h003A; B = 16'h004F; #100;
A = 16'h003A; B = 16'h0050; #100;
A = 16'h003A; B = 16'h0051; #100;
A = 16'h003A; B = 16'h0052; #100;
A = 16'h003A; B = 16'h0053; #100;
A = 16'h003A; B = 16'h0054; #100;
A = 16'h003A; B = 16'h0055; #100;
A = 16'h003A; B = 16'h0056; #100;
A = 16'h003A; B = 16'h0057; #100;
A = 16'h003A; B = 16'h0058; #100;
A = 16'h003A; B = 16'h0059; #100;
A = 16'h003A; B = 16'h005A; #100;
A = 16'h003A; B = 16'h005B; #100;
A = 16'h003A; B = 16'h005C; #100;
A = 16'h003A; B = 16'h005D; #100;
A = 16'h003A; B = 16'h005E; #100;
A = 16'h003A; B = 16'h005F; #100;
A = 16'h003A; B = 16'h0060; #100;
A = 16'h003A; B = 16'h0061; #100;
A = 16'h003A; B = 16'h0062; #100;
A = 16'h003A; B = 16'h0063; #100;
A = 16'h003A; B = 16'h0064; #100;
A = 16'h003A; B = 16'h0065; #100;
A = 16'h003A; B = 16'h0066; #100;
A = 16'h003A; B = 16'h0067; #100;
A = 16'h003A; B = 16'h0068; #100;
A = 16'h003A; B = 16'h0069; #100;
A = 16'h003A; B = 16'h006A; #100;
A = 16'h003A; B = 16'h006B; #100;
A = 16'h003A; B = 16'h006C; #100;
A = 16'h003A; B = 16'h006D; #100;
A = 16'h003A; B = 16'h006E; #100;
A = 16'h003A; B = 16'h006F; #100;
A = 16'h003A; B = 16'h0070; #100;
A = 16'h003A; B = 16'h0071; #100;
A = 16'h003A; B = 16'h0072; #100;
A = 16'h003A; B = 16'h0073; #100;
A = 16'h003A; B = 16'h0074; #100;
A = 16'h003A; B = 16'h0075; #100;
A = 16'h003A; B = 16'h0076; #100;
A = 16'h003A; B = 16'h0077; #100;
A = 16'h003A; B = 16'h0078; #100;
A = 16'h003A; B = 16'h0079; #100;
A = 16'h003A; B = 16'h007A; #100;
A = 16'h003A; B = 16'h007B; #100;
A = 16'h003A; B = 16'h007C; #100;
A = 16'h003A; B = 16'h007D; #100;
A = 16'h003A; B = 16'h007E; #100;
A = 16'h003A; B = 16'h007F; #100;
A = 16'h003A; B = 16'h0080; #100;
A = 16'h003A; B = 16'h0081; #100;
A = 16'h003A; B = 16'h0082; #100;
A = 16'h003A; B = 16'h0083; #100;
A = 16'h003A; B = 16'h0084; #100;
A = 16'h003A; B = 16'h0085; #100;
A = 16'h003A; B = 16'h0086; #100;
A = 16'h003A; B = 16'h0087; #100;
A = 16'h003A; B = 16'h0088; #100;
A = 16'h003A; B = 16'h0089; #100;
A = 16'h003A; B = 16'h008A; #100;
A = 16'h003A; B = 16'h008B; #100;
A = 16'h003A; B = 16'h008C; #100;
A = 16'h003A; B = 16'h008D; #100;
A = 16'h003A; B = 16'h008E; #100;
A = 16'h003A; B = 16'h008F; #100;
A = 16'h003A; B = 16'h0090; #100;
A = 16'h003A; B = 16'h0091; #100;
A = 16'h003A; B = 16'h0092; #100;
A = 16'h003A; B = 16'h0093; #100;
A = 16'h003A; B = 16'h0094; #100;
A = 16'h003A; B = 16'h0095; #100;
A = 16'h003A; B = 16'h0096; #100;
A = 16'h003A; B = 16'h0097; #100;
A = 16'h003A; B = 16'h0098; #100;
A = 16'h003A; B = 16'h0099; #100;
A = 16'h003A; B = 16'h009A; #100;
A = 16'h003A; B = 16'h009B; #100;
A = 16'h003A; B = 16'h009C; #100;
A = 16'h003A; B = 16'h009D; #100;
A = 16'h003A; B = 16'h009E; #100;
A = 16'h003A; B = 16'h009F; #100;
A = 16'h003A; B = 16'h00A0; #100;
A = 16'h003A; B = 16'h00A1; #100;
A = 16'h003A; B = 16'h00A2; #100;
A = 16'h003A; B = 16'h00A3; #100;
A = 16'h003A; B = 16'h00A4; #100;
A = 16'h003A; B = 16'h00A5; #100;
A = 16'h003A; B = 16'h00A6; #100;
A = 16'h003A; B = 16'h00A7; #100;
A = 16'h003A; B = 16'h00A8; #100;
A = 16'h003A; B = 16'h00A9; #100;
A = 16'h003A; B = 16'h00AA; #100;
A = 16'h003A; B = 16'h00AB; #100;
A = 16'h003A; B = 16'h00AC; #100;
A = 16'h003A; B = 16'h00AD; #100;
A = 16'h003A; B = 16'h00AE; #100;
A = 16'h003A; B = 16'h00AF; #100;
A = 16'h003A; B = 16'h00B0; #100;
A = 16'h003A; B = 16'h00B1; #100;
A = 16'h003A; B = 16'h00B2; #100;
A = 16'h003A; B = 16'h00B3; #100;
A = 16'h003A; B = 16'h00B4; #100;
A = 16'h003A; B = 16'h00B5; #100;
A = 16'h003A; B = 16'h00B6; #100;
A = 16'h003A; B = 16'h00B7; #100;
A = 16'h003A; B = 16'h00B8; #100;
A = 16'h003A; B = 16'h00B9; #100;
A = 16'h003A; B = 16'h00BA; #100;
A = 16'h003A; B = 16'h00BB; #100;
A = 16'h003A; B = 16'h00BC; #100;
A = 16'h003A; B = 16'h00BD; #100;
A = 16'h003A; B = 16'h00BE; #100;
A = 16'h003A; B = 16'h00BF; #100;
A = 16'h003A; B = 16'h00C0; #100;
A = 16'h003A; B = 16'h00C1; #100;
A = 16'h003A; B = 16'h00C2; #100;
A = 16'h003A; B = 16'h00C3; #100;
A = 16'h003A; B = 16'h00C4; #100;
A = 16'h003A; B = 16'h00C5; #100;
A = 16'h003A; B = 16'h00C6; #100;
A = 16'h003A; B = 16'h00C7; #100;
A = 16'h003A; B = 16'h00C8; #100;
A = 16'h003A; B = 16'h00C9; #100;
A = 16'h003A; B = 16'h00CA; #100;
A = 16'h003A; B = 16'h00CB; #100;
A = 16'h003A; B = 16'h00CC; #100;
A = 16'h003A; B = 16'h00CD; #100;
A = 16'h003A; B = 16'h00CE; #100;
A = 16'h003A; B = 16'h00CF; #100;
A = 16'h003A; B = 16'h00D0; #100;
A = 16'h003A; B = 16'h00D1; #100;
A = 16'h003A; B = 16'h00D2; #100;
A = 16'h003A; B = 16'h00D3; #100;
A = 16'h003A; B = 16'h00D4; #100;
A = 16'h003A; B = 16'h00D5; #100;
A = 16'h003A; B = 16'h00D6; #100;
A = 16'h003A; B = 16'h00D7; #100;
A = 16'h003A; B = 16'h00D8; #100;
A = 16'h003A; B = 16'h00D9; #100;
A = 16'h003A; B = 16'h00DA; #100;
A = 16'h003A; B = 16'h00DB; #100;
A = 16'h003A; B = 16'h00DC; #100;
A = 16'h003A; B = 16'h00DD; #100;
A = 16'h003A; B = 16'h00DE; #100;
A = 16'h003A; B = 16'h00DF; #100;
A = 16'h003A; B = 16'h00E0; #100;
A = 16'h003A; B = 16'h00E1; #100;
A = 16'h003A; B = 16'h00E2; #100;
A = 16'h003A; B = 16'h00E3; #100;
A = 16'h003A; B = 16'h00E4; #100;
A = 16'h003A; B = 16'h00E5; #100;
A = 16'h003A; B = 16'h00E6; #100;
A = 16'h003A; B = 16'h00E7; #100;
A = 16'h003A; B = 16'h00E8; #100;
A = 16'h003A; B = 16'h00E9; #100;
A = 16'h003A; B = 16'h00EA; #100;
A = 16'h003A; B = 16'h00EB; #100;
A = 16'h003A; B = 16'h00EC; #100;
A = 16'h003A; B = 16'h00ED; #100;
A = 16'h003A; B = 16'h00EE; #100;
A = 16'h003A; B = 16'h00EF; #100;
A = 16'h003A; B = 16'h00F0; #100;
A = 16'h003A; B = 16'h00F1; #100;
A = 16'h003A; B = 16'h00F2; #100;
A = 16'h003A; B = 16'h00F3; #100;
A = 16'h003A; B = 16'h00F4; #100;
A = 16'h003A; B = 16'h00F5; #100;
A = 16'h003A; B = 16'h00F6; #100;
A = 16'h003A; B = 16'h00F7; #100;
A = 16'h003A; B = 16'h00F8; #100;
A = 16'h003A; B = 16'h00F9; #100;
A = 16'h003A; B = 16'h00FA; #100;
A = 16'h003A; B = 16'h00FB; #100;
A = 16'h003A; B = 16'h00FC; #100;
A = 16'h003A; B = 16'h00FD; #100;
A = 16'h003A; B = 16'h00FE; #100;
A = 16'h003A; B = 16'h00FF; #100;
A = 16'h003B; B = 16'h000; #100;
A = 16'h003B; B = 16'h001; #100;
A = 16'h003B; B = 16'h002; #100;
A = 16'h003B; B = 16'h003; #100;
A = 16'h003B; B = 16'h004; #100;
A = 16'h003B; B = 16'h005; #100;
A = 16'h003B; B = 16'h006; #100;
A = 16'h003B; B = 16'h007; #100;
A = 16'h003B; B = 16'h008; #100;
A = 16'h003B; B = 16'h009; #100;
A = 16'h003B; B = 16'h00A; #100;
A = 16'h003B; B = 16'h00B; #100;
A = 16'h003B; B = 16'h00C; #100;
A = 16'h003B; B = 16'h00D; #100;
A = 16'h003B; B = 16'h00E; #100;
A = 16'h003B; B = 16'h00F; #100;
A = 16'h003B; B = 16'h0010; #100;
A = 16'h003B; B = 16'h0011; #100;
A = 16'h003B; B = 16'h0012; #100;
A = 16'h003B; B = 16'h0013; #100;
A = 16'h003B; B = 16'h0014; #100;
A = 16'h003B; B = 16'h0015; #100;
A = 16'h003B; B = 16'h0016; #100;
A = 16'h003B; B = 16'h0017; #100;
A = 16'h003B; B = 16'h0018; #100;
A = 16'h003B; B = 16'h0019; #100;
A = 16'h003B; B = 16'h001A; #100;
A = 16'h003B; B = 16'h001B; #100;
A = 16'h003B; B = 16'h001C; #100;
A = 16'h003B; B = 16'h001D; #100;
A = 16'h003B; B = 16'h001E; #100;
A = 16'h003B; B = 16'h001F; #100;
A = 16'h003B; B = 16'h0020; #100;
A = 16'h003B; B = 16'h0021; #100;
A = 16'h003B; B = 16'h0022; #100;
A = 16'h003B; B = 16'h0023; #100;
A = 16'h003B; B = 16'h0024; #100;
A = 16'h003B; B = 16'h0025; #100;
A = 16'h003B; B = 16'h0026; #100;
A = 16'h003B; B = 16'h0027; #100;
A = 16'h003B; B = 16'h0028; #100;
A = 16'h003B; B = 16'h0029; #100;
A = 16'h003B; B = 16'h002A; #100;
A = 16'h003B; B = 16'h002B; #100;
A = 16'h003B; B = 16'h002C; #100;
A = 16'h003B; B = 16'h002D; #100;
A = 16'h003B; B = 16'h002E; #100;
A = 16'h003B; B = 16'h002F; #100;
A = 16'h003B; B = 16'h0030; #100;
A = 16'h003B; B = 16'h0031; #100;
A = 16'h003B; B = 16'h0032; #100;
A = 16'h003B; B = 16'h0033; #100;
A = 16'h003B; B = 16'h0034; #100;
A = 16'h003B; B = 16'h0035; #100;
A = 16'h003B; B = 16'h0036; #100;
A = 16'h003B; B = 16'h0037; #100;
A = 16'h003B; B = 16'h0038; #100;
A = 16'h003B; B = 16'h0039; #100;
A = 16'h003B; B = 16'h003A; #100;
A = 16'h003B; B = 16'h003B; #100;
A = 16'h003B; B = 16'h003C; #100;
A = 16'h003B; B = 16'h003D; #100;
A = 16'h003B; B = 16'h003E; #100;
A = 16'h003B; B = 16'h003F; #100;
A = 16'h003B; B = 16'h0040; #100;
A = 16'h003B; B = 16'h0041; #100;
A = 16'h003B; B = 16'h0042; #100;
A = 16'h003B; B = 16'h0043; #100;
A = 16'h003B; B = 16'h0044; #100;
A = 16'h003B; B = 16'h0045; #100;
A = 16'h003B; B = 16'h0046; #100;
A = 16'h003B; B = 16'h0047; #100;
A = 16'h003B; B = 16'h0048; #100;
A = 16'h003B; B = 16'h0049; #100;
A = 16'h003B; B = 16'h004A; #100;
A = 16'h003B; B = 16'h004B; #100;
A = 16'h003B; B = 16'h004C; #100;
A = 16'h003B; B = 16'h004D; #100;
A = 16'h003B; B = 16'h004E; #100;
A = 16'h003B; B = 16'h004F; #100;
A = 16'h003B; B = 16'h0050; #100;
A = 16'h003B; B = 16'h0051; #100;
A = 16'h003B; B = 16'h0052; #100;
A = 16'h003B; B = 16'h0053; #100;
A = 16'h003B; B = 16'h0054; #100;
A = 16'h003B; B = 16'h0055; #100;
A = 16'h003B; B = 16'h0056; #100;
A = 16'h003B; B = 16'h0057; #100;
A = 16'h003B; B = 16'h0058; #100;
A = 16'h003B; B = 16'h0059; #100;
A = 16'h003B; B = 16'h005A; #100;
A = 16'h003B; B = 16'h005B; #100;
A = 16'h003B; B = 16'h005C; #100;
A = 16'h003B; B = 16'h005D; #100;
A = 16'h003B; B = 16'h005E; #100;
A = 16'h003B; B = 16'h005F; #100;
A = 16'h003B; B = 16'h0060; #100;
A = 16'h003B; B = 16'h0061; #100;
A = 16'h003B; B = 16'h0062; #100;
A = 16'h003B; B = 16'h0063; #100;
A = 16'h003B; B = 16'h0064; #100;
A = 16'h003B; B = 16'h0065; #100;
A = 16'h003B; B = 16'h0066; #100;
A = 16'h003B; B = 16'h0067; #100;
A = 16'h003B; B = 16'h0068; #100;
A = 16'h003B; B = 16'h0069; #100;
A = 16'h003B; B = 16'h006A; #100;
A = 16'h003B; B = 16'h006B; #100;
A = 16'h003B; B = 16'h006C; #100;
A = 16'h003B; B = 16'h006D; #100;
A = 16'h003B; B = 16'h006E; #100;
A = 16'h003B; B = 16'h006F; #100;
A = 16'h003B; B = 16'h0070; #100;
A = 16'h003B; B = 16'h0071; #100;
A = 16'h003B; B = 16'h0072; #100;
A = 16'h003B; B = 16'h0073; #100;
A = 16'h003B; B = 16'h0074; #100;
A = 16'h003B; B = 16'h0075; #100;
A = 16'h003B; B = 16'h0076; #100;
A = 16'h003B; B = 16'h0077; #100;
A = 16'h003B; B = 16'h0078; #100;
A = 16'h003B; B = 16'h0079; #100;
A = 16'h003B; B = 16'h007A; #100;
A = 16'h003B; B = 16'h007B; #100;
A = 16'h003B; B = 16'h007C; #100;
A = 16'h003B; B = 16'h007D; #100;
A = 16'h003B; B = 16'h007E; #100;
A = 16'h003B; B = 16'h007F; #100;
A = 16'h003B; B = 16'h0080; #100;
A = 16'h003B; B = 16'h0081; #100;
A = 16'h003B; B = 16'h0082; #100;
A = 16'h003B; B = 16'h0083; #100;
A = 16'h003B; B = 16'h0084; #100;
A = 16'h003B; B = 16'h0085; #100;
A = 16'h003B; B = 16'h0086; #100;
A = 16'h003B; B = 16'h0087; #100;
A = 16'h003B; B = 16'h0088; #100;
A = 16'h003B; B = 16'h0089; #100;
A = 16'h003B; B = 16'h008A; #100;
A = 16'h003B; B = 16'h008B; #100;
A = 16'h003B; B = 16'h008C; #100;
A = 16'h003B; B = 16'h008D; #100;
A = 16'h003B; B = 16'h008E; #100;
A = 16'h003B; B = 16'h008F; #100;
A = 16'h003B; B = 16'h0090; #100;
A = 16'h003B; B = 16'h0091; #100;
A = 16'h003B; B = 16'h0092; #100;
A = 16'h003B; B = 16'h0093; #100;
A = 16'h003B; B = 16'h0094; #100;
A = 16'h003B; B = 16'h0095; #100;
A = 16'h003B; B = 16'h0096; #100;
A = 16'h003B; B = 16'h0097; #100;
A = 16'h003B; B = 16'h0098; #100;
A = 16'h003B; B = 16'h0099; #100;
A = 16'h003B; B = 16'h009A; #100;
A = 16'h003B; B = 16'h009B; #100;
A = 16'h003B; B = 16'h009C; #100;
A = 16'h003B; B = 16'h009D; #100;
A = 16'h003B; B = 16'h009E; #100;
A = 16'h003B; B = 16'h009F; #100;
A = 16'h003B; B = 16'h00A0; #100;
A = 16'h003B; B = 16'h00A1; #100;
A = 16'h003B; B = 16'h00A2; #100;
A = 16'h003B; B = 16'h00A3; #100;
A = 16'h003B; B = 16'h00A4; #100;
A = 16'h003B; B = 16'h00A5; #100;
A = 16'h003B; B = 16'h00A6; #100;
A = 16'h003B; B = 16'h00A7; #100;
A = 16'h003B; B = 16'h00A8; #100;
A = 16'h003B; B = 16'h00A9; #100;
A = 16'h003B; B = 16'h00AA; #100;
A = 16'h003B; B = 16'h00AB; #100;
A = 16'h003B; B = 16'h00AC; #100;
A = 16'h003B; B = 16'h00AD; #100;
A = 16'h003B; B = 16'h00AE; #100;
A = 16'h003B; B = 16'h00AF; #100;
A = 16'h003B; B = 16'h00B0; #100;
A = 16'h003B; B = 16'h00B1; #100;
A = 16'h003B; B = 16'h00B2; #100;
A = 16'h003B; B = 16'h00B3; #100;
A = 16'h003B; B = 16'h00B4; #100;
A = 16'h003B; B = 16'h00B5; #100;
A = 16'h003B; B = 16'h00B6; #100;
A = 16'h003B; B = 16'h00B7; #100;
A = 16'h003B; B = 16'h00B8; #100;
A = 16'h003B; B = 16'h00B9; #100;
A = 16'h003B; B = 16'h00BA; #100;
A = 16'h003B; B = 16'h00BB; #100;
A = 16'h003B; B = 16'h00BC; #100;
A = 16'h003B; B = 16'h00BD; #100;
A = 16'h003B; B = 16'h00BE; #100;
A = 16'h003B; B = 16'h00BF; #100;
A = 16'h003B; B = 16'h00C0; #100;
A = 16'h003B; B = 16'h00C1; #100;
A = 16'h003B; B = 16'h00C2; #100;
A = 16'h003B; B = 16'h00C3; #100;
A = 16'h003B; B = 16'h00C4; #100;
A = 16'h003B; B = 16'h00C5; #100;
A = 16'h003B; B = 16'h00C6; #100;
A = 16'h003B; B = 16'h00C7; #100;
A = 16'h003B; B = 16'h00C8; #100;
A = 16'h003B; B = 16'h00C9; #100;
A = 16'h003B; B = 16'h00CA; #100;
A = 16'h003B; B = 16'h00CB; #100;
A = 16'h003B; B = 16'h00CC; #100;
A = 16'h003B; B = 16'h00CD; #100;
A = 16'h003B; B = 16'h00CE; #100;
A = 16'h003B; B = 16'h00CF; #100;
A = 16'h003B; B = 16'h00D0; #100;
A = 16'h003B; B = 16'h00D1; #100;
A = 16'h003B; B = 16'h00D2; #100;
A = 16'h003B; B = 16'h00D3; #100;
A = 16'h003B; B = 16'h00D4; #100;
A = 16'h003B; B = 16'h00D5; #100;
A = 16'h003B; B = 16'h00D6; #100;
A = 16'h003B; B = 16'h00D7; #100;
A = 16'h003B; B = 16'h00D8; #100;
A = 16'h003B; B = 16'h00D9; #100;
A = 16'h003B; B = 16'h00DA; #100;
A = 16'h003B; B = 16'h00DB; #100;
A = 16'h003B; B = 16'h00DC; #100;
A = 16'h003B; B = 16'h00DD; #100;
A = 16'h003B; B = 16'h00DE; #100;
A = 16'h003B; B = 16'h00DF; #100;
A = 16'h003B; B = 16'h00E0; #100;
A = 16'h003B; B = 16'h00E1; #100;
A = 16'h003B; B = 16'h00E2; #100;
A = 16'h003B; B = 16'h00E3; #100;
A = 16'h003B; B = 16'h00E4; #100;
A = 16'h003B; B = 16'h00E5; #100;
A = 16'h003B; B = 16'h00E6; #100;
A = 16'h003B; B = 16'h00E7; #100;
A = 16'h003B; B = 16'h00E8; #100;
A = 16'h003B; B = 16'h00E9; #100;
A = 16'h003B; B = 16'h00EA; #100;
A = 16'h003B; B = 16'h00EB; #100;
A = 16'h003B; B = 16'h00EC; #100;
A = 16'h003B; B = 16'h00ED; #100;
A = 16'h003B; B = 16'h00EE; #100;
A = 16'h003B; B = 16'h00EF; #100;
A = 16'h003B; B = 16'h00F0; #100;
A = 16'h003B; B = 16'h00F1; #100;
A = 16'h003B; B = 16'h00F2; #100;
A = 16'h003B; B = 16'h00F3; #100;
A = 16'h003B; B = 16'h00F4; #100;
A = 16'h003B; B = 16'h00F5; #100;
A = 16'h003B; B = 16'h00F6; #100;
A = 16'h003B; B = 16'h00F7; #100;
A = 16'h003B; B = 16'h00F8; #100;
A = 16'h003B; B = 16'h00F9; #100;
A = 16'h003B; B = 16'h00FA; #100;
A = 16'h003B; B = 16'h00FB; #100;
A = 16'h003B; B = 16'h00FC; #100;
A = 16'h003B; B = 16'h00FD; #100;
A = 16'h003B; B = 16'h00FE; #100;
A = 16'h003B; B = 16'h00FF; #100;
A = 16'h003C; B = 16'h000; #100;
A = 16'h003C; B = 16'h001; #100;
A = 16'h003C; B = 16'h002; #100;
A = 16'h003C; B = 16'h003; #100;
A = 16'h003C; B = 16'h004; #100;
A = 16'h003C; B = 16'h005; #100;
A = 16'h003C; B = 16'h006; #100;
A = 16'h003C; B = 16'h007; #100;
A = 16'h003C; B = 16'h008; #100;
A = 16'h003C; B = 16'h009; #100;
A = 16'h003C; B = 16'h00A; #100;
A = 16'h003C; B = 16'h00B; #100;
A = 16'h003C; B = 16'h00C; #100;
A = 16'h003C; B = 16'h00D; #100;
A = 16'h003C; B = 16'h00E; #100;
A = 16'h003C; B = 16'h00F; #100;
A = 16'h003C; B = 16'h0010; #100;
A = 16'h003C; B = 16'h0011; #100;
A = 16'h003C; B = 16'h0012; #100;
A = 16'h003C; B = 16'h0013; #100;
A = 16'h003C; B = 16'h0014; #100;
A = 16'h003C; B = 16'h0015; #100;
A = 16'h003C; B = 16'h0016; #100;
A = 16'h003C; B = 16'h0017; #100;
A = 16'h003C; B = 16'h0018; #100;
A = 16'h003C; B = 16'h0019; #100;
A = 16'h003C; B = 16'h001A; #100;
A = 16'h003C; B = 16'h001B; #100;
A = 16'h003C; B = 16'h001C; #100;
A = 16'h003C; B = 16'h001D; #100;
A = 16'h003C; B = 16'h001E; #100;
A = 16'h003C; B = 16'h001F; #100;
A = 16'h003C; B = 16'h0020; #100;
A = 16'h003C; B = 16'h0021; #100;
A = 16'h003C; B = 16'h0022; #100;
A = 16'h003C; B = 16'h0023; #100;
A = 16'h003C; B = 16'h0024; #100;
A = 16'h003C; B = 16'h0025; #100;
A = 16'h003C; B = 16'h0026; #100;
A = 16'h003C; B = 16'h0027; #100;
A = 16'h003C; B = 16'h0028; #100;
A = 16'h003C; B = 16'h0029; #100;
A = 16'h003C; B = 16'h002A; #100;
A = 16'h003C; B = 16'h002B; #100;
A = 16'h003C; B = 16'h002C; #100;
A = 16'h003C; B = 16'h002D; #100;
A = 16'h003C; B = 16'h002E; #100;
A = 16'h003C; B = 16'h002F; #100;
A = 16'h003C; B = 16'h0030; #100;
A = 16'h003C; B = 16'h0031; #100;
A = 16'h003C; B = 16'h0032; #100;
A = 16'h003C; B = 16'h0033; #100;
A = 16'h003C; B = 16'h0034; #100;
A = 16'h003C; B = 16'h0035; #100;
A = 16'h003C; B = 16'h0036; #100;
A = 16'h003C; B = 16'h0037; #100;
A = 16'h003C; B = 16'h0038; #100;
A = 16'h003C; B = 16'h0039; #100;
A = 16'h003C; B = 16'h003A; #100;
A = 16'h003C; B = 16'h003B; #100;
A = 16'h003C; B = 16'h003C; #100;
A = 16'h003C; B = 16'h003D; #100;
A = 16'h003C; B = 16'h003E; #100;
A = 16'h003C; B = 16'h003F; #100;
A = 16'h003C; B = 16'h0040; #100;
A = 16'h003C; B = 16'h0041; #100;
A = 16'h003C; B = 16'h0042; #100;
A = 16'h003C; B = 16'h0043; #100;
A = 16'h003C; B = 16'h0044; #100;
A = 16'h003C; B = 16'h0045; #100;
A = 16'h003C; B = 16'h0046; #100;
A = 16'h003C; B = 16'h0047; #100;
A = 16'h003C; B = 16'h0048; #100;
A = 16'h003C; B = 16'h0049; #100;
A = 16'h003C; B = 16'h004A; #100;
A = 16'h003C; B = 16'h004B; #100;
A = 16'h003C; B = 16'h004C; #100;
A = 16'h003C; B = 16'h004D; #100;
A = 16'h003C; B = 16'h004E; #100;
A = 16'h003C; B = 16'h004F; #100;
A = 16'h003C; B = 16'h0050; #100;
A = 16'h003C; B = 16'h0051; #100;
A = 16'h003C; B = 16'h0052; #100;
A = 16'h003C; B = 16'h0053; #100;
A = 16'h003C; B = 16'h0054; #100;
A = 16'h003C; B = 16'h0055; #100;
A = 16'h003C; B = 16'h0056; #100;
A = 16'h003C; B = 16'h0057; #100;
A = 16'h003C; B = 16'h0058; #100;
A = 16'h003C; B = 16'h0059; #100;
A = 16'h003C; B = 16'h005A; #100;
A = 16'h003C; B = 16'h005B; #100;
A = 16'h003C; B = 16'h005C; #100;
A = 16'h003C; B = 16'h005D; #100;
A = 16'h003C; B = 16'h005E; #100;
A = 16'h003C; B = 16'h005F; #100;
A = 16'h003C; B = 16'h0060; #100;
A = 16'h003C; B = 16'h0061; #100;
A = 16'h003C; B = 16'h0062; #100;
A = 16'h003C; B = 16'h0063; #100;
A = 16'h003C; B = 16'h0064; #100;
A = 16'h003C; B = 16'h0065; #100;
A = 16'h003C; B = 16'h0066; #100;
A = 16'h003C; B = 16'h0067; #100;
A = 16'h003C; B = 16'h0068; #100;
A = 16'h003C; B = 16'h0069; #100;
A = 16'h003C; B = 16'h006A; #100;
A = 16'h003C; B = 16'h006B; #100;
A = 16'h003C; B = 16'h006C; #100;
A = 16'h003C; B = 16'h006D; #100;
A = 16'h003C; B = 16'h006E; #100;
A = 16'h003C; B = 16'h006F; #100;
A = 16'h003C; B = 16'h0070; #100;
A = 16'h003C; B = 16'h0071; #100;
A = 16'h003C; B = 16'h0072; #100;
A = 16'h003C; B = 16'h0073; #100;
A = 16'h003C; B = 16'h0074; #100;
A = 16'h003C; B = 16'h0075; #100;
A = 16'h003C; B = 16'h0076; #100;
A = 16'h003C; B = 16'h0077; #100;
A = 16'h003C; B = 16'h0078; #100;
A = 16'h003C; B = 16'h0079; #100;
A = 16'h003C; B = 16'h007A; #100;
A = 16'h003C; B = 16'h007B; #100;
A = 16'h003C; B = 16'h007C; #100;
A = 16'h003C; B = 16'h007D; #100;
A = 16'h003C; B = 16'h007E; #100;
A = 16'h003C; B = 16'h007F; #100;
A = 16'h003C; B = 16'h0080; #100;
A = 16'h003C; B = 16'h0081; #100;
A = 16'h003C; B = 16'h0082; #100;
A = 16'h003C; B = 16'h0083; #100;
A = 16'h003C; B = 16'h0084; #100;
A = 16'h003C; B = 16'h0085; #100;
A = 16'h003C; B = 16'h0086; #100;
A = 16'h003C; B = 16'h0087; #100;
A = 16'h003C; B = 16'h0088; #100;
A = 16'h003C; B = 16'h0089; #100;
A = 16'h003C; B = 16'h008A; #100;
A = 16'h003C; B = 16'h008B; #100;
A = 16'h003C; B = 16'h008C; #100;
A = 16'h003C; B = 16'h008D; #100;
A = 16'h003C; B = 16'h008E; #100;
A = 16'h003C; B = 16'h008F; #100;
A = 16'h003C; B = 16'h0090; #100;
A = 16'h003C; B = 16'h0091; #100;
A = 16'h003C; B = 16'h0092; #100;
A = 16'h003C; B = 16'h0093; #100;
A = 16'h003C; B = 16'h0094; #100;
A = 16'h003C; B = 16'h0095; #100;
A = 16'h003C; B = 16'h0096; #100;
A = 16'h003C; B = 16'h0097; #100;
A = 16'h003C; B = 16'h0098; #100;
A = 16'h003C; B = 16'h0099; #100;
A = 16'h003C; B = 16'h009A; #100;
A = 16'h003C; B = 16'h009B; #100;
A = 16'h003C; B = 16'h009C; #100;
A = 16'h003C; B = 16'h009D; #100;
A = 16'h003C; B = 16'h009E; #100;
A = 16'h003C; B = 16'h009F; #100;
A = 16'h003C; B = 16'h00A0; #100;
A = 16'h003C; B = 16'h00A1; #100;
A = 16'h003C; B = 16'h00A2; #100;
A = 16'h003C; B = 16'h00A3; #100;
A = 16'h003C; B = 16'h00A4; #100;
A = 16'h003C; B = 16'h00A5; #100;
A = 16'h003C; B = 16'h00A6; #100;
A = 16'h003C; B = 16'h00A7; #100;
A = 16'h003C; B = 16'h00A8; #100;
A = 16'h003C; B = 16'h00A9; #100;
A = 16'h003C; B = 16'h00AA; #100;
A = 16'h003C; B = 16'h00AB; #100;
A = 16'h003C; B = 16'h00AC; #100;
A = 16'h003C; B = 16'h00AD; #100;
A = 16'h003C; B = 16'h00AE; #100;
A = 16'h003C; B = 16'h00AF; #100;
A = 16'h003C; B = 16'h00B0; #100;
A = 16'h003C; B = 16'h00B1; #100;
A = 16'h003C; B = 16'h00B2; #100;
A = 16'h003C; B = 16'h00B3; #100;
A = 16'h003C; B = 16'h00B4; #100;
A = 16'h003C; B = 16'h00B5; #100;
A = 16'h003C; B = 16'h00B6; #100;
A = 16'h003C; B = 16'h00B7; #100;
A = 16'h003C; B = 16'h00B8; #100;
A = 16'h003C; B = 16'h00B9; #100;
A = 16'h003C; B = 16'h00BA; #100;
A = 16'h003C; B = 16'h00BB; #100;
A = 16'h003C; B = 16'h00BC; #100;
A = 16'h003C; B = 16'h00BD; #100;
A = 16'h003C; B = 16'h00BE; #100;
A = 16'h003C; B = 16'h00BF; #100;
A = 16'h003C; B = 16'h00C0; #100;
A = 16'h003C; B = 16'h00C1; #100;
A = 16'h003C; B = 16'h00C2; #100;
A = 16'h003C; B = 16'h00C3; #100;
A = 16'h003C; B = 16'h00C4; #100;
A = 16'h003C; B = 16'h00C5; #100;
A = 16'h003C; B = 16'h00C6; #100;
A = 16'h003C; B = 16'h00C7; #100;
A = 16'h003C; B = 16'h00C8; #100;
A = 16'h003C; B = 16'h00C9; #100;
A = 16'h003C; B = 16'h00CA; #100;
A = 16'h003C; B = 16'h00CB; #100;
A = 16'h003C; B = 16'h00CC; #100;
A = 16'h003C; B = 16'h00CD; #100;
A = 16'h003C; B = 16'h00CE; #100;
A = 16'h003C; B = 16'h00CF; #100;
A = 16'h003C; B = 16'h00D0; #100;
A = 16'h003C; B = 16'h00D1; #100;
A = 16'h003C; B = 16'h00D2; #100;
A = 16'h003C; B = 16'h00D3; #100;
A = 16'h003C; B = 16'h00D4; #100;
A = 16'h003C; B = 16'h00D5; #100;
A = 16'h003C; B = 16'h00D6; #100;
A = 16'h003C; B = 16'h00D7; #100;
A = 16'h003C; B = 16'h00D8; #100;
A = 16'h003C; B = 16'h00D9; #100;
A = 16'h003C; B = 16'h00DA; #100;
A = 16'h003C; B = 16'h00DB; #100;
A = 16'h003C; B = 16'h00DC; #100;
A = 16'h003C; B = 16'h00DD; #100;
A = 16'h003C; B = 16'h00DE; #100;
A = 16'h003C; B = 16'h00DF; #100;
A = 16'h003C; B = 16'h00E0; #100;
A = 16'h003C; B = 16'h00E1; #100;
A = 16'h003C; B = 16'h00E2; #100;
A = 16'h003C; B = 16'h00E3; #100;
A = 16'h003C; B = 16'h00E4; #100;
A = 16'h003C; B = 16'h00E5; #100;
A = 16'h003C; B = 16'h00E6; #100;
A = 16'h003C; B = 16'h00E7; #100;
A = 16'h003C; B = 16'h00E8; #100;
A = 16'h003C; B = 16'h00E9; #100;
A = 16'h003C; B = 16'h00EA; #100;
A = 16'h003C; B = 16'h00EB; #100;
A = 16'h003C; B = 16'h00EC; #100;
A = 16'h003C; B = 16'h00ED; #100;
A = 16'h003C; B = 16'h00EE; #100;
A = 16'h003C; B = 16'h00EF; #100;
A = 16'h003C; B = 16'h00F0; #100;
A = 16'h003C; B = 16'h00F1; #100;
A = 16'h003C; B = 16'h00F2; #100;
A = 16'h003C; B = 16'h00F3; #100;
A = 16'h003C; B = 16'h00F4; #100;
A = 16'h003C; B = 16'h00F5; #100;
A = 16'h003C; B = 16'h00F6; #100;
A = 16'h003C; B = 16'h00F7; #100;
A = 16'h003C; B = 16'h00F8; #100;
A = 16'h003C; B = 16'h00F9; #100;
A = 16'h003C; B = 16'h00FA; #100;
A = 16'h003C; B = 16'h00FB; #100;
A = 16'h003C; B = 16'h00FC; #100;
A = 16'h003C; B = 16'h00FD; #100;
A = 16'h003C; B = 16'h00FE; #100;
A = 16'h003C; B = 16'h00FF; #100;
A = 16'h003D; B = 16'h000; #100;
A = 16'h003D; B = 16'h001; #100;
A = 16'h003D; B = 16'h002; #100;
A = 16'h003D; B = 16'h003; #100;
A = 16'h003D; B = 16'h004; #100;
A = 16'h003D; B = 16'h005; #100;
A = 16'h003D; B = 16'h006; #100;
A = 16'h003D; B = 16'h007; #100;
A = 16'h003D; B = 16'h008; #100;
A = 16'h003D; B = 16'h009; #100;
A = 16'h003D; B = 16'h00A; #100;
A = 16'h003D; B = 16'h00B; #100;
A = 16'h003D; B = 16'h00C; #100;
A = 16'h003D; B = 16'h00D; #100;
A = 16'h003D; B = 16'h00E; #100;
A = 16'h003D; B = 16'h00F; #100;
A = 16'h003D; B = 16'h0010; #100;
A = 16'h003D; B = 16'h0011; #100;
A = 16'h003D; B = 16'h0012; #100;
A = 16'h003D; B = 16'h0013; #100;
A = 16'h003D; B = 16'h0014; #100;
A = 16'h003D; B = 16'h0015; #100;
A = 16'h003D; B = 16'h0016; #100;
A = 16'h003D; B = 16'h0017; #100;
A = 16'h003D; B = 16'h0018; #100;
A = 16'h003D; B = 16'h0019; #100;
A = 16'h003D; B = 16'h001A; #100;
A = 16'h003D; B = 16'h001B; #100;
A = 16'h003D; B = 16'h001C; #100;
A = 16'h003D; B = 16'h001D; #100;
A = 16'h003D; B = 16'h001E; #100;
A = 16'h003D; B = 16'h001F; #100;
A = 16'h003D; B = 16'h0020; #100;
A = 16'h003D; B = 16'h0021; #100;
A = 16'h003D; B = 16'h0022; #100;
A = 16'h003D; B = 16'h0023; #100;
A = 16'h003D; B = 16'h0024; #100;
A = 16'h003D; B = 16'h0025; #100;
A = 16'h003D; B = 16'h0026; #100;
A = 16'h003D; B = 16'h0027; #100;
A = 16'h003D; B = 16'h0028; #100;
A = 16'h003D; B = 16'h0029; #100;
A = 16'h003D; B = 16'h002A; #100;
A = 16'h003D; B = 16'h002B; #100;
A = 16'h003D; B = 16'h002C; #100;
A = 16'h003D; B = 16'h002D; #100;
A = 16'h003D; B = 16'h002E; #100;
A = 16'h003D; B = 16'h002F; #100;
A = 16'h003D; B = 16'h0030; #100;
A = 16'h003D; B = 16'h0031; #100;
A = 16'h003D; B = 16'h0032; #100;
A = 16'h003D; B = 16'h0033; #100;
A = 16'h003D; B = 16'h0034; #100;
A = 16'h003D; B = 16'h0035; #100;
A = 16'h003D; B = 16'h0036; #100;
A = 16'h003D; B = 16'h0037; #100;
A = 16'h003D; B = 16'h0038; #100;
A = 16'h003D; B = 16'h0039; #100;
A = 16'h003D; B = 16'h003A; #100;
A = 16'h003D; B = 16'h003B; #100;
A = 16'h003D; B = 16'h003C; #100;
A = 16'h003D; B = 16'h003D; #100;
A = 16'h003D; B = 16'h003E; #100;
A = 16'h003D; B = 16'h003F; #100;
A = 16'h003D; B = 16'h0040; #100;
A = 16'h003D; B = 16'h0041; #100;
A = 16'h003D; B = 16'h0042; #100;
A = 16'h003D; B = 16'h0043; #100;
A = 16'h003D; B = 16'h0044; #100;
A = 16'h003D; B = 16'h0045; #100;
A = 16'h003D; B = 16'h0046; #100;
A = 16'h003D; B = 16'h0047; #100;
A = 16'h003D; B = 16'h0048; #100;
A = 16'h003D; B = 16'h0049; #100;
A = 16'h003D; B = 16'h004A; #100;
A = 16'h003D; B = 16'h004B; #100;
A = 16'h003D; B = 16'h004C; #100;
A = 16'h003D; B = 16'h004D; #100;
A = 16'h003D; B = 16'h004E; #100;
A = 16'h003D; B = 16'h004F; #100;
A = 16'h003D; B = 16'h0050; #100;
A = 16'h003D; B = 16'h0051; #100;
A = 16'h003D; B = 16'h0052; #100;
A = 16'h003D; B = 16'h0053; #100;
A = 16'h003D; B = 16'h0054; #100;
A = 16'h003D; B = 16'h0055; #100;
A = 16'h003D; B = 16'h0056; #100;
A = 16'h003D; B = 16'h0057; #100;
A = 16'h003D; B = 16'h0058; #100;
A = 16'h003D; B = 16'h0059; #100;
A = 16'h003D; B = 16'h005A; #100;
A = 16'h003D; B = 16'h005B; #100;
A = 16'h003D; B = 16'h005C; #100;
A = 16'h003D; B = 16'h005D; #100;
A = 16'h003D; B = 16'h005E; #100;
A = 16'h003D; B = 16'h005F; #100;
A = 16'h003D; B = 16'h0060; #100;
A = 16'h003D; B = 16'h0061; #100;
A = 16'h003D; B = 16'h0062; #100;
A = 16'h003D; B = 16'h0063; #100;
A = 16'h003D; B = 16'h0064; #100;
A = 16'h003D; B = 16'h0065; #100;
A = 16'h003D; B = 16'h0066; #100;
A = 16'h003D; B = 16'h0067; #100;
A = 16'h003D; B = 16'h0068; #100;
A = 16'h003D; B = 16'h0069; #100;
A = 16'h003D; B = 16'h006A; #100;
A = 16'h003D; B = 16'h006B; #100;
A = 16'h003D; B = 16'h006C; #100;
A = 16'h003D; B = 16'h006D; #100;
A = 16'h003D; B = 16'h006E; #100;
A = 16'h003D; B = 16'h006F; #100;
A = 16'h003D; B = 16'h0070; #100;
A = 16'h003D; B = 16'h0071; #100;
A = 16'h003D; B = 16'h0072; #100;
A = 16'h003D; B = 16'h0073; #100;
A = 16'h003D; B = 16'h0074; #100;
A = 16'h003D; B = 16'h0075; #100;
A = 16'h003D; B = 16'h0076; #100;
A = 16'h003D; B = 16'h0077; #100;
A = 16'h003D; B = 16'h0078; #100;
A = 16'h003D; B = 16'h0079; #100;
A = 16'h003D; B = 16'h007A; #100;
A = 16'h003D; B = 16'h007B; #100;
A = 16'h003D; B = 16'h007C; #100;
A = 16'h003D; B = 16'h007D; #100;
A = 16'h003D; B = 16'h007E; #100;
A = 16'h003D; B = 16'h007F; #100;
A = 16'h003D; B = 16'h0080; #100;
A = 16'h003D; B = 16'h0081; #100;
A = 16'h003D; B = 16'h0082; #100;
A = 16'h003D; B = 16'h0083; #100;
A = 16'h003D; B = 16'h0084; #100;
A = 16'h003D; B = 16'h0085; #100;
A = 16'h003D; B = 16'h0086; #100;
A = 16'h003D; B = 16'h0087; #100;
A = 16'h003D; B = 16'h0088; #100;
A = 16'h003D; B = 16'h0089; #100;
A = 16'h003D; B = 16'h008A; #100;
A = 16'h003D; B = 16'h008B; #100;
A = 16'h003D; B = 16'h008C; #100;
A = 16'h003D; B = 16'h008D; #100;
A = 16'h003D; B = 16'h008E; #100;
A = 16'h003D; B = 16'h008F; #100;
A = 16'h003D; B = 16'h0090; #100;
A = 16'h003D; B = 16'h0091; #100;
A = 16'h003D; B = 16'h0092; #100;
A = 16'h003D; B = 16'h0093; #100;
A = 16'h003D; B = 16'h0094; #100;
A = 16'h003D; B = 16'h0095; #100;
A = 16'h003D; B = 16'h0096; #100;
A = 16'h003D; B = 16'h0097; #100;
A = 16'h003D; B = 16'h0098; #100;
A = 16'h003D; B = 16'h0099; #100;
A = 16'h003D; B = 16'h009A; #100;
A = 16'h003D; B = 16'h009B; #100;
A = 16'h003D; B = 16'h009C; #100;
A = 16'h003D; B = 16'h009D; #100;
A = 16'h003D; B = 16'h009E; #100;
A = 16'h003D; B = 16'h009F; #100;
A = 16'h003D; B = 16'h00A0; #100;
A = 16'h003D; B = 16'h00A1; #100;
A = 16'h003D; B = 16'h00A2; #100;
A = 16'h003D; B = 16'h00A3; #100;
A = 16'h003D; B = 16'h00A4; #100;
A = 16'h003D; B = 16'h00A5; #100;
A = 16'h003D; B = 16'h00A6; #100;
A = 16'h003D; B = 16'h00A7; #100;
A = 16'h003D; B = 16'h00A8; #100;
A = 16'h003D; B = 16'h00A9; #100;
A = 16'h003D; B = 16'h00AA; #100;
A = 16'h003D; B = 16'h00AB; #100;
A = 16'h003D; B = 16'h00AC; #100;
A = 16'h003D; B = 16'h00AD; #100;
A = 16'h003D; B = 16'h00AE; #100;
A = 16'h003D; B = 16'h00AF; #100;
A = 16'h003D; B = 16'h00B0; #100;
A = 16'h003D; B = 16'h00B1; #100;
A = 16'h003D; B = 16'h00B2; #100;
A = 16'h003D; B = 16'h00B3; #100;
A = 16'h003D; B = 16'h00B4; #100;
A = 16'h003D; B = 16'h00B5; #100;
A = 16'h003D; B = 16'h00B6; #100;
A = 16'h003D; B = 16'h00B7; #100;
A = 16'h003D; B = 16'h00B8; #100;
A = 16'h003D; B = 16'h00B9; #100;
A = 16'h003D; B = 16'h00BA; #100;
A = 16'h003D; B = 16'h00BB; #100;
A = 16'h003D; B = 16'h00BC; #100;
A = 16'h003D; B = 16'h00BD; #100;
A = 16'h003D; B = 16'h00BE; #100;
A = 16'h003D; B = 16'h00BF; #100;
A = 16'h003D; B = 16'h00C0; #100;
A = 16'h003D; B = 16'h00C1; #100;
A = 16'h003D; B = 16'h00C2; #100;
A = 16'h003D; B = 16'h00C3; #100;
A = 16'h003D; B = 16'h00C4; #100;
A = 16'h003D; B = 16'h00C5; #100;
A = 16'h003D; B = 16'h00C6; #100;
A = 16'h003D; B = 16'h00C7; #100;
A = 16'h003D; B = 16'h00C8; #100;
A = 16'h003D; B = 16'h00C9; #100;
A = 16'h003D; B = 16'h00CA; #100;
A = 16'h003D; B = 16'h00CB; #100;
A = 16'h003D; B = 16'h00CC; #100;
A = 16'h003D; B = 16'h00CD; #100;
A = 16'h003D; B = 16'h00CE; #100;
A = 16'h003D; B = 16'h00CF; #100;
A = 16'h003D; B = 16'h00D0; #100;
A = 16'h003D; B = 16'h00D1; #100;
A = 16'h003D; B = 16'h00D2; #100;
A = 16'h003D; B = 16'h00D3; #100;
A = 16'h003D; B = 16'h00D4; #100;
A = 16'h003D; B = 16'h00D5; #100;
A = 16'h003D; B = 16'h00D6; #100;
A = 16'h003D; B = 16'h00D7; #100;
A = 16'h003D; B = 16'h00D8; #100;
A = 16'h003D; B = 16'h00D9; #100;
A = 16'h003D; B = 16'h00DA; #100;
A = 16'h003D; B = 16'h00DB; #100;
A = 16'h003D; B = 16'h00DC; #100;
A = 16'h003D; B = 16'h00DD; #100;
A = 16'h003D; B = 16'h00DE; #100;
A = 16'h003D; B = 16'h00DF; #100;
A = 16'h003D; B = 16'h00E0; #100;
A = 16'h003D; B = 16'h00E1; #100;
A = 16'h003D; B = 16'h00E2; #100;
A = 16'h003D; B = 16'h00E3; #100;
A = 16'h003D; B = 16'h00E4; #100;
A = 16'h003D; B = 16'h00E5; #100;
A = 16'h003D; B = 16'h00E6; #100;
A = 16'h003D; B = 16'h00E7; #100;
A = 16'h003D; B = 16'h00E8; #100;
A = 16'h003D; B = 16'h00E9; #100;
A = 16'h003D; B = 16'h00EA; #100;
A = 16'h003D; B = 16'h00EB; #100;
A = 16'h003D; B = 16'h00EC; #100;
A = 16'h003D; B = 16'h00ED; #100;
A = 16'h003D; B = 16'h00EE; #100;
A = 16'h003D; B = 16'h00EF; #100;
A = 16'h003D; B = 16'h00F0; #100;
A = 16'h003D; B = 16'h00F1; #100;
A = 16'h003D; B = 16'h00F2; #100;
A = 16'h003D; B = 16'h00F3; #100;
A = 16'h003D; B = 16'h00F4; #100;
A = 16'h003D; B = 16'h00F5; #100;
A = 16'h003D; B = 16'h00F6; #100;
A = 16'h003D; B = 16'h00F7; #100;
A = 16'h003D; B = 16'h00F8; #100;
A = 16'h003D; B = 16'h00F9; #100;
A = 16'h003D; B = 16'h00FA; #100;
A = 16'h003D; B = 16'h00FB; #100;
A = 16'h003D; B = 16'h00FC; #100;
A = 16'h003D; B = 16'h00FD; #100;
A = 16'h003D; B = 16'h00FE; #100;
A = 16'h003D; B = 16'h00FF; #100;
A = 16'h003E; B = 16'h000; #100;
A = 16'h003E; B = 16'h001; #100;
A = 16'h003E; B = 16'h002; #100;
A = 16'h003E; B = 16'h003; #100;
A = 16'h003E; B = 16'h004; #100;
A = 16'h003E; B = 16'h005; #100;
A = 16'h003E; B = 16'h006; #100;
A = 16'h003E; B = 16'h007; #100;
A = 16'h003E; B = 16'h008; #100;
A = 16'h003E; B = 16'h009; #100;
A = 16'h003E; B = 16'h00A; #100;
A = 16'h003E; B = 16'h00B; #100;
A = 16'h003E; B = 16'h00C; #100;
A = 16'h003E; B = 16'h00D; #100;
A = 16'h003E; B = 16'h00E; #100;
A = 16'h003E; B = 16'h00F; #100;
A = 16'h003E; B = 16'h0010; #100;
A = 16'h003E; B = 16'h0011; #100;
A = 16'h003E; B = 16'h0012; #100;
A = 16'h003E; B = 16'h0013; #100;
A = 16'h003E; B = 16'h0014; #100;
A = 16'h003E; B = 16'h0015; #100;
A = 16'h003E; B = 16'h0016; #100;
A = 16'h003E; B = 16'h0017; #100;
A = 16'h003E; B = 16'h0018; #100;
A = 16'h003E; B = 16'h0019; #100;
A = 16'h003E; B = 16'h001A; #100;
A = 16'h003E; B = 16'h001B; #100;
A = 16'h003E; B = 16'h001C; #100;
A = 16'h003E; B = 16'h001D; #100;
A = 16'h003E; B = 16'h001E; #100;
A = 16'h003E; B = 16'h001F; #100;
A = 16'h003E; B = 16'h0020; #100;
A = 16'h003E; B = 16'h0021; #100;
A = 16'h003E; B = 16'h0022; #100;
A = 16'h003E; B = 16'h0023; #100;
A = 16'h003E; B = 16'h0024; #100;
A = 16'h003E; B = 16'h0025; #100;
A = 16'h003E; B = 16'h0026; #100;
A = 16'h003E; B = 16'h0027; #100;
A = 16'h003E; B = 16'h0028; #100;
A = 16'h003E; B = 16'h0029; #100;
A = 16'h003E; B = 16'h002A; #100;
A = 16'h003E; B = 16'h002B; #100;
A = 16'h003E; B = 16'h002C; #100;
A = 16'h003E; B = 16'h002D; #100;
A = 16'h003E; B = 16'h002E; #100;
A = 16'h003E; B = 16'h002F; #100;
A = 16'h003E; B = 16'h0030; #100;
A = 16'h003E; B = 16'h0031; #100;
A = 16'h003E; B = 16'h0032; #100;
A = 16'h003E; B = 16'h0033; #100;
A = 16'h003E; B = 16'h0034; #100;
A = 16'h003E; B = 16'h0035; #100;
A = 16'h003E; B = 16'h0036; #100;
A = 16'h003E; B = 16'h0037; #100;
A = 16'h003E; B = 16'h0038; #100;
A = 16'h003E; B = 16'h0039; #100;
A = 16'h003E; B = 16'h003A; #100;
A = 16'h003E; B = 16'h003B; #100;
A = 16'h003E; B = 16'h003C; #100;
A = 16'h003E; B = 16'h003D; #100;
A = 16'h003E; B = 16'h003E; #100;
A = 16'h003E; B = 16'h003F; #100;
A = 16'h003E; B = 16'h0040; #100;
A = 16'h003E; B = 16'h0041; #100;
A = 16'h003E; B = 16'h0042; #100;
A = 16'h003E; B = 16'h0043; #100;
A = 16'h003E; B = 16'h0044; #100;
A = 16'h003E; B = 16'h0045; #100;
A = 16'h003E; B = 16'h0046; #100;
A = 16'h003E; B = 16'h0047; #100;
A = 16'h003E; B = 16'h0048; #100;
A = 16'h003E; B = 16'h0049; #100;
A = 16'h003E; B = 16'h004A; #100;
A = 16'h003E; B = 16'h004B; #100;
A = 16'h003E; B = 16'h004C; #100;
A = 16'h003E; B = 16'h004D; #100;
A = 16'h003E; B = 16'h004E; #100;
A = 16'h003E; B = 16'h004F; #100;
A = 16'h003E; B = 16'h0050; #100;
A = 16'h003E; B = 16'h0051; #100;
A = 16'h003E; B = 16'h0052; #100;
A = 16'h003E; B = 16'h0053; #100;
A = 16'h003E; B = 16'h0054; #100;
A = 16'h003E; B = 16'h0055; #100;
A = 16'h003E; B = 16'h0056; #100;
A = 16'h003E; B = 16'h0057; #100;
A = 16'h003E; B = 16'h0058; #100;
A = 16'h003E; B = 16'h0059; #100;
A = 16'h003E; B = 16'h005A; #100;
A = 16'h003E; B = 16'h005B; #100;
A = 16'h003E; B = 16'h005C; #100;
A = 16'h003E; B = 16'h005D; #100;
A = 16'h003E; B = 16'h005E; #100;
A = 16'h003E; B = 16'h005F; #100;
A = 16'h003E; B = 16'h0060; #100;
A = 16'h003E; B = 16'h0061; #100;
A = 16'h003E; B = 16'h0062; #100;
A = 16'h003E; B = 16'h0063; #100;
A = 16'h003E; B = 16'h0064; #100;
A = 16'h003E; B = 16'h0065; #100;
A = 16'h003E; B = 16'h0066; #100;
A = 16'h003E; B = 16'h0067; #100;
A = 16'h003E; B = 16'h0068; #100;
A = 16'h003E; B = 16'h0069; #100;
A = 16'h003E; B = 16'h006A; #100;
A = 16'h003E; B = 16'h006B; #100;
A = 16'h003E; B = 16'h006C; #100;
A = 16'h003E; B = 16'h006D; #100;
A = 16'h003E; B = 16'h006E; #100;
A = 16'h003E; B = 16'h006F; #100;
A = 16'h003E; B = 16'h0070; #100;
A = 16'h003E; B = 16'h0071; #100;
A = 16'h003E; B = 16'h0072; #100;
A = 16'h003E; B = 16'h0073; #100;
A = 16'h003E; B = 16'h0074; #100;
A = 16'h003E; B = 16'h0075; #100;
A = 16'h003E; B = 16'h0076; #100;
A = 16'h003E; B = 16'h0077; #100;
A = 16'h003E; B = 16'h0078; #100;
A = 16'h003E; B = 16'h0079; #100;
A = 16'h003E; B = 16'h007A; #100;
A = 16'h003E; B = 16'h007B; #100;
A = 16'h003E; B = 16'h007C; #100;
A = 16'h003E; B = 16'h007D; #100;
A = 16'h003E; B = 16'h007E; #100;
A = 16'h003E; B = 16'h007F; #100;
A = 16'h003E; B = 16'h0080; #100;
A = 16'h003E; B = 16'h0081; #100;
A = 16'h003E; B = 16'h0082; #100;
A = 16'h003E; B = 16'h0083; #100;
A = 16'h003E; B = 16'h0084; #100;
A = 16'h003E; B = 16'h0085; #100;
A = 16'h003E; B = 16'h0086; #100;
A = 16'h003E; B = 16'h0087; #100;
A = 16'h003E; B = 16'h0088; #100;
A = 16'h003E; B = 16'h0089; #100;
A = 16'h003E; B = 16'h008A; #100;
A = 16'h003E; B = 16'h008B; #100;
A = 16'h003E; B = 16'h008C; #100;
A = 16'h003E; B = 16'h008D; #100;
A = 16'h003E; B = 16'h008E; #100;
A = 16'h003E; B = 16'h008F; #100;
A = 16'h003E; B = 16'h0090; #100;
A = 16'h003E; B = 16'h0091; #100;
A = 16'h003E; B = 16'h0092; #100;
A = 16'h003E; B = 16'h0093; #100;
A = 16'h003E; B = 16'h0094; #100;
A = 16'h003E; B = 16'h0095; #100;
A = 16'h003E; B = 16'h0096; #100;
A = 16'h003E; B = 16'h0097; #100;
A = 16'h003E; B = 16'h0098; #100;
A = 16'h003E; B = 16'h0099; #100;
A = 16'h003E; B = 16'h009A; #100;
A = 16'h003E; B = 16'h009B; #100;
A = 16'h003E; B = 16'h009C; #100;
A = 16'h003E; B = 16'h009D; #100;
A = 16'h003E; B = 16'h009E; #100;
A = 16'h003E; B = 16'h009F; #100;
A = 16'h003E; B = 16'h00A0; #100;
A = 16'h003E; B = 16'h00A1; #100;
A = 16'h003E; B = 16'h00A2; #100;
A = 16'h003E; B = 16'h00A3; #100;
A = 16'h003E; B = 16'h00A4; #100;
A = 16'h003E; B = 16'h00A5; #100;
A = 16'h003E; B = 16'h00A6; #100;
A = 16'h003E; B = 16'h00A7; #100;
A = 16'h003E; B = 16'h00A8; #100;
A = 16'h003E; B = 16'h00A9; #100;
A = 16'h003E; B = 16'h00AA; #100;
A = 16'h003E; B = 16'h00AB; #100;
A = 16'h003E; B = 16'h00AC; #100;
A = 16'h003E; B = 16'h00AD; #100;
A = 16'h003E; B = 16'h00AE; #100;
A = 16'h003E; B = 16'h00AF; #100;
A = 16'h003E; B = 16'h00B0; #100;
A = 16'h003E; B = 16'h00B1; #100;
A = 16'h003E; B = 16'h00B2; #100;
A = 16'h003E; B = 16'h00B3; #100;
A = 16'h003E; B = 16'h00B4; #100;
A = 16'h003E; B = 16'h00B5; #100;
A = 16'h003E; B = 16'h00B6; #100;
A = 16'h003E; B = 16'h00B7; #100;
A = 16'h003E; B = 16'h00B8; #100;
A = 16'h003E; B = 16'h00B9; #100;
A = 16'h003E; B = 16'h00BA; #100;
A = 16'h003E; B = 16'h00BB; #100;
A = 16'h003E; B = 16'h00BC; #100;
A = 16'h003E; B = 16'h00BD; #100;
A = 16'h003E; B = 16'h00BE; #100;
A = 16'h003E; B = 16'h00BF; #100;
A = 16'h003E; B = 16'h00C0; #100;
A = 16'h003E; B = 16'h00C1; #100;
A = 16'h003E; B = 16'h00C2; #100;
A = 16'h003E; B = 16'h00C3; #100;
A = 16'h003E; B = 16'h00C4; #100;
A = 16'h003E; B = 16'h00C5; #100;
A = 16'h003E; B = 16'h00C6; #100;
A = 16'h003E; B = 16'h00C7; #100;
A = 16'h003E; B = 16'h00C8; #100;
A = 16'h003E; B = 16'h00C9; #100;
A = 16'h003E; B = 16'h00CA; #100;
A = 16'h003E; B = 16'h00CB; #100;
A = 16'h003E; B = 16'h00CC; #100;
A = 16'h003E; B = 16'h00CD; #100;
A = 16'h003E; B = 16'h00CE; #100;
A = 16'h003E; B = 16'h00CF; #100;
A = 16'h003E; B = 16'h00D0; #100;
A = 16'h003E; B = 16'h00D1; #100;
A = 16'h003E; B = 16'h00D2; #100;
A = 16'h003E; B = 16'h00D3; #100;
A = 16'h003E; B = 16'h00D4; #100;
A = 16'h003E; B = 16'h00D5; #100;
A = 16'h003E; B = 16'h00D6; #100;
A = 16'h003E; B = 16'h00D7; #100;
A = 16'h003E; B = 16'h00D8; #100;
A = 16'h003E; B = 16'h00D9; #100;
A = 16'h003E; B = 16'h00DA; #100;
A = 16'h003E; B = 16'h00DB; #100;
A = 16'h003E; B = 16'h00DC; #100;
A = 16'h003E; B = 16'h00DD; #100;
A = 16'h003E; B = 16'h00DE; #100;
A = 16'h003E; B = 16'h00DF; #100;
A = 16'h003E; B = 16'h00E0; #100;
A = 16'h003E; B = 16'h00E1; #100;
A = 16'h003E; B = 16'h00E2; #100;
A = 16'h003E; B = 16'h00E3; #100;
A = 16'h003E; B = 16'h00E4; #100;
A = 16'h003E; B = 16'h00E5; #100;
A = 16'h003E; B = 16'h00E6; #100;
A = 16'h003E; B = 16'h00E7; #100;
A = 16'h003E; B = 16'h00E8; #100;
A = 16'h003E; B = 16'h00E9; #100;
A = 16'h003E; B = 16'h00EA; #100;
A = 16'h003E; B = 16'h00EB; #100;
A = 16'h003E; B = 16'h00EC; #100;
A = 16'h003E; B = 16'h00ED; #100;
A = 16'h003E; B = 16'h00EE; #100;
A = 16'h003E; B = 16'h00EF; #100;
A = 16'h003E; B = 16'h00F0; #100;
A = 16'h003E; B = 16'h00F1; #100;
A = 16'h003E; B = 16'h00F2; #100;
A = 16'h003E; B = 16'h00F3; #100;
A = 16'h003E; B = 16'h00F4; #100;
A = 16'h003E; B = 16'h00F5; #100;
A = 16'h003E; B = 16'h00F6; #100;
A = 16'h003E; B = 16'h00F7; #100;
A = 16'h003E; B = 16'h00F8; #100;
A = 16'h003E; B = 16'h00F9; #100;
A = 16'h003E; B = 16'h00FA; #100;
A = 16'h003E; B = 16'h00FB; #100;
A = 16'h003E; B = 16'h00FC; #100;
A = 16'h003E; B = 16'h00FD; #100;
A = 16'h003E; B = 16'h00FE; #100;
A = 16'h003E; B = 16'h00FF; #100;
A = 16'h003F; B = 16'h000; #100;
A = 16'h003F; B = 16'h001; #100;
A = 16'h003F; B = 16'h002; #100;
A = 16'h003F; B = 16'h003; #100;
A = 16'h003F; B = 16'h004; #100;
A = 16'h003F; B = 16'h005; #100;
A = 16'h003F; B = 16'h006; #100;
A = 16'h003F; B = 16'h007; #100;
A = 16'h003F; B = 16'h008; #100;
A = 16'h003F; B = 16'h009; #100;
A = 16'h003F; B = 16'h00A; #100;
A = 16'h003F; B = 16'h00B; #100;
A = 16'h003F; B = 16'h00C; #100;
A = 16'h003F; B = 16'h00D; #100;
A = 16'h003F; B = 16'h00E; #100;
A = 16'h003F; B = 16'h00F; #100;
A = 16'h003F; B = 16'h0010; #100;
A = 16'h003F; B = 16'h0011; #100;
A = 16'h003F; B = 16'h0012; #100;
A = 16'h003F; B = 16'h0013; #100;
A = 16'h003F; B = 16'h0014; #100;
A = 16'h003F; B = 16'h0015; #100;
A = 16'h003F; B = 16'h0016; #100;
A = 16'h003F; B = 16'h0017; #100;
A = 16'h003F; B = 16'h0018; #100;
A = 16'h003F; B = 16'h0019; #100;
A = 16'h003F; B = 16'h001A; #100;
A = 16'h003F; B = 16'h001B; #100;
A = 16'h003F; B = 16'h001C; #100;
A = 16'h003F; B = 16'h001D; #100;
A = 16'h003F; B = 16'h001E; #100;
A = 16'h003F; B = 16'h001F; #100;
A = 16'h003F; B = 16'h0020; #100;
A = 16'h003F; B = 16'h0021; #100;
A = 16'h003F; B = 16'h0022; #100;
A = 16'h003F; B = 16'h0023; #100;
A = 16'h003F; B = 16'h0024; #100;
A = 16'h003F; B = 16'h0025; #100;
A = 16'h003F; B = 16'h0026; #100;
A = 16'h003F; B = 16'h0027; #100;
A = 16'h003F; B = 16'h0028; #100;
A = 16'h003F; B = 16'h0029; #100;
A = 16'h003F; B = 16'h002A; #100;
A = 16'h003F; B = 16'h002B; #100;
A = 16'h003F; B = 16'h002C; #100;
A = 16'h003F; B = 16'h002D; #100;
A = 16'h003F; B = 16'h002E; #100;
A = 16'h003F; B = 16'h002F; #100;
A = 16'h003F; B = 16'h0030; #100;
A = 16'h003F; B = 16'h0031; #100;
A = 16'h003F; B = 16'h0032; #100;
A = 16'h003F; B = 16'h0033; #100;
A = 16'h003F; B = 16'h0034; #100;
A = 16'h003F; B = 16'h0035; #100;
A = 16'h003F; B = 16'h0036; #100;
A = 16'h003F; B = 16'h0037; #100;
A = 16'h003F; B = 16'h0038; #100;
A = 16'h003F; B = 16'h0039; #100;
A = 16'h003F; B = 16'h003A; #100;
A = 16'h003F; B = 16'h003B; #100;
A = 16'h003F; B = 16'h003C; #100;
A = 16'h003F; B = 16'h003D; #100;
A = 16'h003F; B = 16'h003E; #100;
A = 16'h003F; B = 16'h003F; #100;
A = 16'h003F; B = 16'h0040; #100;
A = 16'h003F; B = 16'h0041; #100;
A = 16'h003F; B = 16'h0042; #100;
A = 16'h003F; B = 16'h0043; #100;
A = 16'h003F; B = 16'h0044; #100;
A = 16'h003F; B = 16'h0045; #100;
A = 16'h003F; B = 16'h0046; #100;
A = 16'h003F; B = 16'h0047; #100;
A = 16'h003F; B = 16'h0048; #100;
A = 16'h003F; B = 16'h0049; #100;
A = 16'h003F; B = 16'h004A; #100;
A = 16'h003F; B = 16'h004B; #100;
A = 16'h003F; B = 16'h004C; #100;
A = 16'h003F; B = 16'h004D; #100;
A = 16'h003F; B = 16'h004E; #100;
A = 16'h003F; B = 16'h004F; #100;
A = 16'h003F; B = 16'h0050; #100;
A = 16'h003F; B = 16'h0051; #100;
A = 16'h003F; B = 16'h0052; #100;
A = 16'h003F; B = 16'h0053; #100;
A = 16'h003F; B = 16'h0054; #100;
A = 16'h003F; B = 16'h0055; #100;
A = 16'h003F; B = 16'h0056; #100;
A = 16'h003F; B = 16'h0057; #100;
A = 16'h003F; B = 16'h0058; #100;
A = 16'h003F; B = 16'h0059; #100;
A = 16'h003F; B = 16'h005A; #100;
A = 16'h003F; B = 16'h005B; #100;
A = 16'h003F; B = 16'h005C; #100;
A = 16'h003F; B = 16'h005D; #100;
A = 16'h003F; B = 16'h005E; #100;
A = 16'h003F; B = 16'h005F; #100;
A = 16'h003F; B = 16'h0060; #100;
A = 16'h003F; B = 16'h0061; #100;
A = 16'h003F; B = 16'h0062; #100;
A = 16'h003F; B = 16'h0063; #100;
A = 16'h003F; B = 16'h0064; #100;
A = 16'h003F; B = 16'h0065; #100;
A = 16'h003F; B = 16'h0066; #100;
A = 16'h003F; B = 16'h0067; #100;
A = 16'h003F; B = 16'h0068; #100;
A = 16'h003F; B = 16'h0069; #100;
A = 16'h003F; B = 16'h006A; #100;
A = 16'h003F; B = 16'h006B; #100;
A = 16'h003F; B = 16'h006C; #100;
A = 16'h003F; B = 16'h006D; #100;
A = 16'h003F; B = 16'h006E; #100;
A = 16'h003F; B = 16'h006F; #100;
A = 16'h003F; B = 16'h0070; #100;
A = 16'h003F; B = 16'h0071; #100;
A = 16'h003F; B = 16'h0072; #100;
A = 16'h003F; B = 16'h0073; #100;
A = 16'h003F; B = 16'h0074; #100;
A = 16'h003F; B = 16'h0075; #100;
A = 16'h003F; B = 16'h0076; #100;
A = 16'h003F; B = 16'h0077; #100;
A = 16'h003F; B = 16'h0078; #100;
A = 16'h003F; B = 16'h0079; #100;
A = 16'h003F; B = 16'h007A; #100;
A = 16'h003F; B = 16'h007B; #100;
A = 16'h003F; B = 16'h007C; #100;
A = 16'h003F; B = 16'h007D; #100;
A = 16'h003F; B = 16'h007E; #100;
A = 16'h003F; B = 16'h007F; #100;
A = 16'h003F; B = 16'h0080; #100;
A = 16'h003F; B = 16'h0081; #100;
A = 16'h003F; B = 16'h0082; #100;
A = 16'h003F; B = 16'h0083; #100;
A = 16'h003F; B = 16'h0084; #100;
A = 16'h003F; B = 16'h0085; #100;
A = 16'h003F; B = 16'h0086; #100;
A = 16'h003F; B = 16'h0087; #100;
A = 16'h003F; B = 16'h0088; #100;
A = 16'h003F; B = 16'h0089; #100;
A = 16'h003F; B = 16'h008A; #100;
A = 16'h003F; B = 16'h008B; #100;
A = 16'h003F; B = 16'h008C; #100;
A = 16'h003F; B = 16'h008D; #100;
A = 16'h003F; B = 16'h008E; #100;
A = 16'h003F; B = 16'h008F; #100;
A = 16'h003F; B = 16'h0090; #100;
A = 16'h003F; B = 16'h0091; #100;
A = 16'h003F; B = 16'h0092; #100;
A = 16'h003F; B = 16'h0093; #100;
A = 16'h003F; B = 16'h0094; #100;
A = 16'h003F; B = 16'h0095; #100;
A = 16'h003F; B = 16'h0096; #100;
A = 16'h003F; B = 16'h0097; #100;
A = 16'h003F; B = 16'h0098; #100;
A = 16'h003F; B = 16'h0099; #100;
A = 16'h003F; B = 16'h009A; #100;
A = 16'h003F; B = 16'h009B; #100;
A = 16'h003F; B = 16'h009C; #100;
A = 16'h003F; B = 16'h009D; #100;
A = 16'h003F; B = 16'h009E; #100;
A = 16'h003F; B = 16'h009F; #100;
A = 16'h003F; B = 16'h00A0; #100;
A = 16'h003F; B = 16'h00A1; #100;
A = 16'h003F; B = 16'h00A2; #100;
A = 16'h003F; B = 16'h00A3; #100;
A = 16'h003F; B = 16'h00A4; #100;
A = 16'h003F; B = 16'h00A5; #100;
A = 16'h003F; B = 16'h00A6; #100;
A = 16'h003F; B = 16'h00A7; #100;
A = 16'h003F; B = 16'h00A8; #100;
A = 16'h003F; B = 16'h00A9; #100;
A = 16'h003F; B = 16'h00AA; #100;
A = 16'h003F; B = 16'h00AB; #100;
A = 16'h003F; B = 16'h00AC; #100;
A = 16'h003F; B = 16'h00AD; #100;
A = 16'h003F; B = 16'h00AE; #100;
A = 16'h003F; B = 16'h00AF; #100;
A = 16'h003F; B = 16'h00B0; #100;
A = 16'h003F; B = 16'h00B1; #100;
A = 16'h003F; B = 16'h00B2; #100;
A = 16'h003F; B = 16'h00B3; #100;
A = 16'h003F; B = 16'h00B4; #100;
A = 16'h003F; B = 16'h00B5; #100;
A = 16'h003F; B = 16'h00B6; #100;
A = 16'h003F; B = 16'h00B7; #100;
A = 16'h003F; B = 16'h00B8; #100;
A = 16'h003F; B = 16'h00B9; #100;
A = 16'h003F; B = 16'h00BA; #100;
A = 16'h003F; B = 16'h00BB; #100;
A = 16'h003F; B = 16'h00BC; #100;
A = 16'h003F; B = 16'h00BD; #100;
A = 16'h003F; B = 16'h00BE; #100;
A = 16'h003F; B = 16'h00BF; #100;
A = 16'h003F; B = 16'h00C0; #100;
A = 16'h003F; B = 16'h00C1; #100;
A = 16'h003F; B = 16'h00C2; #100;
A = 16'h003F; B = 16'h00C3; #100;
A = 16'h003F; B = 16'h00C4; #100;
A = 16'h003F; B = 16'h00C5; #100;
A = 16'h003F; B = 16'h00C6; #100;
A = 16'h003F; B = 16'h00C7; #100;
A = 16'h003F; B = 16'h00C8; #100;
A = 16'h003F; B = 16'h00C9; #100;
A = 16'h003F; B = 16'h00CA; #100;
A = 16'h003F; B = 16'h00CB; #100;
A = 16'h003F; B = 16'h00CC; #100;
A = 16'h003F; B = 16'h00CD; #100;
A = 16'h003F; B = 16'h00CE; #100;
A = 16'h003F; B = 16'h00CF; #100;
A = 16'h003F; B = 16'h00D0; #100;
A = 16'h003F; B = 16'h00D1; #100;
A = 16'h003F; B = 16'h00D2; #100;
A = 16'h003F; B = 16'h00D3; #100;
A = 16'h003F; B = 16'h00D4; #100;
A = 16'h003F; B = 16'h00D5; #100;
A = 16'h003F; B = 16'h00D6; #100;
A = 16'h003F; B = 16'h00D7; #100;
A = 16'h003F; B = 16'h00D8; #100;
A = 16'h003F; B = 16'h00D9; #100;
A = 16'h003F; B = 16'h00DA; #100;
A = 16'h003F; B = 16'h00DB; #100;
A = 16'h003F; B = 16'h00DC; #100;
A = 16'h003F; B = 16'h00DD; #100;
A = 16'h003F; B = 16'h00DE; #100;
A = 16'h003F; B = 16'h00DF; #100;
A = 16'h003F; B = 16'h00E0; #100;
A = 16'h003F; B = 16'h00E1; #100;
A = 16'h003F; B = 16'h00E2; #100;
A = 16'h003F; B = 16'h00E3; #100;
A = 16'h003F; B = 16'h00E4; #100;
A = 16'h003F; B = 16'h00E5; #100;
A = 16'h003F; B = 16'h00E6; #100;
A = 16'h003F; B = 16'h00E7; #100;
A = 16'h003F; B = 16'h00E8; #100;
A = 16'h003F; B = 16'h00E9; #100;
A = 16'h003F; B = 16'h00EA; #100;
A = 16'h003F; B = 16'h00EB; #100;
A = 16'h003F; B = 16'h00EC; #100;
A = 16'h003F; B = 16'h00ED; #100;
A = 16'h003F; B = 16'h00EE; #100;
A = 16'h003F; B = 16'h00EF; #100;
A = 16'h003F; B = 16'h00F0; #100;
A = 16'h003F; B = 16'h00F1; #100;
A = 16'h003F; B = 16'h00F2; #100;
A = 16'h003F; B = 16'h00F3; #100;
A = 16'h003F; B = 16'h00F4; #100;
A = 16'h003F; B = 16'h00F5; #100;
A = 16'h003F; B = 16'h00F6; #100;
A = 16'h003F; B = 16'h00F7; #100;
A = 16'h003F; B = 16'h00F8; #100;
A = 16'h003F; B = 16'h00F9; #100;
A = 16'h003F; B = 16'h00FA; #100;
A = 16'h003F; B = 16'h00FB; #100;
A = 16'h003F; B = 16'h00FC; #100;
A = 16'h003F; B = 16'h00FD; #100;
A = 16'h003F; B = 16'h00FE; #100;
A = 16'h003F; B = 16'h00FF; #100;
A = 16'h0040; B = 16'h000; #100;
A = 16'h0040; B = 16'h001; #100;
A = 16'h0040; B = 16'h002; #100;
A = 16'h0040; B = 16'h003; #100;
A = 16'h0040; B = 16'h004; #100;
A = 16'h0040; B = 16'h005; #100;
A = 16'h0040; B = 16'h006; #100;
A = 16'h0040; B = 16'h007; #100;
A = 16'h0040; B = 16'h008; #100;
A = 16'h0040; B = 16'h009; #100;
A = 16'h0040; B = 16'h00A; #100;
A = 16'h0040; B = 16'h00B; #100;
A = 16'h0040; B = 16'h00C; #100;
A = 16'h0040; B = 16'h00D; #100;
A = 16'h0040; B = 16'h00E; #100;
A = 16'h0040; B = 16'h00F; #100;
A = 16'h0040; B = 16'h0010; #100;
A = 16'h0040; B = 16'h0011; #100;
A = 16'h0040; B = 16'h0012; #100;
A = 16'h0040; B = 16'h0013; #100;
A = 16'h0040; B = 16'h0014; #100;
A = 16'h0040; B = 16'h0015; #100;
A = 16'h0040; B = 16'h0016; #100;
A = 16'h0040; B = 16'h0017; #100;
A = 16'h0040; B = 16'h0018; #100;
A = 16'h0040; B = 16'h0019; #100;
A = 16'h0040; B = 16'h001A; #100;
A = 16'h0040; B = 16'h001B; #100;
A = 16'h0040; B = 16'h001C; #100;
A = 16'h0040; B = 16'h001D; #100;
A = 16'h0040; B = 16'h001E; #100;
A = 16'h0040; B = 16'h001F; #100;
A = 16'h0040; B = 16'h0020; #100;
A = 16'h0040; B = 16'h0021; #100;
A = 16'h0040; B = 16'h0022; #100;
A = 16'h0040; B = 16'h0023; #100;
A = 16'h0040; B = 16'h0024; #100;
A = 16'h0040; B = 16'h0025; #100;
A = 16'h0040; B = 16'h0026; #100;
A = 16'h0040; B = 16'h0027; #100;
A = 16'h0040; B = 16'h0028; #100;
A = 16'h0040; B = 16'h0029; #100;
A = 16'h0040; B = 16'h002A; #100;
A = 16'h0040; B = 16'h002B; #100;
A = 16'h0040; B = 16'h002C; #100;
A = 16'h0040; B = 16'h002D; #100;
A = 16'h0040; B = 16'h002E; #100;
A = 16'h0040; B = 16'h002F; #100;
A = 16'h0040; B = 16'h0030; #100;
A = 16'h0040; B = 16'h0031; #100;
A = 16'h0040; B = 16'h0032; #100;
A = 16'h0040; B = 16'h0033; #100;
A = 16'h0040; B = 16'h0034; #100;
A = 16'h0040; B = 16'h0035; #100;
A = 16'h0040; B = 16'h0036; #100;
A = 16'h0040; B = 16'h0037; #100;
A = 16'h0040; B = 16'h0038; #100;
A = 16'h0040; B = 16'h0039; #100;
A = 16'h0040; B = 16'h003A; #100;
A = 16'h0040; B = 16'h003B; #100;
A = 16'h0040; B = 16'h003C; #100;
A = 16'h0040; B = 16'h003D; #100;
A = 16'h0040; B = 16'h003E; #100;
A = 16'h0040; B = 16'h003F; #100;
A = 16'h0040; B = 16'h0040; #100;
A = 16'h0040; B = 16'h0041; #100;
A = 16'h0040; B = 16'h0042; #100;
A = 16'h0040; B = 16'h0043; #100;
A = 16'h0040; B = 16'h0044; #100;
A = 16'h0040; B = 16'h0045; #100;
A = 16'h0040; B = 16'h0046; #100;
A = 16'h0040; B = 16'h0047; #100;
A = 16'h0040; B = 16'h0048; #100;
A = 16'h0040; B = 16'h0049; #100;
A = 16'h0040; B = 16'h004A; #100;
A = 16'h0040; B = 16'h004B; #100;
A = 16'h0040; B = 16'h004C; #100;
A = 16'h0040; B = 16'h004D; #100;
A = 16'h0040; B = 16'h004E; #100;
A = 16'h0040; B = 16'h004F; #100;
A = 16'h0040; B = 16'h0050; #100;
A = 16'h0040; B = 16'h0051; #100;
A = 16'h0040; B = 16'h0052; #100;
A = 16'h0040; B = 16'h0053; #100;
A = 16'h0040; B = 16'h0054; #100;
A = 16'h0040; B = 16'h0055; #100;
A = 16'h0040; B = 16'h0056; #100;
A = 16'h0040; B = 16'h0057; #100;
A = 16'h0040; B = 16'h0058; #100;
A = 16'h0040; B = 16'h0059; #100;
A = 16'h0040; B = 16'h005A; #100;
A = 16'h0040; B = 16'h005B; #100;
A = 16'h0040; B = 16'h005C; #100;
A = 16'h0040; B = 16'h005D; #100;
A = 16'h0040; B = 16'h005E; #100;
A = 16'h0040; B = 16'h005F; #100;
A = 16'h0040; B = 16'h0060; #100;
A = 16'h0040; B = 16'h0061; #100;
A = 16'h0040; B = 16'h0062; #100;
A = 16'h0040; B = 16'h0063; #100;
A = 16'h0040; B = 16'h0064; #100;
A = 16'h0040; B = 16'h0065; #100;
A = 16'h0040; B = 16'h0066; #100;
A = 16'h0040; B = 16'h0067; #100;
A = 16'h0040; B = 16'h0068; #100;
A = 16'h0040; B = 16'h0069; #100;
A = 16'h0040; B = 16'h006A; #100;
A = 16'h0040; B = 16'h006B; #100;
A = 16'h0040; B = 16'h006C; #100;
A = 16'h0040; B = 16'h006D; #100;
A = 16'h0040; B = 16'h006E; #100;
A = 16'h0040; B = 16'h006F; #100;
A = 16'h0040; B = 16'h0070; #100;
A = 16'h0040; B = 16'h0071; #100;
A = 16'h0040; B = 16'h0072; #100;
A = 16'h0040; B = 16'h0073; #100;
A = 16'h0040; B = 16'h0074; #100;
A = 16'h0040; B = 16'h0075; #100;
A = 16'h0040; B = 16'h0076; #100;
A = 16'h0040; B = 16'h0077; #100;
A = 16'h0040; B = 16'h0078; #100;
A = 16'h0040; B = 16'h0079; #100;
A = 16'h0040; B = 16'h007A; #100;
A = 16'h0040; B = 16'h007B; #100;
A = 16'h0040; B = 16'h007C; #100;
A = 16'h0040; B = 16'h007D; #100;
A = 16'h0040; B = 16'h007E; #100;
A = 16'h0040; B = 16'h007F; #100;
A = 16'h0040; B = 16'h0080; #100;
A = 16'h0040; B = 16'h0081; #100;
A = 16'h0040; B = 16'h0082; #100;
A = 16'h0040; B = 16'h0083; #100;
A = 16'h0040; B = 16'h0084; #100;
A = 16'h0040; B = 16'h0085; #100;
A = 16'h0040; B = 16'h0086; #100;
A = 16'h0040; B = 16'h0087; #100;
A = 16'h0040; B = 16'h0088; #100;
A = 16'h0040; B = 16'h0089; #100;
A = 16'h0040; B = 16'h008A; #100;
A = 16'h0040; B = 16'h008B; #100;
A = 16'h0040; B = 16'h008C; #100;
A = 16'h0040; B = 16'h008D; #100;
A = 16'h0040; B = 16'h008E; #100;
A = 16'h0040; B = 16'h008F; #100;
A = 16'h0040; B = 16'h0090; #100;
A = 16'h0040; B = 16'h0091; #100;
A = 16'h0040; B = 16'h0092; #100;
A = 16'h0040; B = 16'h0093; #100;
A = 16'h0040; B = 16'h0094; #100;
A = 16'h0040; B = 16'h0095; #100;
A = 16'h0040; B = 16'h0096; #100;
A = 16'h0040; B = 16'h0097; #100;
A = 16'h0040; B = 16'h0098; #100;
A = 16'h0040; B = 16'h0099; #100;
A = 16'h0040; B = 16'h009A; #100;
A = 16'h0040; B = 16'h009B; #100;
A = 16'h0040; B = 16'h009C; #100;
A = 16'h0040; B = 16'h009D; #100;
A = 16'h0040; B = 16'h009E; #100;
A = 16'h0040; B = 16'h009F; #100;
A = 16'h0040; B = 16'h00A0; #100;
A = 16'h0040; B = 16'h00A1; #100;
A = 16'h0040; B = 16'h00A2; #100;
A = 16'h0040; B = 16'h00A3; #100;
A = 16'h0040; B = 16'h00A4; #100;
A = 16'h0040; B = 16'h00A5; #100;
A = 16'h0040; B = 16'h00A6; #100;
A = 16'h0040; B = 16'h00A7; #100;
A = 16'h0040; B = 16'h00A8; #100;
A = 16'h0040; B = 16'h00A9; #100;
A = 16'h0040; B = 16'h00AA; #100;
A = 16'h0040; B = 16'h00AB; #100;
A = 16'h0040; B = 16'h00AC; #100;
A = 16'h0040; B = 16'h00AD; #100;
A = 16'h0040; B = 16'h00AE; #100;
A = 16'h0040; B = 16'h00AF; #100;
A = 16'h0040; B = 16'h00B0; #100;
A = 16'h0040; B = 16'h00B1; #100;
A = 16'h0040; B = 16'h00B2; #100;
A = 16'h0040; B = 16'h00B3; #100;
A = 16'h0040; B = 16'h00B4; #100;
A = 16'h0040; B = 16'h00B5; #100;
A = 16'h0040; B = 16'h00B6; #100;
A = 16'h0040; B = 16'h00B7; #100;
A = 16'h0040; B = 16'h00B8; #100;
A = 16'h0040; B = 16'h00B9; #100;
A = 16'h0040; B = 16'h00BA; #100;
A = 16'h0040; B = 16'h00BB; #100;
A = 16'h0040; B = 16'h00BC; #100;
A = 16'h0040; B = 16'h00BD; #100;
A = 16'h0040; B = 16'h00BE; #100;
A = 16'h0040; B = 16'h00BF; #100;
A = 16'h0040; B = 16'h00C0; #100;
A = 16'h0040; B = 16'h00C1; #100;
A = 16'h0040; B = 16'h00C2; #100;
A = 16'h0040; B = 16'h00C3; #100;
A = 16'h0040; B = 16'h00C4; #100;
A = 16'h0040; B = 16'h00C5; #100;
A = 16'h0040; B = 16'h00C6; #100;
A = 16'h0040; B = 16'h00C7; #100;
A = 16'h0040; B = 16'h00C8; #100;
A = 16'h0040; B = 16'h00C9; #100;
A = 16'h0040; B = 16'h00CA; #100;
A = 16'h0040; B = 16'h00CB; #100;
A = 16'h0040; B = 16'h00CC; #100;
A = 16'h0040; B = 16'h00CD; #100;
A = 16'h0040; B = 16'h00CE; #100;
A = 16'h0040; B = 16'h00CF; #100;
A = 16'h0040; B = 16'h00D0; #100;
A = 16'h0040; B = 16'h00D1; #100;
A = 16'h0040; B = 16'h00D2; #100;
A = 16'h0040; B = 16'h00D3; #100;
A = 16'h0040; B = 16'h00D4; #100;
A = 16'h0040; B = 16'h00D5; #100;
A = 16'h0040; B = 16'h00D6; #100;
A = 16'h0040; B = 16'h00D7; #100;
A = 16'h0040; B = 16'h00D8; #100;
A = 16'h0040; B = 16'h00D9; #100;
A = 16'h0040; B = 16'h00DA; #100;
A = 16'h0040; B = 16'h00DB; #100;
A = 16'h0040; B = 16'h00DC; #100;
A = 16'h0040; B = 16'h00DD; #100;
A = 16'h0040; B = 16'h00DE; #100;
A = 16'h0040; B = 16'h00DF; #100;
A = 16'h0040; B = 16'h00E0; #100;
A = 16'h0040; B = 16'h00E1; #100;
A = 16'h0040; B = 16'h00E2; #100;
A = 16'h0040; B = 16'h00E3; #100;
A = 16'h0040; B = 16'h00E4; #100;
A = 16'h0040; B = 16'h00E5; #100;
A = 16'h0040; B = 16'h00E6; #100;
A = 16'h0040; B = 16'h00E7; #100;
A = 16'h0040; B = 16'h00E8; #100;
A = 16'h0040; B = 16'h00E9; #100;
A = 16'h0040; B = 16'h00EA; #100;
A = 16'h0040; B = 16'h00EB; #100;
A = 16'h0040; B = 16'h00EC; #100;
A = 16'h0040; B = 16'h00ED; #100;
A = 16'h0040; B = 16'h00EE; #100;
A = 16'h0040; B = 16'h00EF; #100;
A = 16'h0040; B = 16'h00F0; #100;
A = 16'h0040; B = 16'h00F1; #100;
A = 16'h0040; B = 16'h00F2; #100;
A = 16'h0040; B = 16'h00F3; #100;
A = 16'h0040; B = 16'h00F4; #100;
A = 16'h0040; B = 16'h00F5; #100;
A = 16'h0040; B = 16'h00F6; #100;
A = 16'h0040; B = 16'h00F7; #100;
A = 16'h0040; B = 16'h00F8; #100;
A = 16'h0040; B = 16'h00F9; #100;
A = 16'h0040; B = 16'h00FA; #100;
A = 16'h0040; B = 16'h00FB; #100;
A = 16'h0040; B = 16'h00FC; #100;
A = 16'h0040; B = 16'h00FD; #100;
A = 16'h0040; B = 16'h00FE; #100;
A = 16'h0040; B = 16'h00FF; #100;
A = 16'h0041; B = 16'h000; #100;
A = 16'h0041; B = 16'h001; #100;
A = 16'h0041; B = 16'h002; #100;
A = 16'h0041; B = 16'h003; #100;
A = 16'h0041; B = 16'h004; #100;
A = 16'h0041; B = 16'h005; #100;
A = 16'h0041; B = 16'h006; #100;
A = 16'h0041; B = 16'h007; #100;
A = 16'h0041; B = 16'h008; #100;
A = 16'h0041; B = 16'h009; #100;
A = 16'h0041; B = 16'h00A; #100;
A = 16'h0041; B = 16'h00B; #100;
A = 16'h0041; B = 16'h00C; #100;
A = 16'h0041; B = 16'h00D; #100;
A = 16'h0041; B = 16'h00E; #100;
A = 16'h0041; B = 16'h00F; #100;
A = 16'h0041; B = 16'h0010; #100;
A = 16'h0041; B = 16'h0011; #100;
A = 16'h0041; B = 16'h0012; #100;
A = 16'h0041; B = 16'h0013; #100;
A = 16'h0041; B = 16'h0014; #100;
A = 16'h0041; B = 16'h0015; #100;
A = 16'h0041; B = 16'h0016; #100;
A = 16'h0041; B = 16'h0017; #100;
A = 16'h0041; B = 16'h0018; #100;
A = 16'h0041; B = 16'h0019; #100;
A = 16'h0041; B = 16'h001A; #100;
A = 16'h0041; B = 16'h001B; #100;
A = 16'h0041; B = 16'h001C; #100;
A = 16'h0041; B = 16'h001D; #100;
A = 16'h0041; B = 16'h001E; #100;
A = 16'h0041; B = 16'h001F; #100;
A = 16'h0041; B = 16'h0020; #100;
A = 16'h0041; B = 16'h0021; #100;
A = 16'h0041; B = 16'h0022; #100;
A = 16'h0041; B = 16'h0023; #100;
A = 16'h0041; B = 16'h0024; #100;
A = 16'h0041; B = 16'h0025; #100;
A = 16'h0041; B = 16'h0026; #100;
A = 16'h0041; B = 16'h0027; #100;
A = 16'h0041; B = 16'h0028; #100;
A = 16'h0041; B = 16'h0029; #100;
A = 16'h0041; B = 16'h002A; #100;
A = 16'h0041; B = 16'h002B; #100;
A = 16'h0041; B = 16'h002C; #100;
A = 16'h0041; B = 16'h002D; #100;
A = 16'h0041; B = 16'h002E; #100;
A = 16'h0041; B = 16'h002F; #100;
A = 16'h0041; B = 16'h0030; #100;
A = 16'h0041; B = 16'h0031; #100;
A = 16'h0041; B = 16'h0032; #100;
A = 16'h0041; B = 16'h0033; #100;
A = 16'h0041; B = 16'h0034; #100;
A = 16'h0041; B = 16'h0035; #100;
A = 16'h0041; B = 16'h0036; #100;
A = 16'h0041; B = 16'h0037; #100;
A = 16'h0041; B = 16'h0038; #100;
A = 16'h0041; B = 16'h0039; #100;
A = 16'h0041; B = 16'h003A; #100;
A = 16'h0041; B = 16'h003B; #100;
A = 16'h0041; B = 16'h003C; #100;
A = 16'h0041; B = 16'h003D; #100;
A = 16'h0041; B = 16'h003E; #100;
A = 16'h0041; B = 16'h003F; #100;
A = 16'h0041; B = 16'h0040; #100;
A = 16'h0041; B = 16'h0041; #100;
A = 16'h0041; B = 16'h0042; #100;
A = 16'h0041; B = 16'h0043; #100;
A = 16'h0041; B = 16'h0044; #100;
A = 16'h0041; B = 16'h0045; #100;
A = 16'h0041; B = 16'h0046; #100;
A = 16'h0041; B = 16'h0047; #100;
A = 16'h0041; B = 16'h0048; #100;
A = 16'h0041; B = 16'h0049; #100;
A = 16'h0041; B = 16'h004A; #100;
A = 16'h0041; B = 16'h004B; #100;
A = 16'h0041; B = 16'h004C; #100;
A = 16'h0041; B = 16'h004D; #100;
A = 16'h0041; B = 16'h004E; #100;
A = 16'h0041; B = 16'h004F; #100;
A = 16'h0041; B = 16'h0050; #100;
A = 16'h0041; B = 16'h0051; #100;
A = 16'h0041; B = 16'h0052; #100;
A = 16'h0041; B = 16'h0053; #100;
A = 16'h0041; B = 16'h0054; #100;
A = 16'h0041; B = 16'h0055; #100;
A = 16'h0041; B = 16'h0056; #100;
A = 16'h0041; B = 16'h0057; #100;
A = 16'h0041; B = 16'h0058; #100;
A = 16'h0041; B = 16'h0059; #100;
A = 16'h0041; B = 16'h005A; #100;
A = 16'h0041; B = 16'h005B; #100;
A = 16'h0041; B = 16'h005C; #100;
A = 16'h0041; B = 16'h005D; #100;
A = 16'h0041; B = 16'h005E; #100;
A = 16'h0041; B = 16'h005F; #100;
A = 16'h0041; B = 16'h0060; #100;
A = 16'h0041; B = 16'h0061; #100;
A = 16'h0041; B = 16'h0062; #100;
A = 16'h0041; B = 16'h0063; #100;
A = 16'h0041; B = 16'h0064; #100;
A = 16'h0041; B = 16'h0065; #100;
A = 16'h0041; B = 16'h0066; #100;
A = 16'h0041; B = 16'h0067; #100;
A = 16'h0041; B = 16'h0068; #100;
A = 16'h0041; B = 16'h0069; #100;
A = 16'h0041; B = 16'h006A; #100;
A = 16'h0041; B = 16'h006B; #100;
A = 16'h0041; B = 16'h006C; #100;
A = 16'h0041; B = 16'h006D; #100;
A = 16'h0041; B = 16'h006E; #100;
A = 16'h0041; B = 16'h006F; #100;
A = 16'h0041; B = 16'h0070; #100;
A = 16'h0041; B = 16'h0071; #100;
A = 16'h0041; B = 16'h0072; #100;
A = 16'h0041; B = 16'h0073; #100;
A = 16'h0041; B = 16'h0074; #100;
A = 16'h0041; B = 16'h0075; #100;
A = 16'h0041; B = 16'h0076; #100;
A = 16'h0041; B = 16'h0077; #100;
A = 16'h0041; B = 16'h0078; #100;
A = 16'h0041; B = 16'h0079; #100;
A = 16'h0041; B = 16'h007A; #100;
A = 16'h0041; B = 16'h007B; #100;
A = 16'h0041; B = 16'h007C; #100;
A = 16'h0041; B = 16'h007D; #100;
A = 16'h0041; B = 16'h007E; #100;
A = 16'h0041; B = 16'h007F; #100;
A = 16'h0041; B = 16'h0080; #100;
A = 16'h0041; B = 16'h0081; #100;
A = 16'h0041; B = 16'h0082; #100;
A = 16'h0041; B = 16'h0083; #100;
A = 16'h0041; B = 16'h0084; #100;
A = 16'h0041; B = 16'h0085; #100;
A = 16'h0041; B = 16'h0086; #100;
A = 16'h0041; B = 16'h0087; #100;
A = 16'h0041; B = 16'h0088; #100;
A = 16'h0041; B = 16'h0089; #100;
A = 16'h0041; B = 16'h008A; #100;
A = 16'h0041; B = 16'h008B; #100;
A = 16'h0041; B = 16'h008C; #100;
A = 16'h0041; B = 16'h008D; #100;
A = 16'h0041; B = 16'h008E; #100;
A = 16'h0041; B = 16'h008F; #100;
A = 16'h0041; B = 16'h0090; #100;
A = 16'h0041; B = 16'h0091; #100;
A = 16'h0041; B = 16'h0092; #100;
A = 16'h0041; B = 16'h0093; #100;
A = 16'h0041; B = 16'h0094; #100;
A = 16'h0041; B = 16'h0095; #100;
A = 16'h0041; B = 16'h0096; #100;
A = 16'h0041; B = 16'h0097; #100;
A = 16'h0041; B = 16'h0098; #100;
A = 16'h0041; B = 16'h0099; #100;
A = 16'h0041; B = 16'h009A; #100;
A = 16'h0041; B = 16'h009B; #100;
A = 16'h0041; B = 16'h009C; #100;
A = 16'h0041; B = 16'h009D; #100;
A = 16'h0041; B = 16'h009E; #100;
A = 16'h0041; B = 16'h009F; #100;
A = 16'h0041; B = 16'h00A0; #100;
A = 16'h0041; B = 16'h00A1; #100;
A = 16'h0041; B = 16'h00A2; #100;
A = 16'h0041; B = 16'h00A3; #100;
A = 16'h0041; B = 16'h00A4; #100;
A = 16'h0041; B = 16'h00A5; #100;
A = 16'h0041; B = 16'h00A6; #100;
A = 16'h0041; B = 16'h00A7; #100;
A = 16'h0041; B = 16'h00A8; #100;
A = 16'h0041; B = 16'h00A9; #100;
A = 16'h0041; B = 16'h00AA; #100;
A = 16'h0041; B = 16'h00AB; #100;
A = 16'h0041; B = 16'h00AC; #100;
A = 16'h0041; B = 16'h00AD; #100;
A = 16'h0041; B = 16'h00AE; #100;
A = 16'h0041; B = 16'h00AF; #100;
A = 16'h0041; B = 16'h00B0; #100;
A = 16'h0041; B = 16'h00B1; #100;
A = 16'h0041; B = 16'h00B2; #100;
A = 16'h0041; B = 16'h00B3; #100;
A = 16'h0041; B = 16'h00B4; #100;
A = 16'h0041; B = 16'h00B5; #100;
A = 16'h0041; B = 16'h00B6; #100;
A = 16'h0041; B = 16'h00B7; #100;
A = 16'h0041; B = 16'h00B8; #100;
A = 16'h0041; B = 16'h00B9; #100;
A = 16'h0041; B = 16'h00BA; #100;
A = 16'h0041; B = 16'h00BB; #100;
A = 16'h0041; B = 16'h00BC; #100;
A = 16'h0041; B = 16'h00BD; #100;
A = 16'h0041; B = 16'h00BE; #100;
A = 16'h0041; B = 16'h00BF; #100;
A = 16'h0041; B = 16'h00C0; #100;
A = 16'h0041; B = 16'h00C1; #100;
A = 16'h0041; B = 16'h00C2; #100;
A = 16'h0041; B = 16'h00C3; #100;
A = 16'h0041; B = 16'h00C4; #100;
A = 16'h0041; B = 16'h00C5; #100;
A = 16'h0041; B = 16'h00C6; #100;
A = 16'h0041; B = 16'h00C7; #100;
A = 16'h0041; B = 16'h00C8; #100;
A = 16'h0041; B = 16'h00C9; #100;
A = 16'h0041; B = 16'h00CA; #100;
A = 16'h0041; B = 16'h00CB; #100;
A = 16'h0041; B = 16'h00CC; #100;
A = 16'h0041; B = 16'h00CD; #100;
A = 16'h0041; B = 16'h00CE; #100;
A = 16'h0041; B = 16'h00CF; #100;
A = 16'h0041; B = 16'h00D0; #100;
A = 16'h0041; B = 16'h00D1; #100;
A = 16'h0041; B = 16'h00D2; #100;
A = 16'h0041; B = 16'h00D3; #100;
A = 16'h0041; B = 16'h00D4; #100;
A = 16'h0041; B = 16'h00D5; #100;
A = 16'h0041; B = 16'h00D6; #100;
A = 16'h0041; B = 16'h00D7; #100;
A = 16'h0041; B = 16'h00D8; #100;
A = 16'h0041; B = 16'h00D9; #100;
A = 16'h0041; B = 16'h00DA; #100;
A = 16'h0041; B = 16'h00DB; #100;
A = 16'h0041; B = 16'h00DC; #100;
A = 16'h0041; B = 16'h00DD; #100;
A = 16'h0041; B = 16'h00DE; #100;
A = 16'h0041; B = 16'h00DF; #100;
A = 16'h0041; B = 16'h00E0; #100;
A = 16'h0041; B = 16'h00E1; #100;
A = 16'h0041; B = 16'h00E2; #100;
A = 16'h0041; B = 16'h00E3; #100;
A = 16'h0041; B = 16'h00E4; #100;
A = 16'h0041; B = 16'h00E5; #100;
A = 16'h0041; B = 16'h00E6; #100;
A = 16'h0041; B = 16'h00E7; #100;
A = 16'h0041; B = 16'h00E8; #100;
A = 16'h0041; B = 16'h00E9; #100;
A = 16'h0041; B = 16'h00EA; #100;
A = 16'h0041; B = 16'h00EB; #100;
A = 16'h0041; B = 16'h00EC; #100;
A = 16'h0041; B = 16'h00ED; #100;
A = 16'h0041; B = 16'h00EE; #100;
A = 16'h0041; B = 16'h00EF; #100;
A = 16'h0041; B = 16'h00F0; #100;
A = 16'h0041; B = 16'h00F1; #100;
A = 16'h0041; B = 16'h00F2; #100;
A = 16'h0041; B = 16'h00F3; #100;
A = 16'h0041; B = 16'h00F4; #100;
A = 16'h0041; B = 16'h00F5; #100;
A = 16'h0041; B = 16'h00F6; #100;
A = 16'h0041; B = 16'h00F7; #100;
A = 16'h0041; B = 16'h00F8; #100;
A = 16'h0041; B = 16'h00F9; #100;
A = 16'h0041; B = 16'h00FA; #100;
A = 16'h0041; B = 16'h00FB; #100;
A = 16'h0041; B = 16'h00FC; #100;
A = 16'h0041; B = 16'h00FD; #100;
A = 16'h0041; B = 16'h00FE; #100;
A = 16'h0041; B = 16'h00FF; #100;
A = 16'h0042; B = 16'h000; #100;
A = 16'h0042; B = 16'h001; #100;
A = 16'h0042; B = 16'h002; #100;
A = 16'h0042; B = 16'h003; #100;
A = 16'h0042; B = 16'h004; #100;
A = 16'h0042; B = 16'h005; #100;
A = 16'h0042; B = 16'h006; #100;
A = 16'h0042; B = 16'h007; #100;
A = 16'h0042; B = 16'h008; #100;
A = 16'h0042; B = 16'h009; #100;
A = 16'h0042; B = 16'h00A; #100;
A = 16'h0042; B = 16'h00B; #100;
A = 16'h0042; B = 16'h00C; #100;
A = 16'h0042; B = 16'h00D; #100;
A = 16'h0042; B = 16'h00E; #100;
A = 16'h0042; B = 16'h00F; #100;
A = 16'h0042; B = 16'h0010; #100;
A = 16'h0042; B = 16'h0011; #100;
A = 16'h0042; B = 16'h0012; #100;
A = 16'h0042; B = 16'h0013; #100;
A = 16'h0042; B = 16'h0014; #100;
A = 16'h0042; B = 16'h0015; #100;
A = 16'h0042; B = 16'h0016; #100;
A = 16'h0042; B = 16'h0017; #100;
A = 16'h0042; B = 16'h0018; #100;
A = 16'h0042; B = 16'h0019; #100;
A = 16'h0042; B = 16'h001A; #100;
A = 16'h0042; B = 16'h001B; #100;
A = 16'h0042; B = 16'h001C; #100;
A = 16'h0042; B = 16'h001D; #100;
A = 16'h0042; B = 16'h001E; #100;
A = 16'h0042; B = 16'h001F; #100;
A = 16'h0042; B = 16'h0020; #100;
A = 16'h0042; B = 16'h0021; #100;
A = 16'h0042; B = 16'h0022; #100;
A = 16'h0042; B = 16'h0023; #100;
A = 16'h0042; B = 16'h0024; #100;
A = 16'h0042; B = 16'h0025; #100;
A = 16'h0042; B = 16'h0026; #100;
A = 16'h0042; B = 16'h0027; #100;
A = 16'h0042; B = 16'h0028; #100;
A = 16'h0042; B = 16'h0029; #100;
A = 16'h0042; B = 16'h002A; #100;
A = 16'h0042; B = 16'h002B; #100;
A = 16'h0042; B = 16'h002C; #100;
A = 16'h0042; B = 16'h002D; #100;
A = 16'h0042; B = 16'h002E; #100;
A = 16'h0042; B = 16'h002F; #100;
A = 16'h0042; B = 16'h0030; #100;
A = 16'h0042; B = 16'h0031; #100;
A = 16'h0042; B = 16'h0032; #100;
A = 16'h0042; B = 16'h0033; #100;
A = 16'h0042; B = 16'h0034; #100;
A = 16'h0042; B = 16'h0035; #100;
A = 16'h0042; B = 16'h0036; #100;
A = 16'h0042; B = 16'h0037; #100;
A = 16'h0042; B = 16'h0038; #100;
A = 16'h0042; B = 16'h0039; #100;
A = 16'h0042; B = 16'h003A; #100;
A = 16'h0042; B = 16'h003B; #100;
A = 16'h0042; B = 16'h003C; #100;
A = 16'h0042; B = 16'h003D; #100;
A = 16'h0042; B = 16'h003E; #100;
A = 16'h0042; B = 16'h003F; #100;
A = 16'h0042; B = 16'h0040; #100;
A = 16'h0042; B = 16'h0041; #100;
A = 16'h0042; B = 16'h0042; #100;
A = 16'h0042; B = 16'h0043; #100;
A = 16'h0042; B = 16'h0044; #100;
A = 16'h0042; B = 16'h0045; #100;
A = 16'h0042; B = 16'h0046; #100;
A = 16'h0042; B = 16'h0047; #100;
A = 16'h0042; B = 16'h0048; #100;
A = 16'h0042; B = 16'h0049; #100;
A = 16'h0042; B = 16'h004A; #100;
A = 16'h0042; B = 16'h004B; #100;
A = 16'h0042; B = 16'h004C; #100;
A = 16'h0042; B = 16'h004D; #100;
A = 16'h0042; B = 16'h004E; #100;
A = 16'h0042; B = 16'h004F; #100;
A = 16'h0042; B = 16'h0050; #100;
A = 16'h0042; B = 16'h0051; #100;
A = 16'h0042; B = 16'h0052; #100;
A = 16'h0042; B = 16'h0053; #100;
A = 16'h0042; B = 16'h0054; #100;
A = 16'h0042; B = 16'h0055; #100;
A = 16'h0042; B = 16'h0056; #100;
A = 16'h0042; B = 16'h0057; #100;
A = 16'h0042; B = 16'h0058; #100;
A = 16'h0042; B = 16'h0059; #100;
A = 16'h0042; B = 16'h005A; #100;
A = 16'h0042; B = 16'h005B; #100;
A = 16'h0042; B = 16'h005C; #100;
A = 16'h0042; B = 16'h005D; #100;
A = 16'h0042; B = 16'h005E; #100;
A = 16'h0042; B = 16'h005F; #100;
A = 16'h0042; B = 16'h0060; #100;
A = 16'h0042; B = 16'h0061; #100;
A = 16'h0042; B = 16'h0062; #100;
A = 16'h0042; B = 16'h0063; #100;
A = 16'h0042; B = 16'h0064; #100;
A = 16'h0042; B = 16'h0065; #100;
A = 16'h0042; B = 16'h0066; #100;
A = 16'h0042; B = 16'h0067; #100;
A = 16'h0042; B = 16'h0068; #100;
A = 16'h0042; B = 16'h0069; #100;
A = 16'h0042; B = 16'h006A; #100;
A = 16'h0042; B = 16'h006B; #100;
A = 16'h0042; B = 16'h006C; #100;
A = 16'h0042; B = 16'h006D; #100;
A = 16'h0042; B = 16'h006E; #100;
A = 16'h0042; B = 16'h006F; #100;
A = 16'h0042; B = 16'h0070; #100;
A = 16'h0042; B = 16'h0071; #100;
A = 16'h0042; B = 16'h0072; #100;
A = 16'h0042; B = 16'h0073; #100;
A = 16'h0042; B = 16'h0074; #100;
A = 16'h0042; B = 16'h0075; #100;
A = 16'h0042; B = 16'h0076; #100;
A = 16'h0042; B = 16'h0077; #100;
A = 16'h0042; B = 16'h0078; #100;
A = 16'h0042; B = 16'h0079; #100;
A = 16'h0042; B = 16'h007A; #100;
A = 16'h0042; B = 16'h007B; #100;
A = 16'h0042; B = 16'h007C; #100;
A = 16'h0042; B = 16'h007D; #100;
A = 16'h0042; B = 16'h007E; #100;
A = 16'h0042; B = 16'h007F; #100;
A = 16'h0042; B = 16'h0080; #100;
A = 16'h0042; B = 16'h0081; #100;
A = 16'h0042; B = 16'h0082; #100;
A = 16'h0042; B = 16'h0083; #100;
A = 16'h0042; B = 16'h0084; #100;
A = 16'h0042; B = 16'h0085; #100;
A = 16'h0042; B = 16'h0086; #100;
A = 16'h0042; B = 16'h0087; #100;
A = 16'h0042; B = 16'h0088; #100;
A = 16'h0042; B = 16'h0089; #100;
A = 16'h0042; B = 16'h008A; #100;
A = 16'h0042; B = 16'h008B; #100;
A = 16'h0042; B = 16'h008C; #100;
A = 16'h0042; B = 16'h008D; #100;
A = 16'h0042; B = 16'h008E; #100;
A = 16'h0042; B = 16'h008F; #100;
A = 16'h0042; B = 16'h0090; #100;
A = 16'h0042; B = 16'h0091; #100;
A = 16'h0042; B = 16'h0092; #100;
A = 16'h0042; B = 16'h0093; #100;
A = 16'h0042; B = 16'h0094; #100;
A = 16'h0042; B = 16'h0095; #100;
A = 16'h0042; B = 16'h0096; #100;
A = 16'h0042; B = 16'h0097; #100;
A = 16'h0042; B = 16'h0098; #100;
A = 16'h0042; B = 16'h0099; #100;
A = 16'h0042; B = 16'h009A; #100;
A = 16'h0042; B = 16'h009B; #100;
A = 16'h0042; B = 16'h009C; #100;
A = 16'h0042; B = 16'h009D; #100;
A = 16'h0042; B = 16'h009E; #100;
A = 16'h0042; B = 16'h009F; #100;
A = 16'h0042; B = 16'h00A0; #100;
A = 16'h0042; B = 16'h00A1; #100;
A = 16'h0042; B = 16'h00A2; #100;
A = 16'h0042; B = 16'h00A3; #100;
A = 16'h0042; B = 16'h00A4; #100;
A = 16'h0042; B = 16'h00A5; #100;
A = 16'h0042; B = 16'h00A6; #100;
A = 16'h0042; B = 16'h00A7; #100;
A = 16'h0042; B = 16'h00A8; #100;
A = 16'h0042; B = 16'h00A9; #100;
A = 16'h0042; B = 16'h00AA; #100;
A = 16'h0042; B = 16'h00AB; #100;
A = 16'h0042; B = 16'h00AC; #100;
A = 16'h0042; B = 16'h00AD; #100;
A = 16'h0042; B = 16'h00AE; #100;
A = 16'h0042; B = 16'h00AF; #100;
A = 16'h0042; B = 16'h00B0; #100;
A = 16'h0042; B = 16'h00B1; #100;
A = 16'h0042; B = 16'h00B2; #100;
A = 16'h0042; B = 16'h00B3; #100;
A = 16'h0042; B = 16'h00B4; #100;
A = 16'h0042; B = 16'h00B5; #100;
A = 16'h0042; B = 16'h00B6; #100;
A = 16'h0042; B = 16'h00B7; #100;
A = 16'h0042; B = 16'h00B8; #100;
A = 16'h0042; B = 16'h00B9; #100;
A = 16'h0042; B = 16'h00BA; #100;
A = 16'h0042; B = 16'h00BB; #100;
A = 16'h0042; B = 16'h00BC; #100;
A = 16'h0042; B = 16'h00BD; #100;
A = 16'h0042; B = 16'h00BE; #100;
A = 16'h0042; B = 16'h00BF; #100;
A = 16'h0042; B = 16'h00C0; #100;
A = 16'h0042; B = 16'h00C1; #100;
A = 16'h0042; B = 16'h00C2; #100;
A = 16'h0042; B = 16'h00C3; #100;
A = 16'h0042; B = 16'h00C4; #100;
A = 16'h0042; B = 16'h00C5; #100;
A = 16'h0042; B = 16'h00C6; #100;
A = 16'h0042; B = 16'h00C7; #100;
A = 16'h0042; B = 16'h00C8; #100;
A = 16'h0042; B = 16'h00C9; #100;
A = 16'h0042; B = 16'h00CA; #100;
A = 16'h0042; B = 16'h00CB; #100;
A = 16'h0042; B = 16'h00CC; #100;
A = 16'h0042; B = 16'h00CD; #100;
A = 16'h0042; B = 16'h00CE; #100;
A = 16'h0042; B = 16'h00CF; #100;
A = 16'h0042; B = 16'h00D0; #100;
A = 16'h0042; B = 16'h00D1; #100;
A = 16'h0042; B = 16'h00D2; #100;
A = 16'h0042; B = 16'h00D3; #100;
A = 16'h0042; B = 16'h00D4; #100;
A = 16'h0042; B = 16'h00D5; #100;
A = 16'h0042; B = 16'h00D6; #100;
A = 16'h0042; B = 16'h00D7; #100;
A = 16'h0042; B = 16'h00D8; #100;
A = 16'h0042; B = 16'h00D9; #100;
A = 16'h0042; B = 16'h00DA; #100;
A = 16'h0042; B = 16'h00DB; #100;
A = 16'h0042; B = 16'h00DC; #100;
A = 16'h0042; B = 16'h00DD; #100;
A = 16'h0042; B = 16'h00DE; #100;
A = 16'h0042; B = 16'h00DF; #100;
A = 16'h0042; B = 16'h00E0; #100;
A = 16'h0042; B = 16'h00E1; #100;
A = 16'h0042; B = 16'h00E2; #100;
A = 16'h0042; B = 16'h00E3; #100;
A = 16'h0042; B = 16'h00E4; #100;
A = 16'h0042; B = 16'h00E5; #100;
A = 16'h0042; B = 16'h00E6; #100;
A = 16'h0042; B = 16'h00E7; #100;
A = 16'h0042; B = 16'h00E8; #100;
A = 16'h0042; B = 16'h00E9; #100;
A = 16'h0042; B = 16'h00EA; #100;
A = 16'h0042; B = 16'h00EB; #100;
A = 16'h0042; B = 16'h00EC; #100;
A = 16'h0042; B = 16'h00ED; #100;
A = 16'h0042; B = 16'h00EE; #100;
A = 16'h0042; B = 16'h00EF; #100;
A = 16'h0042; B = 16'h00F0; #100;
A = 16'h0042; B = 16'h00F1; #100;
A = 16'h0042; B = 16'h00F2; #100;
A = 16'h0042; B = 16'h00F3; #100;
A = 16'h0042; B = 16'h00F4; #100;
A = 16'h0042; B = 16'h00F5; #100;
A = 16'h0042; B = 16'h00F6; #100;
A = 16'h0042; B = 16'h00F7; #100;
A = 16'h0042; B = 16'h00F8; #100;
A = 16'h0042; B = 16'h00F9; #100;
A = 16'h0042; B = 16'h00FA; #100;
A = 16'h0042; B = 16'h00FB; #100;
A = 16'h0042; B = 16'h00FC; #100;
A = 16'h0042; B = 16'h00FD; #100;
A = 16'h0042; B = 16'h00FE; #100;
A = 16'h0042; B = 16'h00FF; #100;
A = 16'h0043; B = 16'h000; #100;
A = 16'h0043; B = 16'h001; #100;
A = 16'h0043; B = 16'h002; #100;
A = 16'h0043; B = 16'h003; #100;
A = 16'h0043; B = 16'h004; #100;
A = 16'h0043; B = 16'h005; #100;
A = 16'h0043; B = 16'h006; #100;
A = 16'h0043; B = 16'h007; #100;
A = 16'h0043; B = 16'h008; #100;
A = 16'h0043; B = 16'h009; #100;
A = 16'h0043; B = 16'h00A; #100;
A = 16'h0043; B = 16'h00B; #100;
A = 16'h0043; B = 16'h00C; #100;
A = 16'h0043; B = 16'h00D; #100;
A = 16'h0043; B = 16'h00E; #100;
A = 16'h0043; B = 16'h00F; #100;
A = 16'h0043; B = 16'h0010; #100;
A = 16'h0043; B = 16'h0011; #100;
A = 16'h0043; B = 16'h0012; #100;
A = 16'h0043; B = 16'h0013; #100;
A = 16'h0043; B = 16'h0014; #100;
A = 16'h0043; B = 16'h0015; #100;
A = 16'h0043; B = 16'h0016; #100;
A = 16'h0043; B = 16'h0017; #100;
A = 16'h0043; B = 16'h0018; #100;
A = 16'h0043; B = 16'h0019; #100;
A = 16'h0043; B = 16'h001A; #100;
A = 16'h0043; B = 16'h001B; #100;
A = 16'h0043; B = 16'h001C; #100;
A = 16'h0043; B = 16'h001D; #100;
A = 16'h0043; B = 16'h001E; #100;
A = 16'h0043; B = 16'h001F; #100;
A = 16'h0043; B = 16'h0020; #100;
A = 16'h0043; B = 16'h0021; #100;
A = 16'h0043; B = 16'h0022; #100;
A = 16'h0043; B = 16'h0023; #100;
A = 16'h0043; B = 16'h0024; #100;
A = 16'h0043; B = 16'h0025; #100;
A = 16'h0043; B = 16'h0026; #100;
A = 16'h0043; B = 16'h0027; #100;
A = 16'h0043; B = 16'h0028; #100;
A = 16'h0043; B = 16'h0029; #100;
A = 16'h0043; B = 16'h002A; #100;
A = 16'h0043; B = 16'h002B; #100;
A = 16'h0043; B = 16'h002C; #100;
A = 16'h0043; B = 16'h002D; #100;
A = 16'h0043; B = 16'h002E; #100;
A = 16'h0043; B = 16'h002F; #100;
A = 16'h0043; B = 16'h0030; #100;
A = 16'h0043; B = 16'h0031; #100;
A = 16'h0043; B = 16'h0032; #100;
A = 16'h0043; B = 16'h0033; #100;
A = 16'h0043; B = 16'h0034; #100;
A = 16'h0043; B = 16'h0035; #100;
A = 16'h0043; B = 16'h0036; #100;
A = 16'h0043; B = 16'h0037; #100;
A = 16'h0043; B = 16'h0038; #100;
A = 16'h0043; B = 16'h0039; #100;
A = 16'h0043; B = 16'h003A; #100;
A = 16'h0043; B = 16'h003B; #100;
A = 16'h0043; B = 16'h003C; #100;
A = 16'h0043; B = 16'h003D; #100;
A = 16'h0043; B = 16'h003E; #100;
A = 16'h0043; B = 16'h003F; #100;
A = 16'h0043; B = 16'h0040; #100;
A = 16'h0043; B = 16'h0041; #100;
A = 16'h0043; B = 16'h0042; #100;
A = 16'h0043; B = 16'h0043; #100;
A = 16'h0043; B = 16'h0044; #100;
A = 16'h0043; B = 16'h0045; #100;
A = 16'h0043; B = 16'h0046; #100;
A = 16'h0043; B = 16'h0047; #100;
A = 16'h0043; B = 16'h0048; #100;
A = 16'h0043; B = 16'h0049; #100;
A = 16'h0043; B = 16'h004A; #100;
A = 16'h0043; B = 16'h004B; #100;
A = 16'h0043; B = 16'h004C; #100;
A = 16'h0043; B = 16'h004D; #100;
A = 16'h0043; B = 16'h004E; #100;
A = 16'h0043; B = 16'h004F; #100;
A = 16'h0043; B = 16'h0050; #100;
A = 16'h0043; B = 16'h0051; #100;
A = 16'h0043; B = 16'h0052; #100;
A = 16'h0043; B = 16'h0053; #100;
A = 16'h0043; B = 16'h0054; #100;
A = 16'h0043; B = 16'h0055; #100;
A = 16'h0043; B = 16'h0056; #100;
A = 16'h0043; B = 16'h0057; #100;
A = 16'h0043; B = 16'h0058; #100;
A = 16'h0043; B = 16'h0059; #100;
A = 16'h0043; B = 16'h005A; #100;
A = 16'h0043; B = 16'h005B; #100;
A = 16'h0043; B = 16'h005C; #100;
A = 16'h0043; B = 16'h005D; #100;
A = 16'h0043; B = 16'h005E; #100;
A = 16'h0043; B = 16'h005F; #100;
A = 16'h0043; B = 16'h0060; #100;
A = 16'h0043; B = 16'h0061; #100;
A = 16'h0043; B = 16'h0062; #100;
A = 16'h0043; B = 16'h0063; #100;
A = 16'h0043; B = 16'h0064; #100;
A = 16'h0043; B = 16'h0065; #100;
A = 16'h0043; B = 16'h0066; #100;
A = 16'h0043; B = 16'h0067; #100;
A = 16'h0043; B = 16'h0068; #100;
A = 16'h0043; B = 16'h0069; #100;
A = 16'h0043; B = 16'h006A; #100;
A = 16'h0043; B = 16'h006B; #100;
A = 16'h0043; B = 16'h006C; #100;
A = 16'h0043; B = 16'h006D; #100;
A = 16'h0043; B = 16'h006E; #100;
A = 16'h0043; B = 16'h006F; #100;
A = 16'h0043; B = 16'h0070; #100;
A = 16'h0043; B = 16'h0071; #100;
A = 16'h0043; B = 16'h0072; #100;
A = 16'h0043; B = 16'h0073; #100;
A = 16'h0043; B = 16'h0074; #100;
A = 16'h0043; B = 16'h0075; #100;
A = 16'h0043; B = 16'h0076; #100;
A = 16'h0043; B = 16'h0077; #100;
A = 16'h0043; B = 16'h0078; #100;
A = 16'h0043; B = 16'h0079; #100;
A = 16'h0043; B = 16'h007A; #100;
A = 16'h0043; B = 16'h007B; #100;
A = 16'h0043; B = 16'h007C; #100;
A = 16'h0043; B = 16'h007D; #100;
A = 16'h0043; B = 16'h007E; #100;
A = 16'h0043; B = 16'h007F; #100;
A = 16'h0043; B = 16'h0080; #100;
A = 16'h0043; B = 16'h0081; #100;
A = 16'h0043; B = 16'h0082; #100;
A = 16'h0043; B = 16'h0083; #100;
A = 16'h0043; B = 16'h0084; #100;
A = 16'h0043; B = 16'h0085; #100;
A = 16'h0043; B = 16'h0086; #100;
A = 16'h0043; B = 16'h0087; #100;
A = 16'h0043; B = 16'h0088; #100;
A = 16'h0043; B = 16'h0089; #100;
A = 16'h0043; B = 16'h008A; #100;
A = 16'h0043; B = 16'h008B; #100;
A = 16'h0043; B = 16'h008C; #100;
A = 16'h0043; B = 16'h008D; #100;
A = 16'h0043; B = 16'h008E; #100;
A = 16'h0043; B = 16'h008F; #100;
A = 16'h0043; B = 16'h0090; #100;
A = 16'h0043; B = 16'h0091; #100;
A = 16'h0043; B = 16'h0092; #100;
A = 16'h0043; B = 16'h0093; #100;
A = 16'h0043; B = 16'h0094; #100;
A = 16'h0043; B = 16'h0095; #100;
A = 16'h0043; B = 16'h0096; #100;
A = 16'h0043; B = 16'h0097; #100;
A = 16'h0043; B = 16'h0098; #100;
A = 16'h0043; B = 16'h0099; #100;
A = 16'h0043; B = 16'h009A; #100;
A = 16'h0043; B = 16'h009B; #100;
A = 16'h0043; B = 16'h009C; #100;
A = 16'h0043; B = 16'h009D; #100;
A = 16'h0043; B = 16'h009E; #100;
A = 16'h0043; B = 16'h009F; #100;
A = 16'h0043; B = 16'h00A0; #100;
A = 16'h0043; B = 16'h00A1; #100;
A = 16'h0043; B = 16'h00A2; #100;
A = 16'h0043; B = 16'h00A3; #100;
A = 16'h0043; B = 16'h00A4; #100;
A = 16'h0043; B = 16'h00A5; #100;
A = 16'h0043; B = 16'h00A6; #100;
A = 16'h0043; B = 16'h00A7; #100;
A = 16'h0043; B = 16'h00A8; #100;
A = 16'h0043; B = 16'h00A9; #100;
A = 16'h0043; B = 16'h00AA; #100;
A = 16'h0043; B = 16'h00AB; #100;
A = 16'h0043; B = 16'h00AC; #100;
A = 16'h0043; B = 16'h00AD; #100;
A = 16'h0043; B = 16'h00AE; #100;
A = 16'h0043; B = 16'h00AF; #100;
A = 16'h0043; B = 16'h00B0; #100;
A = 16'h0043; B = 16'h00B1; #100;
A = 16'h0043; B = 16'h00B2; #100;
A = 16'h0043; B = 16'h00B3; #100;
A = 16'h0043; B = 16'h00B4; #100;
A = 16'h0043; B = 16'h00B5; #100;
A = 16'h0043; B = 16'h00B6; #100;
A = 16'h0043; B = 16'h00B7; #100;
A = 16'h0043; B = 16'h00B8; #100;
A = 16'h0043; B = 16'h00B9; #100;
A = 16'h0043; B = 16'h00BA; #100;
A = 16'h0043; B = 16'h00BB; #100;
A = 16'h0043; B = 16'h00BC; #100;
A = 16'h0043; B = 16'h00BD; #100;
A = 16'h0043; B = 16'h00BE; #100;
A = 16'h0043; B = 16'h00BF; #100;
A = 16'h0043; B = 16'h00C0; #100;
A = 16'h0043; B = 16'h00C1; #100;
A = 16'h0043; B = 16'h00C2; #100;
A = 16'h0043; B = 16'h00C3; #100;
A = 16'h0043; B = 16'h00C4; #100;
A = 16'h0043; B = 16'h00C5; #100;
A = 16'h0043; B = 16'h00C6; #100;
A = 16'h0043; B = 16'h00C7; #100;
A = 16'h0043; B = 16'h00C8; #100;
A = 16'h0043; B = 16'h00C9; #100;
A = 16'h0043; B = 16'h00CA; #100;
A = 16'h0043; B = 16'h00CB; #100;
A = 16'h0043; B = 16'h00CC; #100;
A = 16'h0043; B = 16'h00CD; #100;
A = 16'h0043; B = 16'h00CE; #100;
A = 16'h0043; B = 16'h00CF; #100;
A = 16'h0043; B = 16'h00D0; #100;
A = 16'h0043; B = 16'h00D1; #100;
A = 16'h0043; B = 16'h00D2; #100;
A = 16'h0043; B = 16'h00D3; #100;
A = 16'h0043; B = 16'h00D4; #100;
A = 16'h0043; B = 16'h00D5; #100;
A = 16'h0043; B = 16'h00D6; #100;
A = 16'h0043; B = 16'h00D7; #100;
A = 16'h0043; B = 16'h00D8; #100;
A = 16'h0043; B = 16'h00D9; #100;
A = 16'h0043; B = 16'h00DA; #100;
A = 16'h0043; B = 16'h00DB; #100;
A = 16'h0043; B = 16'h00DC; #100;
A = 16'h0043; B = 16'h00DD; #100;
A = 16'h0043; B = 16'h00DE; #100;
A = 16'h0043; B = 16'h00DF; #100;
A = 16'h0043; B = 16'h00E0; #100;
A = 16'h0043; B = 16'h00E1; #100;
A = 16'h0043; B = 16'h00E2; #100;
A = 16'h0043; B = 16'h00E3; #100;
A = 16'h0043; B = 16'h00E4; #100;
A = 16'h0043; B = 16'h00E5; #100;
A = 16'h0043; B = 16'h00E6; #100;
A = 16'h0043; B = 16'h00E7; #100;
A = 16'h0043; B = 16'h00E8; #100;
A = 16'h0043; B = 16'h00E9; #100;
A = 16'h0043; B = 16'h00EA; #100;
A = 16'h0043; B = 16'h00EB; #100;
A = 16'h0043; B = 16'h00EC; #100;
A = 16'h0043; B = 16'h00ED; #100;
A = 16'h0043; B = 16'h00EE; #100;
A = 16'h0043; B = 16'h00EF; #100;
A = 16'h0043; B = 16'h00F0; #100;
A = 16'h0043; B = 16'h00F1; #100;
A = 16'h0043; B = 16'h00F2; #100;
A = 16'h0043; B = 16'h00F3; #100;
A = 16'h0043; B = 16'h00F4; #100;
A = 16'h0043; B = 16'h00F5; #100;
A = 16'h0043; B = 16'h00F6; #100;
A = 16'h0043; B = 16'h00F7; #100;
A = 16'h0043; B = 16'h00F8; #100;
A = 16'h0043; B = 16'h00F9; #100;
A = 16'h0043; B = 16'h00FA; #100;
A = 16'h0043; B = 16'h00FB; #100;
A = 16'h0043; B = 16'h00FC; #100;
A = 16'h0043; B = 16'h00FD; #100;
A = 16'h0043; B = 16'h00FE; #100;
A = 16'h0043; B = 16'h00FF; #100;
A = 16'h0044; B = 16'h000; #100;
A = 16'h0044; B = 16'h001; #100;
A = 16'h0044; B = 16'h002; #100;
A = 16'h0044; B = 16'h003; #100;
A = 16'h0044; B = 16'h004; #100;
A = 16'h0044; B = 16'h005; #100;
A = 16'h0044; B = 16'h006; #100;
A = 16'h0044; B = 16'h007; #100;
A = 16'h0044; B = 16'h008; #100;
A = 16'h0044; B = 16'h009; #100;
A = 16'h0044; B = 16'h00A; #100;
A = 16'h0044; B = 16'h00B; #100;
A = 16'h0044; B = 16'h00C; #100;
A = 16'h0044; B = 16'h00D; #100;
A = 16'h0044; B = 16'h00E; #100;
A = 16'h0044; B = 16'h00F; #100;
A = 16'h0044; B = 16'h0010; #100;
A = 16'h0044; B = 16'h0011; #100;
A = 16'h0044; B = 16'h0012; #100;
A = 16'h0044; B = 16'h0013; #100;
A = 16'h0044; B = 16'h0014; #100;
A = 16'h0044; B = 16'h0015; #100;
A = 16'h0044; B = 16'h0016; #100;
A = 16'h0044; B = 16'h0017; #100;
A = 16'h0044; B = 16'h0018; #100;
A = 16'h0044; B = 16'h0019; #100;
A = 16'h0044; B = 16'h001A; #100;
A = 16'h0044; B = 16'h001B; #100;
A = 16'h0044; B = 16'h001C; #100;
A = 16'h0044; B = 16'h001D; #100;
A = 16'h0044; B = 16'h001E; #100;
A = 16'h0044; B = 16'h001F; #100;
A = 16'h0044; B = 16'h0020; #100;
A = 16'h0044; B = 16'h0021; #100;
A = 16'h0044; B = 16'h0022; #100;
A = 16'h0044; B = 16'h0023; #100;
A = 16'h0044; B = 16'h0024; #100;
A = 16'h0044; B = 16'h0025; #100;
A = 16'h0044; B = 16'h0026; #100;
A = 16'h0044; B = 16'h0027; #100;
A = 16'h0044; B = 16'h0028; #100;
A = 16'h0044; B = 16'h0029; #100;
A = 16'h0044; B = 16'h002A; #100;
A = 16'h0044; B = 16'h002B; #100;
A = 16'h0044; B = 16'h002C; #100;
A = 16'h0044; B = 16'h002D; #100;
A = 16'h0044; B = 16'h002E; #100;
A = 16'h0044; B = 16'h002F; #100;
A = 16'h0044; B = 16'h0030; #100;
A = 16'h0044; B = 16'h0031; #100;
A = 16'h0044; B = 16'h0032; #100;
A = 16'h0044; B = 16'h0033; #100;
A = 16'h0044; B = 16'h0034; #100;
A = 16'h0044; B = 16'h0035; #100;
A = 16'h0044; B = 16'h0036; #100;
A = 16'h0044; B = 16'h0037; #100;
A = 16'h0044; B = 16'h0038; #100;
A = 16'h0044; B = 16'h0039; #100;
A = 16'h0044; B = 16'h003A; #100;
A = 16'h0044; B = 16'h003B; #100;
A = 16'h0044; B = 16'h003C; #100;
A = 16'h0044; B = 16'h003D; #100;
A = 16'h0044; B = 16'h003E; #100;
A = 16'h0044; B = 16'h003F; #100;
A = 16'h0044; B = 16'h0040; #100;
A = 16'h0044; B = 16'h0041; #100;
A = 16'h0044; B = 16'h0042; #100;
A = 16'h0044; B = 16'h0043; #100;
A = 16'h0044; B = 16'h0044; #100;
A = 16'h0044; B = 16'h0045; #100;
A = 16'h0044; B = 16'h0046; #100;
A = 16'h0044; B = 16'h0047; #100;
A = 16'h0044; B = 16'h0048; #100;
A = 16'h0044; B = 16'h0049; #100;
A = 16'h0044; B = 16'h004A; #100;
A = 16'h0044; B = 16'h004B; #100;
A = 16'h0044; B = 16'h004C; #100;
A = 16'h0044; B = 16'h004D; #100;
A = 16'h0044; B = 16'h004E; #100;
A = 16'h0044; B = 16'h004F; #100;
A = 16'h0044; B = 16'h0050; #100;
A = 16'h0044; B = 16'h0051; #100;
A = 16'h0044; B = 16'h0052; #100;
A = 16'h0044; B = 16'h0053; #100;
A = 16'h0044; B = 16'h0054; #100;
A = 16'h0044; B = 16'h0055; #100;
A = 16'h0044; B = 16'h0056; #100;
A = 16'h0044; B = 16'h0057; #100;
A = 16'h0044; B = 16'h0058; #100;
A = 16'h0044; B = 16'h0059; #100;
A = 16'h0044; B = 16'h005A; #100;
A = 16'h0044; B = 16'h005B; #100;
A = 16'h0044; B = 16'h005C; #100;
A = 16'h0044; B = 16'h005D; #100;
A = 16'h0044; B = 16'h005E; #100;
A = 16'h0044; B = 16'h005F; #100;
A = 16'h0044; B = 16'h0060; #100;
A = 16'h0044; B = 16'h0061; #100;
A = 16'h0044; B = 16'h0062; #100;
A = 16'h0044; B = 16'h0063; #100;
A = 16'h0044; B = 16'h0064; #100;
A = 16'h0044; B = 16'h0065; #100;
A = 16'h0044; B = 16'h0066; #100;
A = 16'h0044; B = 16'h0067; #100;
A = 16'h0044; B = 16'h0068; #100;
A = 16'h0044; B = 16'h0069; #100;
A = 16'h0044; B = 16'h006A; #100;
A = 16'h0044; B = 16'h006B; #100;
A = 16'h0044; B = 16'h006C; #100;
A = 16'h0044; B = 16'h006D; #100;
A = 16'h0044; B = 16'h006E; #100;
A = 16'h0044; B = 16'h006F; #100;
A = 16'h0044; B = 16'h0070; #100;
A = 16'h0044; B = 16'h0071; #100;
A = 16'h0044; B = 16'h0072; #100;
A = 16'h0044; B = 16'h0073; #100;
A = 16'h0044; B = 16'h0074; #100;
A = 16'h0044; B = 16'h0075; #100;
A = 16'h0044; B = 16'h0076; #100;
A = 16'h0044; B = 16'h0077; #100;
A = 16'h0044; B = 16'h0078; #100;
A = 16'h0044; B = 16'h0079; #100;
A = 16'h0044; B = 16'h007A; #100;
A = 16'h0044; B = 16'h007B; #100;
A = 16'h0044; B = 16'h007C; #100;
A = 16'h0044; B = 16'h007D; #100;
A = 16'h0044; B = 16'h007E; #100;
A = 16'h0044; B = 16'h007F; #100;
A = 16'h0044; B = 16'h0080; #100;
A = 16'h0044; B = 16'h0081; #100;
A = 16'h0044; B = 16'h0082; #100;
A = 16'h0044; B = 16'h0083; #100;
A = 16'h0044; B = 16'h0084; #100;
A = 16'h0044; B = 16'h0085; #100;
A = 16'h0044; B = 16'h0086; #100;
A = 16'h0044; B = 16'h0087; #100;
A = 16'h0044; B = 16'h0088; #100;
A = 16'h0044; B = 16'h0089; #100;
A = 16'h0044; B = 16'h008A; #100;
A = 16'h0044; B = 16'h008B; #100;
A = 16'h0044; B = 16'h008C; #100;
A = 16'h0044; B = 16'h008D; #100;
A = 16'h0044; B = 16'h008E; #100;
A = 16'h0044; B = 16'h008F; #100;
A = 16'h0044; B = 16'h0090; #100;
A = 16'h0044; B = 16'h0091; #100;
A = 16'h0044; B = 16'h0092; #100;
A = 16'h0044; B = 16'h0093; #100;
A = 16'h0044; B = 16'h0094; #100;
A = 16'h0044; B = 16'h0095; #100;
A = 16'h0044; B = 16'h0096; #100;
A = 16'h0044; B = 16'h0097; #100;
A = 16'h0044; B = 16'h0098; #100;
A = 16'h0044; B = 16'h0099; #100;
A = 16'h0044; B = 16'h009A; #100;
A = 16'h0044; B = 16'h009B; #100;
A = 16'h0044; B = 16'h009C; #100;
A = 16'h0044; B = 16'h009D; #100;
A = 16'h0044; B = 16'h009E; #100;
A = 16'h0044; B = 16'h009F; #100;
A = 16'h0044; B = 16'h00A0; #100;
A = 16'h0044; B = 16'h00A1; #100;
A = 16'h0044; B = 16'h00A2; #100;
A = 16'h0044; B = 16'h00A3; #100;
A = 16'h0044; B = 16'h00A4; #100;
A = 16'h0044; B = 16'h00A5; #100;
A = 16'h0044; B = 16'h00A6; #100;
A = 16'h0044; B = 16'h00A7; #100;
A = 16'h0044; B = 16'h00A8; #100;
A = 16'h0044; B = 16'h00A9; #100;
A = 16'h0044; B = 16'h00AA; #100;
A = 16'h0044; B = 16'h00AB; #100;
A = 16'h0044; B = 16'h00AC; #100;
A = 16'h0044; B = 16'h00AD; #100;
A = 16'h0044; B = 16'h00AE; #100;
A = 16'h0044; B = 16'h00AF; #100;
A = 16'h0044; B = 16'h00B0; #100;
A = 16'h0044; B = 16'h00B1; #100;
A = 16'h0044; B = 16'h00B2; #100;
A = 16'h0044; B = 16'h00B3; #100;
A = 16'h0044; B = 16'h00B4; #100;
A = 16'h0044; B = 16'h00B5; #100;
A = 16'h0044; B = 16'h00B6; #100;
A = 16'h0044; B = 16'h00B7; #100;
A = 16'h0044; B = 16'h00B8; #100;
A = 16'h0044; B = 16'h00B9; #100;
A = 16'h0044; B = 16'h00BA; #100;
A = 16'h0044; B = 16'h00BB; #100;
A = 16'h0044; B = 16'h00BC; #100;
A = 16'h0044; B = 16'h00BD; #100;
A = 16'h0044; B = 16'h00BE; #100;
A = 16'h0044; B = 16'h00BF; #100;
A = 16'h0044; B = 16'h00C0; #100;
A = 16'h0044; B = 16'h00C1; #100;
A = 16'h0044; B = 16'h00C2; #100;
A = 16'h0044; B = 16'h00C3; #100;
A = 16'h0044; B = 16'h00C4; #100;
A = 16'h0044; B = 16'h00C5; #100;
A = 16'h0044; B = 16'h00C6; #100;
A = 16'h0044; B = 16'h00C7; #100;
A = 16'h0044; B = 16'h00C8; #100;
A = 16'h0044; B = 16'h00C9; #100;
A = 16'h0044; B = 16'h00CA; #100;
A = 16'h0044; B = 16'h00CB; #100;
A = 16'h0044; B = 16'h00CC; #100;
A = 16'h0044; B = 16'h00CD; #100;
A = 16'h0044; B = 16'h00CE; #100;
A = 16'h0044; B = 16'h00CF; #100;
A = 16'h0044; B = 16'h00D0; #100;
A = 16'h0044; B = 16'h00D1; #100;
A = 16'h0044; B = 16'h00D2; #100;
A = 16'h0044; B = 16'h00D3; #100;
A = 16'h0044; B = 16'h00D4; #100;
A = 16'h0044; B = 16'h00D5; #100;
A = 16'h0044; B = 16'h00D6; #100;
A = 16'h0044; B = 16'h00D7; #100;
A = 16'h0044; B = 16'h00D8; #100;
A = 16'h0044; B = 16'h00D9; #100;
A = 16'h0044; B = 16'h00DA; #100;
A = 16'h0044; B = 16'h00DB; #100;
A = 16'h0044; B = 16'h00DC; #100;
A = 16'h0044; B = 16'h00DD; #100;
A = 16'h0044; B = 16'h00DE; #100;
A = 16'h0044; B = 16'h00DF; #100;
A = 16'h0044; B = 16'h00E0; #100;
A = 16'h0044; B = 16'h00E1; #100;
A = 16'h0044; B = 16'h00E2; #100;
A = 16'h0044; B = 16'h00E3; #100;
A = 16'h0044; B = 16'h00E4; #100;
A = 16'h0044; B = 16'h00E5; #100;
A = 16'h0044; B = 16'h00E6; #100;
A = 16'h0044; B = 16'h00E7; #100;
A = 16'h0044; B = 16'h00E8; #100;
A = 16'h0044; B = 16'h00E9; #100;
A = 16'h0044; B = 16'h00EA; #100;
A = 16'h0044; B = 16'h00EB; #100;
A = 16'h0044; B = 16'h00EC; #100;
A = 16'h0044; B = 16'h00ED; #100;
A = 16'h0044; B = 16'h00EE; #100;
A = 16'h0044; B = 16'h00EF; #100;
A = 16'h0044; B = 16'h00F0; #100;
A = 16'h0044; B = 16'h00F1; #100;
A = 16'h0044; B = 16'h00F2; #100;
A = 16'h0044; B = 16'h00F3; #100;
A = 16'h0044; B = 16'h00F4; #100;
A = 16'h0044; B = 16'h00F5; #100;
A = 16'h0044; B = 16'h00F6; #100;
A = 16'h0044; B = 16'h00F7; #100;
A = 16'h0044; B = 16'h00F8; #100;
A = 16'h0044; B = 16'h00F9; #100;
A = 16'h0044; B = 16'h00FA; #100;
A = 16'h0044; B = 16'h00FB; #100;
A = 16'h0044; B = 16'h00FC; #100;
A = 16'h0044; B = 16'h00FD; #100;
A = 16'h0044; B = 16'h00FE; #100;
A = 16'h0044; B = 16'h00FF; #100;
A = 16'h0045; B = 16'h000; #100;
A = 16'h0045; B = 16'h001; #100;
A = 16'h0045; B = 16'h002; #100;
A = 16'h0045; B = 16'h003; #100;
A = 16'h0045; B = 16'h004; #100;
A = 16'h0045; B = 16'h005; #100;
A = 16'h0045; B = 16'h006; #100;
A = 16'h0045; B = 16'h007; #100;
A = 16'h0045; B = 16'h008; #100;
A = 16'h0045; B = 16'h009; #100;
A = 16'h0045; B = 16'h00A; #100;
A = 16'h0045; B = 16'h00B; #100;
A = 16'h0045; B = 16'h00C; #100;
A = 16'h0045; B = 16'h00D; #100;
A = 16'h0045; B = 16'h00E; #100;
A = 16'h0045; B = 16'h00F; #100;
A = 16'h0045; B = 16'h0010; #100;
A = 16'h0045; B = 16'h0011; #100;
A = 16'h0045; B = 16'h0012; #100;
A = 16'h0045; B = 16'h0013; #100;
A = 16'h0045; B = 16'h0014; #100;
A = 16'h0045; B = 16'h0015; #100;
A = 16'h0045; B = 16'h0016; #100;
A = 16'h0045; B = 16'h0017; #100;
A = 16'h0045; B = 16'h0018; #100;
A = 16'h0045; B = 16'h0019; #100;
A = 16'h0045; B = 16'h001A; #100;
A = 16'h0045; B = 16'h001B; #100;
A = 16'h0045; B = 16'h001C; #100;
A = 16'h0045; B = 16'h001D; #100;
A = 16'h0045; B = 16'h001E; #100;
A = 16'h0045; B = 16'h001F; #100;
A = 16'h0045; B = 16'h0020; #100;
A = 16'h0045; B = 16'h0021; #100;
A = 16'h0045; B = 16'h0022; #100;
A = 16'h0045; B = 16'h0023; #100;
A = 16'h0045; B = 16'h0024; #100;
A = 16'h0045; B = 16'h0025; #100;
A = 16'h0045; B = 16'h0026; #100;
A = 16'h0045; B = 16'h0027; #100;
A = 16'h0045; B = 16'h0028; #100;
A = 16'h0045; B = 16'h0029; #100;
A = 16'h0045; B = 16'h002A; #100;
A = 16'h0045; B = 16'h002B; #100;
A = 16'h0045; B = 16'h002C; #100;
A = 16'h0045; B = 16'h002D; #100;
A = 16'h0045; B = 16'h002E; #100;
A = 16'h0045; B = 16'h002F; #100;
A = 16'h0045; B = 16'h0030; #100;
A = 16'h0045; B = 16'h0031; #100;
A = 16'h0045; B = 16'h0032; #100;
A = 16'h0045; B = 16'h0033; #100;
A = 16'h0045; B = 16'h0034; #100;
A = 16'h0045; B = 16'h0035; #100;
A = 16'h0045; B = 16'h0036; #100;
A = 16'h0045; B = 16'h0037; #100;
A = 16'h0045; B = 16'h0038; #100;
A = 16'h0045; B = 16'h0039; #100;
A = 16'h0045; B = 16'h003A; #100;
A = 16'h0045; B = 16'h003B; #100;
A = 16'h0045; B = 16'h003C; #100;
A = 16'h0045; B = 16'h003D; #100;
A = 16'h0045; B = 16'h003E; #100;
A = 16'h0045; B = 16'h003F; #100;
A = 16'h0045; B = 16'h0040; #100;
A = 16'h0045; B = 16'h0041; #100;
A = 16'h0045; B = 16'h0042; #100;
A = 16'h0045; B = 16'h0043; #100;
A = 16'h0045; B = 16'h0044; #100;
A = 16'h0045; B = 16'h0045; #100;
A = 16'h0045; B = 16'h0046; #100;
A = 16'h0045; B = 16'h0047; #100;
A = 16'h0045; B = 16'h0048; #100;
A = 16'h0045; B = 16'h0049; #100;
A = 16'h0045; B = 16'h004A; #100;
A = 16'h0045; B = 16'h004B; #100;
A = 16'h0045; B = 16'h004C; #100;
A = 16'h0045; B = 16'h004D; #100;
A = 16'h0045; B = 16'h004E; #100;
A = 16'h0045; B = 16'h004F; #100;
A = 16'h0045; B = 16'h0050; #100;
A = 16'h0045; B = 16'h0051; #100;
A = 16'h0045; B = 16'h0052; #100;
A = 16'h0045; B = 16'h0053; #100;
A = 16'h0045; B = 16'h0054; #100;
A = 16'h0045; B = 16'h0055; #100;
A = 16'h0045; B = 16'h0056; #100;
A = 16'h0045; B = 16'h0057; #100;
A = 16'h0045; B = 16'h0058; #100;
A = 16'h0045; B = 16'h0059; #100;
A = 16'h0045; B = 16'h005A; #100;
A = 16'h0045; B = 16'h005B; #100;
A = 16'h0045; B = 16'h005C; #100;
A = 16'h0045; B = 16'h005D; #100;
A = 16'h0045; B = 16'h005E; #100;
A = 16'h0045; B = 16'h005F; #100;
A = 16'h0045; B = 16'h0060; #100;
A = 16'h0045; B = 16'h0061; #100;
A = 16'h0045; B = 16'h0062; #100;
A = 16'h0045; B = 16'h0063; #100;
A = 16'h0045; B = 16'h0064; #100;
A = 16'h0045; B = 16'h0065; #100;
A = 16'h0045; B = 16'h0066; #100;
A = 16'h0045; B = 16'h0067; #100;
A = 16'h0045; B = 16'h0068; #100;
A = 16'h0045; B = 16'h0069; #100;
A = 16'h0045; B = 16'h006A; #100;
A = 16'h0045; B = 16'h006B; #100;
A = 16'h0045; B = 16'h006C; #100;
A = 16'h0045; B = 16'h006D; #100;
A = 16'h0045; B = 16'h006E; #100;
A = 16'h0045; B = 16'h006F; #100;
A = 16'h0045; B = 16'h0070; #100;
A = 16'h0045; B = 16'h0071; #100;
A = 16'h0045; B = 16'h0072; #100;
A = 16'h0045; B = 16'h0073; #100;
A = 16'h0045; B = 16'h0074; #100;
A = 16'h0045; B = 16'h0075; #100;
A = 16'h0045; B = 16'h0076; #100;
A = 16'h0045; B = 16'h0077; #100;
A = 16'h0045; B = 16'h0078; #100;
A = 16'h0045; B = 16'h0079; #100;
A = 16'h0045; B = 16'h007A; #100;
A = 16'h0045; B = 16'h007B; #100;
A = 16'h0045; B = 16'h007C; #100;
A = 16'h0045; B = 16'h007D; #100;
A = 16'h0045; B = 16'h007E; #100;
A = 16'h0045; B = 16'h007F; #100;
A = 16'h0045; B = 16'h0080; #100;
A = 16'h0045; B = 16'h0081; #100;
A = 16'h0045; B = 16'h0082; #100;
A = 16'h0045; B = 16'h0083; #100;
A = 16'h0045; B = 16'h0084; #100;
A = 16'h0045; B = 16'h0085; #100;
A = 16'h0045; B = 16'h0086; #100;
A = 16'h0045; B = 16'h0087; #100;
A = 16'h0045; B = 16'h0088; #100;
A = 16'h0045; B = 16'h0089; #100;
A = 16'h0045; B = 16'h008A; #100;
A = 16'h0045; B = 16'h008B; #100;
A = 16'h0045; B = 16'h008C; #100;
A = 16'h0045; B = 16'h008D; #100;
A = 16'h0045; B = 16'h008E; #100;
A = 16'h0045; B = 16'h008F; #100;
A = 16'h0045; B = 16'h0090; #100;
A = 16'h0045; B = 16'h0091; #100;
A = 16'h0045; B = 16'h0092; #100;
A = 16'h0045; B = 16'h0093; #100;
A = 16'h0045; B = 16'h0094; #100;
A = 16'h0045; B = 16'h0095; #100;
A = 16'h0045; B = 16'h0096; #100;
A = 16'h0045; B = 16'h0097; #100;
A = 16'h0045; B = 16'h0098; #100;
A = 16'h0045; B = 16'h0099; #100;
A = 16'h0045; B = 16'h009A; #100;
A = 16'h0045; B = 16'h009B; #100;
A = 16'h0045; B = 16'h009C; #100;
A = 16'h0045; B = 16'h009D; #100;
A = 16'h0045; B = 16'h009E; #100;
A = 16'h0045; B = 16'h009F; #100;
A = 16'h0045; B = 16'h00A0; #100;
A = 16'h0045; B = 16'h00A1; #100;
A = 16'h0045; B = 16'h00A2; #100;
A = 16'h0045; B = 16'h00A3; #100;
A = 16'h0045; B = 16'h00A4; #100;
A = 16'h0045; B = 16'h00A5; #100;
A = 16'h0045; B = 16'h00A6; #100;
A = 16'h0045; B = 16'h00A7; #100;
A = 16'h0045; B = 16'h00A8; #100;
A = 16'h0045; B = 16'h00A9; #100;
A = 16'h0045; B = 16'h00AA; #100;
A = 16'h0045; B = 16'h00AB; #100;
A = 16'h0045; B = 16'h00AC; #100;
A = 16'h0045; B = 16'h00AD; #100;
A = 16'h0045; B = 16'h00AE; #100;
A = 16'h0045; B = 16'h00AF; #100;
A = 16'h0045; B = 16'h00B0; #100;
A = 16'h0045; B = 16'h00B1; #100;
A = 16'h0045; B = 16'h00B2; #100;
A = 16'h0045; B = 16'h00B3; #100;
A = 16'h0045; B = 16'h00B4; #100;
A = 16'h0045; B = 16'h00B5; #100;
A = 16'h0045; B = 16'h00B6; #100;
A = 16'h0045; B = 16'h00B7; #100;
A = 16'h0045; B = 16'h00B8; #100;
A = 16'h0045; B = 16'h00B9; #100;
A = 16'h0045; B = 16'h00BA; #100;
A = 16'h0045; B = 16'h00BB; #100;
A = 16'h0045; B = 16'h00BC; #100;
A = 16'h0045; B = 16'h00BD; #100;
A = 16'h0045; B = 16'h00BE; #100;
A = 16'h0045; B = 16'h00BF; #100;
A = 16'h0045; B = 16'h00C0; #100;
A = 16'h0045; B = 16'h00C1; #100;
A = 16'h0045; B = 16'h00C2; #100;
A = 16'h0045; B = 16'h00C3; #100;
A = 16'h0045; B = 16'h00C4; #100;
A = 16'h0045; B = 16'h00C5; #100;
A = 16'h0045; B = 16'h00C6; #100;
A = 16'h0045; B = 16'h00C7; #100;
A = 16'h0045; B = 16'h00C8; #100;
A = 16'h0045; B = 16'h00C9; #100;
A = 16'h0045; B = 16'h00CA; #100;
A = 16'h0045; B = 16'h00CB; #100;
A = 16'h0045; B = 16'h00CC; #100;
A = 16'h0045; B = 16'h00CD; #100;
A = 16'h0045; B = 16'h00CE; #100;
A = 16'h0045; B = 16'h00CF; #100;
A = 16'h0045; B = 16'h00D0; #100;
A = 16'h0045; B = 16'h00D1; #100;
A = 16'h0045; B = 16'h00D2; #100;
A = 16'h0045; B = 16'h00D3; #100;
A = 16'h0045; B = 16'h00D4; #100;
A = 16'h0045; B = 16'h00D5; #100;
A = 16'h0045; B = 16'h00D6; #100;
A = 16'h0045; B = 16'h00D7; #100;
A = 16'h0045; B = 16'h00D8; #100;
A = 16'h0045; B = 16'h00D9; #100;
A = 16'h0045; B = 16'h00DA; #100;
A = 16'h0045; B = 16'h00DB; #100;
A = 16'h0045; B = 16'h00DC; #100;
A = 16'h0045; B = 16'h00DD; #100;
A = 16'h0045; B = 16'h00DE; #100;
A = 16'h0045; B = 16'h00DF; #100;
A = 16'h0045; B = 16'h00E0; #100;
A = 16'h0045; B = 16'h00E1; #100;
A = 16'h0045; B = 16'h00E2; #100;
A = 16'h0045; B = 16'h00E3; #100;
A = 16'h0045; B = 16'h00E4; #100;
A = 16'h0045; B = 16'h00E5; #100;
A = 16'h0045; B = 16'h00E6; #100;
A = 16'h0045; B = 16'h00E7; #100;
A = 16'h0045; B = 16'h00E8; #100;
A = 16'h0045; B = 16'h00E9; #100;
A = 16'h0045; B = 16'h00EA; #100;
A = 16'h0045; B = 16'h00EB; #100;
A = 16'h0045; B = 16'h00EC; #100;
A = 16'h0045; B = 16'h00ED; #100;
A = 16'h0045; B = 16'h00EE; #100;
A = 16'h0045; B = 16'h00EF; #100;
A = 16'h0045; B = 16'h00F0; #100;
A = 16'h0045; B = 16'h00F1; #100;
A = 16'h0045; B = 16'h00F2; #100;
A = 16'h0045; B = 16'h00F3; #100;
A = 16'h0045; B = 16'h00F4; #100;
A = 16'h0045; B = 16'h00F5; #100;
A = 16'h0045; B = 16'h00F6; #100;
A = 16'h0045; B = 16'h00F7; #100;
A = 16'h0045; B = 16'h00F8; #100;
A = 16'h0045; B = 16'h00F9; #100;
A = 16'h0045; B = 16'h00FA; #100;
A = 16'h0045; B = 16'h00FB; #100;
A = 16'h0045; B = 16'h00FC; #100;
A = 16'h0045; B = 16'h00FD; #100;
A = 16'h0045; B = 16'h00FE; #100;
A = 16'h0045; B = 16'h00FF; #100;
A = 16'h0046; B = 16'h000; #100;
A = 16'h0046; B = 16'h001; #100;
A = 16'h0046; B = 16'h002; #100;
A = 16'h0046; B = 16'h003; #100;
A = 16'h0046; B = 16'h004; #100;
A = 16'h0046; B = 16'h005; #100;
A = 16'h0046; B = 16'h006; #100;
A = 16'h0046; B = 16'h007; #100;
A = 16'h0046; B = 16'h008; #100;
A = 16'h0046; B = 16'h009; #100;
A = 16'h0046; B = 16'h00A; #100;
A = 16'h0046; B = 16'h00B; #100;
A = 16'h0046; B = 16'h00C; #100;
A = 16'h0046; B = 16'h00D; #100;
A = 16'h0046; B = 16'h00E; #100;
A = 16'h0046; B = 16'h00F; #100;
A = 16'h0046; B = 16'h0010; #100;
A = 16'h0046; B = 16'h0011; #100;
A = 16'h0046; B = 16'h0012; #100;
A = 16'h0046; B = 16'h0013; #100;
A = 16'h0046; B = 16'h0014; #100;
A = 16'h0046; B = 16'h0015; #100;
A = 16'h0046; B = 16'h0016; #100;
A = 16'h0046; B = 16'h0017; #100;
A = 16'h0046; B = 16'h0018; #100;
A = 16'h0046; B = 16'h0019; #100;
A = 16'h0046; B = 16'h001A; #100;
A = 16'h0046; B = 16'h001B; #100;
A = 16'h0046; B = 16'h001C; #100;
A = 16'h0046; B = 16'h001D; #100;
A = 16'h0046; B = 16'h001E; #100;
A = 16'h0046; B = 16'h001F; #100;
A = 16'h0046; B = 16'h0020; #100;
A = 16'h0046; B = 16'h0021; #100;
A = 16'h0046; B = 16'h0022; #100;
A = 16'h0046; B = 16'h0023; #100;
A = 16'h0046; B = 16'h0024; #100;
A = 16'h0046; B = 16'h0025; #100;
A = 16'h0046; B = 16'h0026; #100;
A = 16'h0046; B = 16'h0027; #100;
A = 16'h0046; B = 16'h0028; #100;
A = 16'h0046; B = 16'h0029; #100;
A = 16'h0046; B = 16'h002A; #100;
A = 16'h0046; B = 16'h002B; #100;
A = 16'h0046; B = 16'h002C; #100;
A = 16'h0046; B = 16'h002D; #100;
A = 16'h0046; B = 16'h002E; #100;
A = 16'h0046; B = 16'h002F; #100;
A = 16'h0046; B = 16'h0030; #100;
A = 16'h0046; B = 16'h0031; #100;
A = 16'h0046; B = 16'h0032; #100;
A = 16'h0046; B = 16'h0033; #100;
A = 16'h0046; B = 16'h0034; #100;
A = 16'h0046; B = 16'h0035; #100;
A = 16'h0046; B = 16'h0036; #100;
A = 16'h0046; B = 16'h0037; #100;
A = 16'h0046; B = 16'h0038; #100;
A = 16'h0046; B = 16'h0039; #100;
A = 16'h0046; B = 16'h003A; #100;
A = 16'h0046; B = 16'h003B; #100;
A = 16'h0046; B = 16'h003C; #100;
A = 16'h0046; B = 16'h003D; #100;
A = 16'h0046; B = 16'h003E; #100;
A = 16'h0046; B = 16'h003F; #100;
A = 16'h0046; B = 16'h0040; #100;
A = 16'h0046; B = 16'h0041; #100;
A = 16'h0046; B = 16'h0042; #100;
A = 16'h0046; B = 16'h0043; #100;
A = 16'h0046; B = 16'h0044; #100;
A = 16'h0046; B = 16'h0045; #100;
A = 16'h0046; B = 16'h0046; #100;
A = 16'h0046; B = 16'h0047; #100;
A = 16'h0046; B = 16'h0048; #100;
A = 16'h0046; B = 16'h0049; #100;
A = 16'h0046; B = 16'h004A; #100;
A = 16'h0046; B = 16'h004B; #100;
A = 16'h0046; B = 16'h004C; #100;
A = 16'h0046; B = 16'h004D; #100;
A = 16'h0046; B = 16'h004E; #100;
A = 16'h0046; B = 16'h004F; #100;
A = 16'h0046; B = 16'h0050; #100;
A = 16'h0046; B = 16'h0051; #100;
A = 16'h0046; B = 16'h0052; #100;
A = 16'h0046; B = 16'h0053; #100;
A = 16'h0046; B = 16'h0054; #100;
A = 16'h0046; B = 16'h0055; #100;
A = 16'h0046; B = 16'h0056; #100;
A = 16'h0046; B = 16'h0057; #100;
A = 16'h0046; B = 16'h0058; #100;
A = 16'h0046; B = 16'h0059; #100;
A = 16'h0046; B = 16'h005A; #100;
A = 16'h0046; B = 16'h005B; #100;
A = 16'h0046; B = 16'h005C; #100;
A = 16'h0046; B = 16'h005D; #100;
A = 16'h0046; B = 16'h005E; #100;
A = 16'h0046; B = 16'h005F; #100;
A = 16'h0046; B = 16'h0060; #100;
A = 16'h0046; B = 16'h0061; #100;
A = 16'h0046; B = 16'h0062; #100;
A = 16'h0046; B = 16'h0063; #100;
A = 16'h0046; B = 16'h0064; #100;
A = 16'h0046; B = 16'h0065; #100;
A = 16'h0046; B = 16'h0066; #100;
A = 16'h0046; B = 16'h0067; #100;
A = 16'h0046; B = 16'h0068; #100;
A = 16'h0046; B = 16'h0069; #100;
A = 16'h0046; B = 16'h006A; #100;
A = 16'h0046; B = 16'h006B; #100;
A = 16'h0046; B = 16'h006C; #100;
A = 16'h0046; B = 16'h006D; #100;
A = 16'h0046; B = 16'h006E; #100;
A = 16'h0046; B = 16'h006F; #100;
A = 16'h0046; B = 16'h0070; #100;
A = 16'h0046; B = 16'h0071; #100;
A = 16'h0046; B = 16'h0072; #100;
A = 16'h0046; B = 16'h0073; #100;
A = 16'h0046; B = 16'h0074; #100;
A = 16'h0046; B = 16'h0075; #100;
A = 16'h0046; B = 16'h0076; #100;
A = 16'h0046; B = 16'h0077; #100;
A = 16'h0046; B = 16'h0078; #100;
A = 16'h0046; B = 16'h0079; #100;
A = 16'h0046; B = 16'h007A; #100;
A = 16'h0046; B = 16'h007B; #100;
A = 16'h0046; B = 16'h007C; #100;
A = 16'h0046; B = 16'h007D; #100;
A = 16'h0046; B = 16'h007E; #100;
A = 16'h0046; B = 16'h007F; #100;
A = 16'h0046; B = 16'h0080; #100;
A = 16'h0046; B = 16'h0081; #100;
A = 16'h0046; B = 16'h0082; #100;
A = 16'h0046; B = 16'h0083; #100;
A = 16'h0046; B = 16'h0084; #100;
A = 16'h0046; B = 16'h0085; #100;
A = 16'h0046; B = 16'h0086; #100;
A = 16'h0046; B = 16'h0087; #100;
A = 16'h0046; B = 16'h0088; #100;
A = 16'h0046; B = 16'h0089; #100;
A = 16'h0046; B = 16'h008A; #100;
A = 16'h0046; B = 16'h008B; #100;
A = 16'h0046; B = 16'h008C; #100;
A = 16'h0046; B = 16'h008D; #100;
A = 16'h0046; B = 16'h008E; #100;
A = 16'h0046; B = 16'h008F; #100;
A = 16'h0046; B = 16'h0090; #100;
A = 16'h0046; B = 16'h0091; #100;
A = 16'h0046; B = 16'h0092; #100;
A = 16'h0046; B = 16'h0093; #100;
A = 16'h0046; B = 16'h0094; #100;
A = 16'h0046; B = 16'h0095; #100;
A = 16'h0046; B = 16'h0096; #100;
A = 16'h0046; B = 16'h0097; #100;
A = 16'h0046; B = 16'h0098; #100;
A = 16'h0046; B = 16'h0099; #100;
A = 16'h0046; B = 16'h009A; #100;
A = 16'h0046; B = 16'h009B; #100;
A = 16'h0046; B = 16'h009C; #100;
A = 16'h0046; B = 16'h009D; #100;
A = 16'h0046; B = 16'h009E; #100;
A = 16'h0046; B = 16'h009F; #100;
A = 16'h0046; B = 16'h00A0; #100;
A = 16'h0046; B = 16'h00A1; #100;
A = 16'h0046; B = 16'h00A2; #100;
A = 16'h0046; B = 16'h00A3; #100;
A = 16'h0046; B = 16'h00A4; #100;
A = 16'h0046; B = 16'h00A5; #100;
A = 16'h0046; B = 16'h00A6; #100;
A = 16'h0046; B = 16'h00A7; #100;
A = 16'h0046; B = 16'h00A8; #100;
A = 16'h0046; B = 16'h00A9; #100;
A = 16'h0046; B = 16'h00AA; #100;
A = 16'h0046; B = 16'h00AB; #100;
A = 16'h0046; B = 16'h00AC; #100;
A = 16'h0046; B = 16'h00AD; #100;
A = 16'h0046; B = 16'h00AE; #100;
A = 16'h0046; B = 16'h00AF; #100;
A = 16'h0046; B = 16'h00B0; #100;
A = 16'h0046; B = 16'h00B1; #100;
A = 16'h0046; B = 16'h00B2; #100;
A = 16'h0046; B = 16'h00B3; #100;
A = 16'h0046; B = 16'h00B4; #100;
A = 16'h0046; B = 16'h00B5; #100;
A = 16'h0046; B = 16'h00B6; #100;
A = 16'h0046; B = 16'h00B7; #100;
A = 16'h0046; B = 16'h00B8; #100;
A = 16'h0046; B = 16'h00B9; #100;
A = 16'h0046; B = 16'h00BA; #100;
A = 16'h0046; B = 16'h00BB; #100;
A = 16'h0046; B = 16'h00BC; #100;
A = 16'h0046; B = 16'h00BD; #100;
A = 16'h0046; B = 16'h00BE; #100;
A = 16'h0046; B = 16'h00BF; #100;
A = 16'h0046; B = 16'h00C0; #100;
A = 16'h0046; B = 16'h00C1; #100;
A = 16'h0046; B = 16'h00C2; #100;
A = 16'h0046; B = 16'h00C3; #100;
A = 16'h0046; B = 16'h00C4; #100;
A = 16'h0046; B = 16'h00C5; #100;
A = 16'h0046; B = 16'h00C6; #100;
A = 16'h0046; B = 16'h00C7; #100;
A = 16'h0046; B = 16'h00C8; #100;
A = 16'h0046; B = 16'h00C9; #100;
A = 16'h0046; B = 16'h00CA; #100;
A = 16'h0046; B = 16'h00CB; #100;
A = 16'h0046; B = 16'h00CC; #100;
A = 16'h0046; B = 16'h00CD; #100;
A = 16'h0046; B = 16'h00CE; #100;
A = 16'h0046; B = 16'h00CF; #100;
A = 16'h0046; B = 16'h00D0; #100;
A = 16'h0046; B = 16'h00D1; #100;
A = 16'h0046; B = 16'h00D2; #100;
A = 16'h0046; B = 16'h00D3; #100;
A = 16'h0046; B = 16'h00D4; #100;
A = 16'h0046; B = 16'h00D5; #100;
A = 16'h0046; B = 16'h00D6; #100;
A = 16'h0046; B = 16'h00D7; #100;
A = 16'h0046; B = 16'h00D8; #100;
A = 16'h0046; B = 16'h00D9; #100;
A = 16'h0046; B = 16'h00DA; #100;
A = 16'h0046; B = 16'h00DB; #100;
A = 16'h0046; B = 16'h00DC; #100;
A = 16'h0046; B = 16'h00DD; #100;
A = 16'h0046; B = 16'h00DE; #100;
A = 16'h0046; B = 16'h00DF; #100;
A = 16'h0046; B = 16'h00E0; #100;
A = 16'h0046; B = 16'h00E1; #100;
A = 16'h0046; B = 16'h00E2; #100;
A = 16'h0046; B = 16'h00E3; #100;
A = 16'h0046; B = 16'h00E4; #100;
A = 16'h0046; B = 16'h00E5; #100;
A = 16'h0046; B = 16'h00E6; #100;
A = 16'h0046; B = 16'h00E7; #100;
A = 16'h0046; B = 16'h00E8; #100;
A = 16'h0046; B = 16'h00E9; #100;
A = 16'h0046; B = 16'h00EA; #100;
A = 16'h0046; B = 16'h00EB; #100;
A = 16'h0046; B = 16'h00EC; #100;
A = 16'h0046; B = 16'h00ED; #100;
A = 16'h0046; B = 16'h00EE; #100;
A = 16'h0046; B = 16'h00EF; #100;
A = 16'h0046; B = 16'h00F0; #100;
A = 16'h0046; B = 16'h00F1; #100;
A = 16'h0046; B = 16'h00F2; #100;
A = 16'h0046; B = 16'h00F3; #100;
A = 16'h0046; B = 16'h00F4; #100;
A = 16'h0046; B = 16'h00F5; #100;
A = 16'h0046; B = 16'h00F6; #100;
A = 16'h0046; B = 16'h00F7; #100;
A = 16'h0046; B = 16'h00F8; #100;
A = 16'h0046; B = 16'h00F9; #100;
A = 16'h0046; B = 16'h00FA; #100;
A = 16'h0046; B = 16'h00FB; #100;
A = 16'h0046; B = 16'h00FC; #100;
A = 16'h0046; B = 16'h00FD; #100;
A = 16'h0046; B = 16'h00FE; #100;
A = 16'h0046; B = 16'h00FF; #100;
A = 16'h0047; B = 16'h000; #100;
A = 16'h0047; B = 16'h001; #100;
A = 16'h0047; B = 16'h002; #100;
A = 16'h0047; B = 16'h003; #100;
A = 16'h0047; B = 16'h004; #100;
A = 16'h0047; B = 16'h005; #100;
A = 16'h0047; B = 16'h006; #100;
A = 16'h0047; B = 16'h007; #100;
A = 16'h0047; B = 16'h008; #100;
A = 16'h0047; B = 16'h009; #100;
A = 16'h0047; B = 16'h00A; #100;
A = 16'h0047; B = 16'h00B; #100;
A = 16'h0047; B = 16'h00C; #100;
A = 16'h0047; B = 16'h00D; #100;
A = 16'h0047; B = 16'h00E; #100;
A = 16'h0047; B = 16'h00F; #100;
A = 16'h0047; B = 16'h0010; #100;
A = 16'h0047; B = 16'h0011; #100;
A = 16'h0047; B = 16'h0012; #100;
A = 16'h0047; B = 16'h0013; #100;
A = 16'h0047; B = 16'h0014; #100;
A = 16'h0047; B = 16'h0015; #100;
A = 16'h0047; B = 16'h0016; #100;
A = 16'h0047; B = 16'h0017; #100;
A = 16'h0047; B = 16'h0018; #100;
A = 16'h0047; B = 16'h0019; #100;
A = 16'h0047; B = 16'h001A; #100;
A = 16'h0047; B = 16'h001B; #100;
A = 16'h0047; B = 16'h001C; #100;
A = 16'h0047; B = 16'h001D; #100;
A = 16'h0047; B = 16'h001E; #100;
A = 16'h0047; B = 16'h001F; #100;
A = 16'h0047; B = 16'h0020; #100;
A = 16'h0047; B = 16'h0021; #100;
A = 16'h0047; B = 16'h0022; #100;
A = 16'h0047; B = 16'h0023; #100;
A = 16'h0047; B = 16'h0024; #100;
A = 16'h0047; B = 16'h0025; #100;
A = 16'h0047; B = 16'h0026; #100;
A = 16'h0047; B = 16'h0027; #100;
A = 16'h0047; B = 16'h0028; #100;
A = 16'h0047; B = 16'h0029; #100;
A = 16'h0047; B = 16'h002A; #100;
A = 16'h0047; B = 16'h002B; #100;
A = 16'h0047; B = 16'h002C; #100;
A = 16'h0047; B = 16'h002D; #100;
A = 16'h0047; B = 16'h002E; #100;
A = 16'h0047; B = 16'h002F; #100;
A = 16'h0047; B = 16'h0030; #100;
A = 16'h0047; B = 16'h0031; #100;
A = 16'h0047; B = 16'h0032; #100;
A = 16'h0047; B = 16'h0033; #100;
A = 16'h0047; B = 16'h0034; #100;
A = 16'h0047; B = 16'h0035; #100;
A = 16'h0047; B = 16'h0036; #100;
A = 16'h0047; B = 16'h0037; #100;
A = 16'h0047; B = 16'h0038; #100;
A = 16'h0047; B = 16'h0039; #100;
A = 16'h0047; B = 16'h003A; #100;
A = 16'h0047; B = 16'h003B; #100;
A = 16'h0047; B = 16'h003C; #100;
A = 16'h0047; B = 16'h003D; #100;
A = 16'h0047; B = 16'h003E; #100;
A = 16'h0047; B = 16'h003F; #100;
A = 16'h0047; B = 16'h0040; #100;
A = 16'h0047; B = 16'h0041; #100;
A = 16'h0047; B = 16'h0042; #100;
A = 16'h0047; B = 16'h0043; #100;
A = 16'h0047; B = 16'h0044; #100;
A = 16'h0047; B = 16'h0045; #100;
A = 16'h0047; B = 16'h0046; #100;
A = 16'h0047; B = 16'h0047; #100;
A = 16'h0047; B = 16'h0048; #100;
A = 16'h0047; B = 16'h0049; #100;
A = 16'h0047; B = 16'h004A; #100;
A = 16'h0047; B = 16'h004B; #100;
A = 16'h0047; B = 16'h004C; #100;
A = 16'h0047; B = 16'h004D; #100;
A = 16'h0047; B = 16'h004E; #100;
A = 16'h0047; B = 16'h004F; #100;
A = 16'h0047; B = 16'h0050; #100;
A = 16'h0047; B = 16'h0051; #100;
A = 16'h0047; B = 16'h0052; #100;
A = 16'h0047; B = 16'h0053; #100;
A = 16'h0047; B = 16'h0054; #100;
A = 16'h0047; B = 16'h0055; #100;
A = 16'h0047; B = 16'h0056; #100;
A = 16'h0047; B = 16'h0057; #100;
A = 16'h0047; B = 16'h0058; #100;
A = 16'h0047; B = 16'h0059; #100;
A = 16'h0047; B = 16'h005A; #100;
A = 16'h0047; B = 16'h005B; #100;
A = 16'h0047; B = 16'h005C; #100;
A = 16'h0047; B = 16'h005D; #100;
A = 16'h0047; B = 16'h005E; #100;
A = 16'h0047; B = 16'h005F; #100;
A = 16'h0047; B = 16'h0060; #100;
A = 16'h0047; B = 16'h0061; #100;
A = 16'h0047; B = 16'h0062; #100;
A = 16'h0047; B = 16'h0063; #100;
A = 16'h0047; B = 16'h0064; #100;
A = 16'h0047; B = 16'h0065; #100;
A = 16'h0047; B = 16'h0066; #100;
A = 16'h0047; B = 16'h0067; #100;
A = 16'h0047; B = 16'h0068; #100;
A = 16'h0047; B = 16'h0069; #100;
A = 16'h0047; B = 16'h006A; #100;
A = 16'h0047; B = 16'h006B; #100;
A = 16'h0047; B = 16'h006C; #100;
A = 16'h0047; B = 16'h006D; #100;
A = 16'h0047; B = 16'h006E; #100;
A = 16'h0047; B = 16'h006F; #100;
A = 16'h0047; B = 16'h0070; #100;
A = 16'h0047; B = 16'h0071; #100;
A = 16'h0047; B = 16'h0072; #100;
A = 16'h0047; B = 16'h0073; #100;
A = 16'h0047; B = 16'h0074; #100;
A = 16'h0047; B = 16'h0075; #100;
A = 16'h0047; B = 16'h0076; #100;
A = 16'h0047; B = 16'h0077; #100;
A = 16'h0047; B = 16'h0078; #100;
A = 16'h0047; B = 16'h0079; #100;
A = 16'h0047; B = 16'h007A; #100;
A = 16'h0047; B = 16'h007B; #100;
A = 16'h0047; B = 16'h007C; #100;
A = 16'h0047; B = 16'h007D; #100;
A = 16'h0047; B = 16'h007E; #100;
A = 16'h0047; B = 16'h007F; #100;
A = 16'h0047; B = 16'h0080; #100;
A = 16'h0047; B = 16'h0081; #100;
A = 16'h0047; B = 16'h0082; #100;
A = 16'h0047; B = 16'h0083; #100;
A = 16'h0047; B = 16'h0084; #100;
A = 16'h0047; B = 16'h0085; #100;
A = 16'h0047; B = 16'h0086; #100;
A = 16'h0047; B = 16'h0087; #100;
A = 16'h0047; B = 16'h0088; #100;
A = 16'h0047; B = 16'h0089; #100;
A = 16'h0047; B = 16'h008A; #100;
A = 16'h0047; B = 16'h008B; #100;
A = 16'h0047; B = 16'h008C; #100;
A = 16'h0047; B = 16'h008D; #100;
A = 16'h0047; B = 16'h008E; #100;
A = 16'h0047; B = 16'h008F; #100;
A = 16'h0047; B = 16'h0090; #100;
A = 16'h0047; B = 16'h0091; #100;
A = 16'h0047; B = 16'h0092; #100;
A = 16'h0047; B = 16'h0093; #100;
A = 16'h0047; B = 16'h0094; #100;
A = 16'h0047; B = 16'h0095; #100;
A = 16'h0047; B = 16'h0096; #100;
A = 16'h0047; B = 16'h0097; #100;
A = 16'h0047; B = 16'h0098; #100;
A = 16'h0047; B = 16'h0099; #100;
A = 16'h0047; B = 16'h009A; #100;
A = 16'h0047; B = 16'h009B; #100;
A = 16'h0047; B = 16'h009C; #100;
A = 16'h0047; B = 16'h009D; #100;
A = 16'h0047; B = 16'h009E; #100;
A = 16'h0047; B = 16'h009F; #100;
A = 16'h0047; B = 16'h00A0; #100;
A = 16'h0047; B = 16'h00A1; #100;
A = 16'h0047; B = 16'h00A2; #100;
A = 16'h0047; B = 16'h00A3; #100;
A = 16'h0047; B = 16'h00A4; #100;
A = 16'h0047; B = 16'h00A5; #100;
A = 16'h0047; B = 16'h00A6; #100;
A = 16'h0047; B = 16'h00A7; #100;
A = 16'h0047; B = 16'h00A8; #100;
A = 16'h0047; B = 16'h00A9; #100;
A = 16'h0047; B = 16'h00AA; #100;
A = 16'h0047; B = 16'h00AB; #100;
A = 16'h0047; B = 16'h00AC; #100;
A = 16'h0047; B = 16'h00AD; #100;
A = 16'h0047; B = 16'h00AE; #100;
A = 16'h0047; B = 16'h00AF; #100;
A = 16'h0047; B = 16'h00B0; #100;
A = 16'h0047; B = 16'h00B1; #100;
A = 16'h0047; B = 16'h00B2; #100;
A = 16'h0047; B = 16'h00B3; #100;
A = 16'h0047; B = 16'h00B4; #100;
A = 16'h0047; B = 16'h00B5; #100;
A = 16'h0047; B = 16'h00B6; #100;
A = 16'h0047; B = 16'h00B7; #100;
A = 16'h0047; B = 16'h00B8; #100;
A = 16'h0047; B = 16'h00B9; #100;
A = 16'h0047; B = 16'h00BA; #100;
A = 16'h0047; B = 16'h00BB; #100;
A = 16'h0047; B = 16'h00BC; #100;
A = 16'h0047; B = 16'h00BD; #100;
A = 16'h0047; B = 16'h00BE; #100;
A = 16'h0047; B = 16'h00BF; #100;
A = 16'h0047; B = 16'h00C0; #100;
A = 16'h0047; B = 16'h00C1; #100;
A = 16'h0047; B = 16'h00C2; #100;
A = 16'h0047; B = 16'h00C3; #100;
A = 16'h0047; B = 16'h00C4; #100;
A = 16'h0047; B = 16'h00C5; #100;
A = 16'h0047; B = 16'h00C6; #100;
A = 16'h0047; B = 16'h00C7; #100;
A = 16'h0047; B = 16'h00C8; #100;
A = 16'h0047; B = 16'h00C9; #100;
A = 16'h0047; B = 16'h00CA; #100;
A = 16'h0047; B = 16'h00CB; #100;
A = 16'h0047; B = 16'h00CC; #100;
A = 16'h0047; B = 16'h00CD; #100;
A = 16'h0047; B = 16'h00CE; #100;
A = 16'h0047; B = 16'h00CF; #100;
A = 16'h0047; B = 16'h00D0; #100;
A = 16'h0047; B = 16'h00D1; #100;
A = 16'h0047; B = 16'h00D2; #100;
A = 16'h0047; B = 16'h00D3; #100;
A = 16'h0047; B = 16'h00D4; #100;
A = 16'h0047; B = 16'h00D5; #100;
A = 16'h0047; B = 16'h00D6; #100;
A = 16'h0047; B = 16'h00D7; #100;
A = 16'h0047; B = 16'h00D8; #100;
A = 16'h0047; B = 16'h00D9; #100;
A = 16'h0047; B = 16'h00DA; #100;
A = 16'h0047; B = 16'h00DB; #100;
A = 16'h0047; B = 16'h00DC; #100;
A = 16'h0047; B = 16'h00DD; #100;
A = 16'h0047; B = 16'h00DE; #100;
A = 16'h0047; B = 16'h00DF; #100;
A = 16'h0047; B = 16'h00E0; #100;
A = 16'h0047; B = 16'h00E1; #100;
A = 16'h0047; B = 16'h00E2; #100;
A = 16'h0047; B = 16'h00E3; #100;
A = 16'h0047; B = 16'h00E4; #100;
A = 16'h0047; B = 16'h00E5; #100;
A = 16'h0047; B = 16'h00E6; #100;
A = 16'h0047; B = 16'h00E7; #100;
A = 16'h0047; B = 16'h00E8; #100;
A = 16'h0047; B = 16'h00E9; #100;
A = 16'h0047; B = 16'h00EA; #100;
A = 16'h0047; B = 16'h00EB; #100;
A = 16'h0047; B = 16'h00EC; #100;
A = 16'h0047; B = 16'h00ED; #100;
A = 16'h0047; B = 16'h00EE; #100;
A = 16'h0047; B = 16'h00EF; #100;
A = 16'h0047; B = 16'h00F0; #100;
A = 16'h0047; B = 16'h00F1; #100;
A = 16'h0047; B = 16'h00F2; #100;
A = 16'h0047; B = 16'h00F3; #100;
A = 16'h0047; B = 16'h00F4; #100;
A = 16'h0047; B = 16'h00F5; #100;
A = 16'h0047; B = 16'h00F6; #100;
A = 16'h0047; B = 16'h00F7; #100;
A = 16'h0047; B = 16'h00F8; #100;
A = 16'h0047; B = 16'h00F9; #100;
A = 16'h0047; B = 16'h00FA; #100;
A = 16'h0047; B = 16'h00FB; #100;
A = 16'h0047; B = 16'h00FC; #100;
A = 16'h0047; B = 16'h00FD; #100;
A = 16'h0047; B = 16'h00FE; #100;
A = 16'h0047; B = 16'h00FF; #100;
A = 16'h0048; B = 16'h000; #100;
A = 16'h0048; B = 16'h001; #100;
A = 16'h0048; B = 16'h002; #100;
A = 16'h0048; B = 16'h003; #100;
A = 16'h0048; B = 16'h004; #100;
A = 16'h0048; B = 16'h005; #100;
A = 16'h0048; B = 16'h006; #100;
A = 16'h0048; B = 16'h007; #100;
A = 16'h0048; B = 16'h008; #100;
A = 16'h0048; B = 16'h009; #100;
A = 16'h0048; B = 16'h00A; #100;
A = 16'h0048; B = 16'h00B; #100;
A = 16'h0048; B = 16'h00C; #100;
A = 16'h0048; B = 16'h00D; #100;
A = 16'h0048; B = 16'h00E; #100;
A = 16'h0048; B = 16'h00F; #100;
A = 16'h0048; B = 16'h0010; #100;
A = 16'h0048; B = 16'h0011; #100;
A = 16'h0048; B = 16'h0012; #100;
A = 16'h0048; B = 16'h0013; #100;
A = 16'h0048; B = 16'h0014; #100;
A = 16'h0048; B = 16'h0015; #100;
A = 16'h0048; B = 16'h0016; #100;
A = 16'h0048; B = 16'h0017; #100;
A = 16'h0048; B = 16'h0018; #100;
A = 16'h0048; B = 16'h0019; #100;
A = 16'h0048; B = 16'h001A; #100;
A = 16'h0048; B = 16'h001B; #100;
A = 16'h0048; B = 16'h001C; #100;
A = 16'h0048; B = 16'h001D; #100;
A = 16'h0048; B = 16'h001E; #100;
A = 16'h0048; B = 16'h001F; #100;
A = 16'h0048; B = 16'h0020; #100;
A = 16'h0048; B = 16'h0021; #100;
A = 16'h0048; B = 16'h0022; #100;
A = 16'h0048; B = 16'h0023; #100;
A = 16'h0048; B = 16'h0024; #100;
A = 16'h0048; B = 16'h0025; #100;
A = 16'h0048; B = 16'h0026; #100;
A = 16'h0048; B = 16'h0027; #100;
A = 16'h0048; B = 16'h0028; #100;
A = 16'h0048; B = 16'h0029; #100;
A = 16'h0048; B = 16'h002A; #100;
A = 16'h0048; B = 16'h002B; #100;
A = 16'h0048; B = 16'h002C; #100;
A = 16'h0048; B = 16'h002D; #100;
A = 16'h0048; B = 16'h002E; #100;
A = 16'h0048; B = 16'h002F; #100;
A = 16'h0048; B = 16'h0030; #100;
A = 16'h0048; B = 16'h0031; #100;
A = 16'h0048; B = 16'h0032; #100;
A = 16'h0048; B = 16'h0033; #100;
A = 16'h0048; B = 16'h0034; #100;
A = 16'h0048; B = 16'h0035; #100;
A = 16'h0048; B = 16'h0036; #100;
A = 16'h0048; B = 16'h0037; #100;
A = 16'h0048; B = 16'h0038; #100;
A = 16'h0048; B = 16'h0039; #100;
A = 16'h0048; B = 16'h003A; #100;
A = 16'h0048; B = 16'h003B; #100;
A = 16'h0048; B = 16'h003C; #100;
A = 16'h0048; B = 16'h003D; #100;
A = 16'h0048; B = 16'h003E; #100;
A = 16'h0048; B = 16'h003F; #100;
A = 16'h0048; B = 16'h0040; #100;
A = 16'h0048; B = 16'h0041; #100;
A = 16'h0048; B = 16'h0042; #100;
A = 16'h0048; B = 16'h0043; #100;
A = 16'h0048; B = 16'h0044; #100;
A = 16'h0048; B = 16'h0045; #100;
A = 16'h0048; B = 16'h0046; #100;
A = 16'h0048; B = 16'h0047; #100;
A = 16'h0048; B = 16'h0048; #100;
A = 16'h0048; B = 16'h0049; #100;
A = 16'h0048; B = 16'h004A; #100;
A = 16'h0048; B = 16'h004B; #100;
A = 16'h0048; B = 16'h004C; #100;
A = 16'h0048; B = 16'h004D; #100;
A = 16'h0048; B = 16'h004E; #100;
A = 16'h0048; B = 16'h004F; #100;
A = 16'h0048; B = 16'h0050; #100;
A = 16'h0048; B = 16'h0051; #100;
A = 16'h0048; B = 16'h0052; #100;
A = 16'h0048; B = 16'h0053; #100;
A = 16'h0048; B = 16'h0054; #100;
A = 16'h0048; B = 16'h0055; #100;
A = 16'h0048; B = 16'h0056; #100;
A = 16'h0048; B = 16'h0057; #100;
A = 16'h0048; B = 16'h0058; #100;
A = 16'h0048; B = 16'h0059; #100;
A = 16'h0048; B = 16'h005A; #100;
A = 16'h0048; B = 16'h005B; #100;
A = 16'h0048; B = 16'h005C; #100;
A = 16'h0048; B = 16'h005D; #100;
A = 16'h0048; B = 16'h005E; #100;
A = 16'h0048; B = 16'h005F; #100;
A = 16'h0048; B = 16'h0060; #100;
A = 16'h0048; B = 16'h0061; #100;
A = 16'h0048; B = 16'h0062; #100;
A = 16'h0048; B = 16'h0063; #100;
A = 16'h0048; B = 16'h0064; #100;
A = 16'h0048; B = 16'h0065; #100;
A = 16'h0048; B = 16'h0066; #100;
A = 16'h0048; B = 16'h0067; #100;
A = 16'h0048; B = 16'h0068; #100;
A = 16'h0048; B = 16'h0069; #100;
A = 16'h0048; B = 16'h006A; #100;
A = 16'h0048; B = 16'h006B; #100;
A = 16'h0048; B = 16'h006C; #100;
A = 16'h0048; B = 16'h006D; #100;
A = 16'h0048; B = 16'h006E; #100;
A = 16'h0048; B = 16'h006F; #100;
A = 16'h0048; B = 16'h0070; #100;
A = 16'h0048; B = 16'h0071; #100;
A = 16'h0048; B = 16'h0072; #100;
A = 16'h0048; B = 16'h0073; #100;
A = 16'h0048; B = 16'h0074; #100;
A = 16'h0048; B = 16'h0075; #100;
A = 16'h0048; B = 16'h0076; #100;
A = 16'h0048; B = 16'h0077; #100;
A = 16'h0048; B = 16'h0078; #100;
A = 16'h0048; B = 16'h0079; #100;
A = 16'h0048; B = 16'h007A; #100;
A = 16'h0048; B = 16'h007B; #100;
A = 16'h0048; B = 16'h007C; #100;
A = 16'h0048; B = 16'h007D; #100;
A = 16'h0048; B = 16'h007E; #100;
A = 16'h0048; B = 16'h007F; #100;
A = 16'h0048; B = 16'h0080; #100;
A = 16'h0048; B = 16'h0081; #100;
A = 16'h0048; B = 16'h0082; #100;
A = 16'h0048; B = 16'h0083; #100;
A = 16'h0048; B = 16'h0084; #100;
A = 16'h0048; B = 16'h0085; #100;
A = 16'h0048; B = 16'h0086; #100;
A = 16'h0048; B = 16'h0087; #100;
A = 16'h0048; B = 16'h0088; #100;
A = 16'h0048; B = 16'h0089; #100;
A = 16'h0048; B = 16'h008A; #100;
A = 16'h0048; B = 16'h008B; #100;
A = 16'h0048; B = 16'h008C; #100;
A = 16'h0048; B = 16'h008D; #100;
A = 16'h0048; B = 16'h008E; #100;
A = 16'h0048; B = 16'h008F; #100;
A = 16'h0048; B = 16'h0090; #100;
A = 16'h0048; B = 16'h0091; #100;
A = 16'h0048; B = 16'h0092; #100;
A = 16'h0048; B = 16'h0093; #100;
A = 16'h0048; B = 16'h0094; #100;
A = 16'h0048; B = 16'h0095; #100;
A = 16'h0048; B = 16'h0096; #100;
A = 16'h0048; B = 16'h0097; #100;
A = 16'h0048; B = 16'h0098; #100;
A = 16'h0048; B = 16'h0099; #100;
A = 16'h0048; B = 16'h009A; #100;
A = 16'h0048; B = 16'h009B; #100;
A = 16'h0048; B = 16'h009C; #100;
A = 16'h0048; B = 16'h009D; #100;
A = 16'h0048; B = 16'h009E; #100;
A = 16'h0048; B = 16'h009F; #100;
A = 16'h0048; B = 16'h00A0; #100;
A = 16'h0048; B = 16'h00A1; #100;
A = 16'h0048; B = 16'h00A2; #100;
A = 16'h0048; B = 16'h00A3; #100;
A = 16'h0048; B = 16'h00A4; #100;
A = 16'h0048; B = 16'h00A5; #100;
A = 16'h0048; B = 16'h00A6; #100;
A = 16'h0048; B = 16'h00A7; #100;
A = 16'h0048; B = 16'h00A8; #100;
A = 16'h0048; B = 16'h00A9; #100;
A = 16'h0048; B = 16'h00AA; #100;
A = 16'h0048; B = 16'h00AB; #100;
A = 16'h0048; B = 16'h00AC; #100;
A = 16'h0048; B = 16'h00AD; #100;
A = 16'h0048; B = 16'h00AE; #100;
A = 16'h0048; B = 16'h00AF; #100;
A = 16'h0048; B = 16'h00B0; #100;
A = 16'h0048; B = 16'h00B1; #100;
A = 16'h0048; B = 16'h00B2; #100;
A = 16'h0048; B = 16'h00B3; #100;
A = 16'h0048; B = 16'h00B4; #100;
A = 16'h0048; B = 16'h00B5; #100;
A = 16'h0048; B = 16'h00B6; #100;
A = 16'h0048; B = 16'h00B7; #100;
A = 16'h0048; B = 16'h00B8; #100;
A = 16'h0048; B = 16'h00B9; #100;
A = 16'h0048; B = 16'h00BA; #100;
A = 16'h0048; B = 16'h00BB; #100;
A = 16'h0048; B = 16'h00BC; #100;
A = 16'h0048; B = 16'h00BD; #100;
A = 16'h0048; B = 16'h00BE; #100;
A = 16'h0048; B = 16'h00BF; #100;
A = 16'h0048; B = 16'h00C0; #100;
A = 16'h0048; B = 16'h00C1; #100;
A = 16'h0048; B = 16'h00C2; #100;
A = 16'h0048; B = 16'h00C3; #100;
A = 16'h0048; B = 16'h00C4; #100;
A = 16'h0048; B = 16'h00C5; #100;
A = 16'h0048; B = 16'h00C6; #100;
A = 16'h0048; B = 16'h00C7; #100;
A = 16'h0048; B = 16'h00C8; #100;
A = 16'h0048; B = 16'h00C9; #100;
A = 16'h0048; B = 16'h00CA; #100;
A = 16'h0048; B = 16'h00CB; #100;
A = 16'h0048; B = 16'h00CC; #100;
A = 16'h0048; B = 16'h00CD; #100;
A = 16'h0048; B = 16'h00CE; #100;
A = 16'h0048; B = 16'h00CF; #100;
A = 16'h0048; B = 16'h00D0; #100;
A = 16'h0048; B = 16'h00D1; #100;
A = 16'h0048; B = 16'h00D2; #100;
A = 16'h0048; B = 16'h00D3; #100;
A = 16'h0048; B = 16'h00D4; #100;
A = 16'h0048; B = 16'h00D5; #100;
A = 16'h0048; B = 16'h00D6; #100;
A = 16'h0048; B = 16'h00D7; #100;
A = 16'h0048; B = 16'h00D8; #100;
A = 16'h0048; B = 16'h00D9; #100;
A = 16'h0048; B = 16'h00DA; #100;
A = 16'h0048; B = 16'h00DB; #100;
A = 16'h0048; B = 16'h00DC; #100;
A = 16'h0048; B = 16'h00DD; #100;
A = 16'h0048; B = 16'h00DE; #100;
A = 16'h0048; B = 16'h00DF; #100;
A = 16'h0048; B = 16'h00E0; #100;
A = 16'h0048; B = 16'h00E1; #100;
A = 16'h0048; B = 16'h00E2; #100;
A = 16'h0048; B = 16'h00E3; #100;
A = 16'h0048; B = 16'h00E4; #100;
A = 16'h0048; B = 16'h00E5; #100;
A = 16'h0048; B = 16'h00E6; #100;
A = 16'h0048; B = 16'h00E7; #100;
A = 16'h0048; B = 16'h00E8; #100;
A = 16'h0048; B = 16'h00E9; #100;
A = 16'h0048; B = 16'h00EA; #100;
A = 16'h0048; B = 16'h00EB; #100;
A = 16'h0048; B = 16'h00EC; #100;
A = 16'h0048; B = 16'h00ED; #100;
A = 16'h0048; B = 16'h00EE; #100;
A = 16'h0048; B = 16'h00EF; #100;
A = 16'h0048; B = 16'h00F0; #100;
A = 16'h0048; B = 16'h00F1; #100;
A = 16'h0048; B = 16'h00F2; #100;
A = 16'h0048; B = 16'h00F3; #100;
A = 16'h0048; B = 16'h00F4; #100;
A = 16'h0048; B = 16'h00F5; #100;
A = 16'h0048; B = 16'h00F6; #100;
A = 16'h0048; B = 16'h00F7; #100;
A = 16'h0048; B = 16'h00F8; #100;
A = 16'h0048; B = 16'h00F9; #100;
A = 16'h0048; B = 16'h00FA; #100;
A = 16'h0048; B = 16'h00FB; #100;
A = 16'h0048; B = 16'h00FC; #100;
A = 16'h0048; B = 16'h00FD; #100;
A = 16'h0048; B = 16'h00FE; #100;
A = 16'h0048; B = 16'h00FF; #100;
A = 16'h0049; B = 16'h000; #100;
A = 16'h0049; B = 16'h001; #100;
A = 16'h0049; B = 16'h002; #100;
A = 16'h0049; B = 16'h003; #100;
A = 16'h0049; B = 16'h004; #100;
A = 16'h0049; B = 16'h005; #100;
A = 16'h0049; B = 16'h006; #100;
A = 16'h0049; B = 16'h007; #100;
A = 16'h0049; B = 16'h008; #100;
A = 16'h0049; B = 16'h009; #100;
A = 16'h0049; B = 16'h00A; #100;
A = 16'h0049; B = 16'h00B; #100;
A = 16'h0049; B = 16'h00C; #100;
A = 16'h0049; B = 16'h00D; #100;
A = 16'h0049; B = 16'h00E; #100;
A = 16'h0049; B = 16'h00F; #100;
A = 16'h0049; B = 16'h0010; #100;
A = 16'h0049; B = 16'h0011; #100;
A = 16'h0049; B = 16'h0012; #100;
A = 16'h0049; B = 16'h0013; #100;
A = 16'h0049; B = 16'h0014; #100;
A = 16'h0049; B = 16'h0015; #100;
A = 16'h0049; B = 16'h0016; #100;
A = 16'h0049; B = 16'h0017; #100;
A = 16'h0049; B = 16'h0018; #100;
A = 16'h0049; B = 16'h0019; #100;
A = 16'h0049; B = 16'h001A; #100;
A = 16'h0049; B = 16'h001B; #100;
A = 16'h0049; B = 16'h001C; #100;
A = 16'h0049; B = 16'h001D; #100;
A = 16'h0049; B = 16'h001E; #100;
A = 16'h0049; B = 16'h001F; #100;
A = 16'h0049; B = 16'h0020; #100;
A = 16'h0049; B = 16'h0021; #100;
A = 16'h0049; B = 16'h0022; #100;
A = 16'h0049; B = 16'h0023; #100;
A = 16'h0049; B = 16'h0024; #100;
A = 16'h0049; B = 16'h0025; #100;
A = 16'h0049; B = 16'h0026; #100;
A = 16'h0049; B = 16'h0027; #100;
A = 16'h0049; B = 16'h0028; #100;
A = 16'h0049; B = 16'h0029; #100;
A = 16'h0049; B = 16'h002A; #100;
A = 16'h0049; B = 16'h002B; #100;
A = 16'h0049; B = 16'h002C; #100;
A = 16'h0049; B = 16'h002D; #100;
A = 16'h0049; B = 16'h002E; #100;
A = 16'h0049; B = 16'h002F; #100;
A = 16'h0049; B = 16'h0030; #100;
A = 16'h0049; B = 16'h0031; #100;
A = 16'h0049; B = 16'h0032; #100;
A = 16'h0049; B = 16'h0033; #100;
A = 16'h0049; B = 16'h0034; #100;
A = 16'h0049; B = 16'h0035; #100;
A = 16'h0049; B = 16'h0036; #100;
A = 16'h0049; B = 16'h0037; #100;
A = 16'h0049; B = 16'h0038; #100;
A = 16'h0049; B = 16'h0039; #100;
A = 16'h0049; B = 16'h003A; #100;
A = 16'h0049; B = 16'h003B; #100;
A = 16'h0049; B = 16'h003C; #100;
A = 16'h0049; B = 16'h003D; #100;
A = 16'h0049; B = 16'h003E; #100;
A = 16'h0049; B = 16'h003F; #100;
A = 16'h0049; B = 16'h0040; #100;
A = 16'h0049; B = 16'h0041; #100;
A = 16'h0049; B = 16'h0042; #100;
A = 16'h0049; B = 16'h0043; #100;
A = 16'h0049; B = 16'h0044; #100;
A = 16'h0049; B = 16'h0045; #100;
A = 16'h0049; B = 16'h0046; #100;
A = 16'h0049; B = 16'h0047; #100;
A = 16'h0049; B = 16'h0048; #100;
A = 16'h0049; B = 16'h0049; #100;
A = 16'h0049; B = 16'h004A; #100;
A = 16'h0049; B = 16'h004B; #100;
A = 16'h0049; B = 16'h004C; #100;
A = 16'h0049; B = 16'h004D; #100;
A = 16'h0049; B = 16'h004E; #100;
A = 16'h0049; B = 16'h004F; #100;
A = 16'h0049; B = 16'h0050; #100;
A = 16'h0049; B = 16'h0051; #100;
A = 16'h0049; B = 16'h0052; #100;
A = 16'h0049; B = 16'h0053; #100;
A = 16'h0049; B = 16'h0054; #100;
A = 16'h0049; B = 16'h0055; #100;
A = 16'h0049; B = 16'h0056; #100;
A = 16'h0049; B = 16'h0057; #100;
A = 16'h0049; B = 16'h0058; #100;
A = 16'h0049; B = 16'h0059; #100;
A = 16'h0049; B = 16'h005A; #100;
A = 16'h0049; B = 16'h005B; #100;
A = 16'h0049; B = 16'h005C; #100;
A = 16'h0049; B = 16'h005D; #100;
A = 16'h0049; B = 16'h005E; #100;
A = 16'h0049; B = 16'h005F; #100;
A = 16'h0049; B = 16'h0060; #100;
A = 16'h0049; B = 16'h0061; #100;
A = 16'h0049; B = 16'h0062; #100;
A = 16'h0049; B = 16'h0063; #100;
A = 16'h0049; B = 16'h0064; #100;
A = 16'h0049; B = 16'h0065; #100;
A = 16'h0049; B = 16'h0066; #100;
A = 16'h0049; B = 16'h0067; #100;
A = 16'h0049; B = 16'h0068; #100;
A = 16'h0049; B = 16'h0069; #100;
A = 16'h0049; B = 16'h006A; #100;
A = 16'h0049; B = 16'h006B; #100;
A = 16'h0049; B = 16'h006C; #100;
A = 16'h0049; B = 16'h006D; #100;
A = 16'h0049; B = 16'h006E; #100;
A = 16'h0049; B = 16'h006F; #100;
A = 16'h0049; B = 16'h0070; #100;
A = 16'h0049; B = 16'h0071; #100;
A = 16'h0049; B = 16'h0072; #100;
A = 16'h0049; B = 16'h0073; #100;
A = 16'h0049; B = 16'h0074; #100;
A = 16'h0049; B = 16'h0075; #100;
A = 16'h0049; B = 16'h0076; #100;
A = 16'h0049; B = 16'h0077; #100;
A = 16'h0049; B = 16'h0078; #100;
A = 16'h0049; B = 16'h0079; #100;
A = 16'h0049; B = 16'h007A; #100;
A = 16'h0049; B = 16'h007B; #100;
A = 16'h0049; B = 16'h007C; #100;
A = 16'h0049; B = 16'h007D; #100;
A = 16'h0049; B = 16'h007E; #100;
A = 16'h0049; B = 16'h007F; #100;
A = 16'h0049; B = 16'h0080; #100;
A = 16'h0049; B = 16'h0081; #100;
A = 16'h0049; B = 16'h0082; #100;
A = 16'h0049; B = 16'h0083; #100;
A = 16'h0049; B = 16'h0084; #100;
A = 16'h0049; B = 16'h0085; #100;
A = 16'h0049; B = 16'h0086; #100;
A = 16'h0049; B = 16'h0087; #100;
A = 16'h0049; B = 16'h0088; #100;
A = 16'h0049; B = 16'h0089; #100;
A = 16'h0049; B = 16'h008A; #100;
A = 16'h0049; B = 16'h008B; #100;
A = 16'h0049; B = 16'h008C; #100;
A = 16'h0049; B = 16'h008D; #100;
A = 16'h0049; B = 16'h008E; #100;
A = 16'h0049; B = 16'h008F; #100;
A = 16'h0049; B = 16'h0090; #100;
A = 16'h0049; B = 16'h0091; #100;
A = 16'h0049; B = 16'h0092; #100;
A = 16'h0049; B = 16'h0093; #100;
A = 16'h0049; B = 16'h0094; #100;
A = 16'h0049; B = 16'h0095; #100;
A = 16'h0049; B = 16'h0096; #100;
A = 16'h0049; B = 16'h0097; #100;
A = 16'h0049; B = 16'h0098; #100;
A = 16'h0049; B = 16'h0099; #100;
A = 16'h0049; B = 16'h009A; #100;
A = 16'h0049; B = 16'h009B; #100;
A = 16'h0049; B = 16'h009C; #100;
A = 16'h0049; B = 16'h009D; #100;
A = 16'h0049; B = 16'h009E; #100;
A = 16'h0049; B = 16'h009F; #100;
A = 16'h0049; B = 16'h00A0; #100;
A = 16'h0049; B = 16'h00A1; #100;
A = 16'h0049; B = 16'h00A2; #100;
A = 16'h0049; B = 16'h00A3; #100;
A = 16'h0049; B = 16'h00A4; #100;
A = 16'h0049; B = 16'h00A5; #100;
A = 16'h0049; B = 16'h00A6; #100;
A = 16'h0049; B = 16'h00A7; #100;
A = 16'h0049; B = 16'h00A8; #100;
A = 16'h0049; B = 16'h00A9; #100;
A = 16'h0049; B = 16'h00AA; #100;
A = 16'h0049; B = 16'h00AB; #100;
A = 16'h0049; B = 16'h00AC; #100;
A = 16'h0049; B = 16'h00AD; #100;
A = 16'h0049; B = 16'h00AE; #100;
A = 16'h0049; B = 16'h00AF; #100;
A = 16'h0049; B = 16'h00B0; #100;
A = 16'h0049; B = 16'h00B1; #100;
A = 16'h0049; B = 16'h00B2; #100;
A = 16'h0049; B = 16'h00B3; #100;
A = 16'h0049; B = 16'h00B4; #100;
A = 16'h0049; B = 16'h00B5; #100;
A = 16'h0049; B = 16'h00B6; #100;
A = 16'h0049; B = 16'h00B7; #100;
A = 16'h0049; B = 16'h00B8; #100;
A = 16'h0049; B = 16'h00B9; #100;
A = 16'h0049; B = 16'h00BA; #100;
A = 16'h0049; B = 16'h00BB; #100;
A = 16'h0049; B = 16'h00BC; #100;
A = 16'h0049; B = 16'h00BD; #100;
A = 16'h0049; B = 16'h00BE; #100;
A = 16'h0049; B = 16'h00BF; #100;
A = 16'h0049; B = 16'h00C0; #100;
A = 16'h0049; B = 16'h00C1; #100;
A = 16'h0049; B = 16'h00C2; #100;
A = 16'h0049; B = 16'h00C3; #100;
A = 16'h0049; B = 16'h00C4; #100;
A = 16'h0049; B = 16'h00C5; #100;
A = 16'h0049; B = 16'h00C6; #100;
A = 16'h0049; B = 16'h00C7; #100;
A = 16'h0049; B = 16'h00C8; #100;
A = 16'h0049; B = 16'h00C9; #100;
A = 16'h0049; B = 16'h00CA; #100;
A = 16'h0049; B = 16'h00CB; #100;
A = 16'h0049; B = 16'h00CC; #100;
A = 16'h0049; B = 16'h00CD; #100;
A = 16'h0049; B = 16'h00CE; #100;
A = 16'h0049; B = 16'h00CF; #100;
A = 16'h0049; B = 16'h00D0; #100;
A = 16'h0049; B = 16'h00D1; #100;
A = 16'h0049; B = 16'h00D2; #100;
A = 16'h0049; B = 16'h00D3; #100;
A = 16'h0049; B = 16'h00D4; #100;
A = 16'h0049; B = 16'h00D5; #100;
A = 16'h0049; B = 16'h00D6; #100;
A = 16'h0049; B = 16'h00D7; #100;
A = 16'h0049; B = 16'h00D8; #100;
A = 16'h0049; B = 16'h00D9; #100;
A = 16'h0049; B = 16'h00DA; #100;
A = 16'h0049; B = 16'h00DB; #100;
A = 16'h0049; B = 16'h00DC; #100;
A = 16'h0049; B = 16'h00DD; #100;
A = 16'h0049; B = 16'h00DE; #100;
A = 16'h0049; B = 16'h00DF; #100;
A = 16'h0049; B = 16'h00E0; #100;
A = 16'h0049; B = 16'h00E1; #100;
A = 16'h0049; B = 16'h00E2; #100;
A = 16'h0049; B = 16'h00E3; #100;
A = 16'h0049; B = 16'h00E4; #100;
A = 16'h0049; B = 16'h00E5; #100;
A = 16'h0049; B = 16'h00E6; #100;
A = 16'h0049; B = 16'h00E7; #100;
A = 16'h0049; B = 16'h00E8; #100;
A = 16'h0049; B = 16'h00E9; #100;
A = 16'h0049; B = 16'h00EA; #100;
A = 16'h0049; B = 16'h00EB; #100;
A = 16'h0049; B = 16'h00EC; #100;
A = 16'h0049; B = 16'h00ED; #100;
A = 16'h0049; B = 16'h00EE; #100;
A = 16'h0049; B = 16'h00EF; #100;
A = 16'h0049; B = 16'h00F0; #100;
A = 16'h0049; B = 16'h00F1; #100;
A = 16'h0049; B = 16'h00F2; #100;
A = 16'h0049; B = 16'h00F3; #100;
A = 16'h0049; B = 16'h00F4; #100;
A = 16'h0049; B = 16'h00F5; #100;
A = 16'h0049; B = 16'h00F6; #100;
A = 16'h0049; B = 16'h00F7; #100;
A = 16'h0049; B = 16'h00F8; #100;
A = 16'h0049; B = 16'h00F9; #100;
A = 16'h0049; B = 16'h00FA; #100;
A = 16'h0049; B = 16'h00FB; #100;
A = 16'h0049; B = 16'h00FC; #100;
A = 16'h0049; B = 16'h00FD; #100;
A = 16'h0049; B = 16'h00FE; #100;
A = 16'h0049; B = 16'h00FF; #100;
A = 16'h004A; B = 16'h000; #100;
A = 16'h004A; B = 16'h001; #100;
A = 16'h004A; B = 16'h002; #100;
A = 16'h004A; B = 16'h003; #100;
A = 16'h004A; B = 16'h004; #100;
A = 16'h004A; B = 16'h005; #100;
A = 16'h004A; B = 16'h006; #100;
A = 16'h004A; B = 16'h007; #100;
A = 16'h004A; B = 16'h008; #100;
A = 16'h004A; B = 16'h009; #100;
A = 16'h004A; B = 16'h00A; #100;
A = 16'h004A; B = 16'h00B; #100;
A = 16'h004A; B = 16'h00C; #100;
A = 16'h004A; B = 16'h00D; #100;
A = 16'h004A; B = 16'h00E; #100;
A = 16'h004A; B = 16'h00F; #100;
A = 16'h004A; B = 16'h0010; #100;
A = 16'h004A; B = 16'h0011; #100;
A = 16'h004A; B = 16'h0012; #100;
A = 16'h004A; B = 16'h0013; #100;
A = 16'h004A; B = 16'h0014; #100;
A = 16'h004A; B = 16'h0015; #100;
A = 16'h004A; B = 16'h0016; #100;
A = 16'h004A; B = 16'h0017; #100;
A = 16'h004A; B = 16'h0018; #100;
A = 16'h004A; B = 16'h0019; #100;
A = 16'h004A; B = 16'h001A; #100;
A = 16'h004A; B = 16'h001B; #100;
A = 16'h004A; B = 16'h001C; #100;
A = 16'h004A; B = 16'h001D; #100;
A = 16'h004A; B = 16'h001E; #100;
A = 16'h004A; B = 16'h001F; #100;
A = 16'h004A; B = 16'h0020; #100;
A = 16'h004A; B = 16'h0021; #100;
A = 16'h004A; B = 16'h0022; #100;
A = 16'h004A; B = 16'h0023; #100;
A = 16'h004A; B = 16'h0024; #100;
A = 16'h004A; B = 16'h0025; #100;
A = 16'h004A; B = 16'h0026; #100;
A = 16'h004A; B = 16'h0027; #100;
A = 16'h004A; B = 16'h0028; #100;
A = 16'h004A; B = 16'h0029; #100;
A = 16'h004A; B = 16'h002A; #100;
A = 16'h004A; B = 16'h002B; #100;
A = 16'h004A; B = 16'h002C; #100;
A = 16'h004A; B = 16'h002D; #100;
A = 16'h004A; B = 16'h002E; #100;
A = 16'h004A; B = 16'h002F; #100;
A = 16'h004A; B = 16'h0030; #100;
A = 16'h004A; B = 16'h0031; #100;
A = 16'h004A; B = 16'h0032; #100;
A = 16'h004A; B = 16'h0033; #100;
A = 16'h004A; B = 16'h0034; #100;
A = 16'h004A; B = 16'h0035; #100;
A = 16'h004A; B = 16'h0036; #100;
A = 16'h004A; B = 16'h0037; #100;
A = 16'h004A; B = 16'h0038; #100;
A = 16'h004A; B = 16'h0039; #100;
A = 16'h004A; B = 16'h003A; #100;
A = 16'h004A; B = 16'h003B; #100;
A = 16'h004A; B = 16'h003C; #100;
A = 16'h004A; B = 16'h003D; #100;
A = 16'h004A; B = 16'h003E; #100;
A = 16'h004A; B = 16'h003F; #100;
A = 16'h004A; B = 16'h0040; #100;
A = 16'h004A; B = 16'h0041; #100;
A = 16'h004A; B = 16'h0042; #100;
A = 16'h004A; B = 16'h0043; #100;
A = 16'h004A; B = 16'h0044; #100;
A = 16'h004A; B = 16'h0045; #100;
A = 16'h004A; B = 16'h0046; #100;
A = 16'h004A; B = 16'h0047; #100;
A = 16'h004A; B = 16'h0048; #100;
A = 16'h004A; B = 16'h0049; #100;
A = 16'h004A; B = 16'h004A; #100;
A = 16'h004A; B = 16'h004B; #100;
A = 16'h004A; B = 16'h004C; #100;
A = 16'h004A; B = 16'h004D; #100;
A = 16'h004A; B = 16'h004E; #100;
A = 16'h004A; B = 16'h004F; #100;
A = 16'h004A; B = 16'h0050; #100;
A = 16'h004A; B = 16'h0051; #100;
A = 16'h004A; B = 16'h0052; #100;
A = 16'h004A; B = 16'h0053; #100;
A = 16'h004A; B = 16'h0054; #100;
A = 16'h004A; B = 16'h0055; #100;
A = 16'h004A; B = 16'h0056; #100;
A = 16'h004A; B = 16'h0057; #100;
A = 16'h004A; B = 16'h0058; #100;
A = 16'h004A; B = 16'h0059; #100;
A = 16'h004A; B = 16'h005A; #100;
A = 16'h004A; B = 16'h005B; #100;
A = 16'h004A; B = 16'h005C; #100;
A = 16'h004A; B = 16'h005D; #100;
A = 16'h004A; B = 16'h005E; #100;
A = 16'h004A; B = 16'h005F; #100;
A = 16'h004A; B = 16'h0060; #100;
A = 16'h004A; B = 16'h0061; #100;
A = 16'h004A; B = 16'h0062; #100;
A = 16'h004A; B = 16'h0063; #100;
A = 16'h004A; B = 16'h0064; #100;
A = 16'h004A; B = 16'h0065; #100;
A = 16'h004A; B = 16'h0066; #100;
A = 16'h004A; B = 16'h0067; #100;
A = 16'h004A; B = 16'h0068; #100;
A = 16'h004A; B = 16'h0069; #100;
A = 16'h004A; B = 16'h006A; #100;
A = 16'h004A; B = 16'h006B; #100;
A = 16'h004A; B = 16'h006C; #100;
A = 16'h004A; B = 16'h006D; #100;
A = 16'h004A; B = 16'h006E; #100;
A = 16'h004A; B = 16'h006F; #100;
A = 16'h004A; B = 16'h0070; #100;
A = 16'h004A; B = 16'h0071; #100;
A = 16'h004A; B = 16'h0072; #100;
A = 16'h004A; B = 16'h0073; #100;
A = 16'h004A; B = 16'h0074; #100;
A = 16'h004A; B = 16'h0075; #100;
A = 16'h004A; B = 16'h0076; #100;
A = 16'h004A; B = 16'h0077; #100;
A = 16'h004A; B = 16'h0078; #100;
A = 16'h004A; B = 16'h0079; #100;
A = 16'h004A; B = 16'h007A; #100;
A = 16'h004A; B = 16'h007B; #100;
A = 16'h004A; B = 16'h007C; #100;
A = 16'h004A; B = 16'h007D; #100;
A = 16'h004A; B = 16'h007E; #100;
A = 16'h004A; B = 16'h007F; #100;
A = 16'h004A; B = 16'h0080; #100;
A = 16'h004A; B = 16'h0081; #100;
A = 16'h004A; B = 16'h0082; #100;
A = 16'h004A; B = 16'h0083; #100;
A = 16'h004A; B = 16'h0084; #100;
A = 16'h004A; B = 16'h0085; #100;
A = 16'h004A; B = 16'h0086; #100;
A = 16'h004A; B = 16'h0087; #100;
A = 16'h004A; B = 16'h0088; #100;
A = 16'h004A; B = 16'h0089; #100;
A = 16'h004A; B = 16'h008A; #100;
A = 16'h004A; B = 16'h008B; #100;
A = 16'h004A; B = 16'h008C; #100;
A = 16'h004A; B = 16'h008D; #100;
A = 16'h004A; B = 16'h008E; #100;
A = 16'h004A; B = 16'h008F; #100;
A = 16'h004A; B = 16'h0090; #100;
A = 16'h004A; B = 16'h0091; #100;
A = 16'h004A; B = 16'h0092; #100;
A = 16'h004A; B = 16'h0093; #100;
A = 16'h004A; B = 16'h0094; #100;
A = 16'h004A; B = 16'h0095; #100;
A = 16'h004A; B = 16'h0096; #100;
A = 16'h004A; B = 16'h0097; #100;
A = 16'h004A; B = 16'h0098; #100;
A = 16'h004A; B = 16'h0099; #100;
A = 16'h004A; B = 16'h009A; #100;
A = 16'h004A; B = 16'h009B; #100;
A = 16'h004A; B = 16'h009C; #100;
A = 16'h004A; B = 16'h009D; #100;
A = 16'h004A; B = 16'h009E; #100;
A = 16'h004A; B = 16'h009F; #100;
A = 16'h004A; B = 16'h00A0; #100;
A = 16'h004A; B = 16'h00A1; #100;
A = 16'h004A; B = 16'h00A2; #100;
A = 16'h004A; B = 16'h00A3; #100;
A = 16'h004A; B = 16'h00A4; #100;
A = 16'h004A; B = 16'h00A5; #100;
A = 16'h004A; B = 16'h00A6; #100;
A = 16'h004A; B = 16'h00A7; #100;
A = 16'h004A; B = 16'h00A8; #100;
A = 16'h004A; B = 16'h00A9; #100;
A = 16'h004A; B = 16'h00AA; #100;
A = 16'h004A; B = 16'h00AB; #100;
A = 16'h004A; B = 16'h00AC; #100;
A = 16'h004A; B = 16'h00AD; #100;
A = 16'h004A; B = 16'h00AE; #100;
A = 16'h004A; B = 16'h00AF; #100;
A = 16'h004A; B = 16'h00B0; #100;
A = 16'h004A; B = 16'h00B1; #100;
A = 16'h004A; B = 16'h00B2; #100;
A = 16'h004A; B = 16'h00B3; #100;
A = 16'h004A; B = 16'h00B4; #100;
A = 16'h004A; B = 16'h00B5; #100;
A = 16'h004A; B = 16'h00B6; #100;
A = 16'h004A; B = 16'h00B7; #100;
A = 16'h004A; B = 16'h00B8; #100;
A = 16'h004A; B = 16'h00B9; #100;
A = 16'h004A; B = 16'h00BA; #100;
A = 16'h004A; B = 16'h00BB; #100;
A = 16'h004A; B = 16'h00BC; #100;
A = 16'h004A; B = 16'h00BD; #100;
A = 16'h004A; B = 16'h00BE; #100;
A = 16'h004A; B = 16'h00BF; #100;
A = 16'h004A; B = 16'h00C0; #100;
A = 16'h004A; B = 16'h00C1; #100;
A = 16'h004A; B = 16'h00C2; #100;
A = 16'h004A; B = 16'h00C3; #100;
A = 16'h004A; B = 16'h00C4; #100;
A = 16'h004A; B = 16'h00C5; #100;
A = 16'h004A; B = 16'h00C6; #100;
A = 16'h004A; B = 16'h00C7; #100;
A = 16'h004A; B = 16'h00C8; #100;
A = 16'h004A; B = 16'h00C9; #100;
A = 16'h004A; B = 16'h00CA; #100;
A = 16'h004A; B = 16'h00CB; #100;
A = 16'h004A; B = 16'h00CC; #100;
A = 16'h004A; B = 16'h00CD; #100;
A = 16'h004A; B = 16'h00CE; #100;
A = 16'h004A; B = 16'h00CF; #100;
A = 16'h004A; B = 16'h00D0; #100;
A = 16'h004A; B = 16'h00D1; #100;
A = 16'h004A; B = 16'h00D2; #100;
A = 16'h004A; B = 16'h00D3; #100;
A = 16'h004A; B = 16'h00D4; #100;
A = 16'h004A; B = 16'h00D5; #100;
A = 16'h004A; B = 16'h00D6; #100;
A = 16'h004A; B = 16'h00D7; #100;
A = 16'h004A; B = 16'h00D8; #100;
A = 16'h004A; B = 16'h00D9; #100;
A = 16'h004A; B = 16'h00DA; #100;
A = 16'h004A; B = 16'h00DB; #100;
A = 16'h004A; B = 16'h00DC; #100;
A = 16'h004A; B = 16'h00DD; #100;
A = 16'h004A; B = 16'h00DE; #100;
A = 16'h004A; B = 16'h00DF; #100;
A = 16'h004A; B = 16'h00E0; #100;
A = 16'h004A; B = 16'h00E1; #100;
A = 16'h004A; B = 16'h00E2; #100;
A = 16'h004A; B = 16'h00E3; #100;
A = 16'h004A; B = 16'h00E4; #100;
A = 16'h004A; B = 16'h00E5; #100;
A = 16'h004A; B = 16'h00E6; #100;
A = 16'h004A; B = 16'h00E7; #100;
A = 16'h004A; B = 16'h00E8; #100;
A = 16'h004A; B = 16'h00E9; #100;
A = 16'h004A; B = 16'h00EA; #100;
A = 16'h004A; B = 16'h00EB; #100;
A = 16'h004A; B = 16'h00EC; #100;
A = 16'h004A; B = 16'h00ED; #100;
A = 16'h004A; B = 16'h00EE; #100;
A = 16'h004A; B = 16'h00EF; #100;
A = 16'h004A; B = 16'h00F0; #100;
A = 16'h004A; B = 16'h00F1; #100;
A = 16'h004A; B = 16'h00F2; #100;
A = 16'h004A; B = 16'h00F3; #100;
A = 16'h004A; B = 16'h00F4; #100;
A = 16'h004A; B = 16'h00F5; #100;
A = 16'h004A; B = 16'h00F6; #100;
A = 16'h004A; B = 16'h00F7; #100;
A = 16'h004A; B = 16'h00F8; #100;
A = 16'h004A; B = 16'h00F9; #100;
A = 16'h004A; B = 16'h00FA; #100;
A = 16'h004A; B = 16'h00FB; #100;
A = 16'h004A; B = 16'h00FC; #100;
A = 16'h004A; B = 16'h00FD; #100;
A = 16'h004A; B = 16'h00FE; #100;
A = 16'h004A; B = 16'h00FF; #100;
A = 16'h004B; B = 16'h000; #100;
A = 16'h004B; B = 16'h001; #100;
A = 16'h004B; B = 16'h002; #100;
A = 16'h004B; B = 16'h003; #100;
A = 16'h004B; B = 16'h004; #100;
A = 16'h004B; B = 16'h005; #100;
A = 16'h004B; B = 16'h006; #100;
A = 16'h004B; B = 16'h007; #100;
A = 16'h004B; B = 16'h008; #100;
A = 16'h004B; B = 16'h009; #100;
A = 16'h004B; B = 16'h00A; #100;
A = 16'h004B; B = 16'h00B; #100;
A = 16'h004B; B = 16'h00C; #100;
A = 16'h004B; B = 16'h00D; #100;
A = 16'h004B; B = 16'h00E; #100;
A = 16'h004B; B = 16'h00F; #100;
A = 16'h004B; B = 16'h0010; #100;
A = 16'h004B; B = 16'h0011; #100;
A = 16'h004B; B = 16'h0012; #100;
A = 16'h004B; B = 16'h0013; #100;
A = 16'h004B; B = 16'h0014; #100;
A = 16'h004B; B = 16'h0015; #100;
A = 16'h004B; B = 16'h0016; #100;
A = 16'h004B; B = 16'h0017; #100;
A = 16'h004B; B = 16'h0018; #100;
A = 16'h004B; B = 16'h0019; #100;
A = 16'h004B; B = 16'h001A; #100;
A = 16'h004B; B = 16'h001B; #100;
A = 16'h004B; B = 16'h001C; #100;
A = 16'h004B; B = 16'h001D; #100;
A = 16'h004B; B = 16'h001E; #100;
A = 16'h004B; B = 16'h001F; #100;
A = 16'h004B; B = 16'h0020; #100;
A = 16'h004B; B = 16'h0021; #100;
A = 16'h004B; B = 16'h0022; #100;
A = 16'h004B; B = 16'h0023; #100;
A = 16'h004B; B = 16'h0024; #100;
A = 16'h004B; B = 16'h0025; #100;
A = 16'h004B; B = 16'h0026; #100;
A = 16'h004B; B = 16'h0027; #100;
A = 16'h004B; B = 16'h0028; #100;
A = 16'h004B; B = 16'h0029; #100;
A = 16'h004B; B = 16'h002A; #100;
A = 16'h004B; B = 16'h002B; #100;
A = 16'h004B; B = 16'h002C; #100;
A = 16'h004B; B = 16'h002D; #100;
A = 16'h004B; B = 16'h002E; #100;
A = 16'h004B; B = 16'h002F; #100;
A = 16'h004B; B = 16'h0030; #100;
A = 16'h004B; B = 16'h0031; #100;
A = 16'h004B; B = 16'h0032; #100;
A = 16'h004B; B = 16'h0033; #100;
A = 16'h004B; B = 16'h0034; #100;
A = 16'h004B; B = 16'h0035; #100;
A = 16'h004B; B = 16'h0036; #100;
A = 16'h004B; B = 16'h0037; #100;
A = 16'h004B; B = 16'h0038; #100;
A = 16'h004B; B = 16'h0039; #100;
A = 16'h004B; B = 16'h003A; #100;
A = 16'h004B; B = 16'h003B; #100;
A = 16'h004B; B = 16'h003C; #100;
A = 16'h004B; B = 16'h003D; #100;
A = 16'h004B; B = 16'h003E; #100;
A = 16'h004B; B = 16'h003F; #100;
A = 16'h004B; B = 16'h0040; #100;
A = 16'h004B; B = 16'h0041; #100;
A = 16'h004B; B = 16'h0042; #100;
A = 16'h004B; B = 16'h0043; #100;
A = 16'h004B; B = 16'h0044; #100;
A = 16'h004B; B = 16'h0045; #100;
A = 16'h004B; B = 16'h0046; #100;
A = 16'h004B; B = 16'h0047; #100;
A = 16'h004B; B = 16'h0048; #100;
A = 16'h004B; B = 16'h0049; #100;
A = 16'h004B; B = 16'h004A; #100;
A = 16'h004B; B = 16'h004B; #100;
A = 16'h004B; B = 16'h004C; #100;
A = 16'h004B; B = 16'h004D; #100;
A = 16'h004B; B = 16'h004E; #100;
A = 16'h004B; B = 16'h004F; #100;
A = 16'h004B; B = 16'h0050; #100;
A = 16'h004B; B = 16'h0051; #100;
A = 16'h004B; B = 16'h0052; #100;
A = 16'h004B; B = 16'h0053; #100;
A = 16'h004B; B = 16'h0054; #100;
A = 16'h004B; B = 16'h0055; #100;
A = 16'h004B; B = 16'h0056; #100;
A = 16'h004B; B = 16'h0057; #100;
A = 16'h004B; B = 16'h0058; #100;
A = 16'h004B; B = 16'h0059; #100;
A = 16'h004B; B = 16'h005A; #100;
A = 16'h004B; B = 16'h005B; #100;
A = 16'h004B; B = 16'h005C; #100;
A = 16'h004B; B = 16'h005D; #100;
A = 16'h004B; B = 16'h005E; #100;
A = 16'h004B; B = 16'h005F; #100;
A = 16'h004B; B = 16'h0060; #100;
A = 16'h004B; B = 16'h0061; #100;
A = 16'h004B; B = 16'h0062; #100;
A = 16'h004B; B = 16'h0063; #100;
A = 16'h004B; B = 16'h0064; #100;
A = 16'h004B; B = 16'h0065; #100;
A = 16'h004B; B = 16'h0066; #100;
A = 16'h004B; B = 16'h0067; #100;
A = 16'h004B; B = 16'h0068; #100;
A = 16'h004B; B = 16'h0069; #100;
A = 16'h004B; B = 16'h006A; #100;
A = 16'h004B; B = 16'h006B; #100;
A = 16'h004B; B = 16'h006C; #100;
A = 16'h004B; B = 16'h006D; #100;
A = 16'h004B; B = 16'h006E; #100;
A = 16'h004B; B = 16'h006F; #100;
A = 16'h004B; B = 16'h0070; #100;
A = 16'h004B; B = 16'h0071; #100;
A = 16'h004B; B = 16'h0072; #100;
A = 16'h004B; B = 16'h0073; #100;
A = 16'h004B; B = 16'h0074; #100;
A = 16'h004B; B = 16'h0075; #100;
A = 16'h004B; B = 16'h0076; #100;
A = 16'h004B; B = 16'h0077; #100;
A = 16'h004B; B = 16'h0078; #100;
A = 16'h004B; B = 16'h0079; #100;
A = 16'h004B; B = 16'h007A; #100;
A = 16'h004B; B = 16'h007B; #100;
A = 16'h004B; B = 16'h007C; #100;
A = 16'h004B; B = 16'h007D; #100;
A = 16'h004B; B = 16'h007E; #100;
A = 16'h004B; B = 16'h007F; #100;
A = 16'h004B; B = 16'h0080; #100;
A = 16'h004B; B = 16'h0081; #100;
A = 16'h004B; B = 16'h0082; #100;
A = 16'h004B; B = 16'h0083; #100;
A = 16'h004B; B = 16'h0084; #100;
A = 16'h004B; B = 16'h0085; #100;
A = 16'h004B; B = 16'h0086; #100;
A = 16'h004B; B = 16'h0087; #100;
A = 16'h004B; B = 16'h0088; #100;
A = 16'h004B; B = 16'h0089; #100;
A = 16'h004B; B = 16'h008A; #100;
A = 16'h004B; B = 16'h008B; #100;
A = 16'h004B; B = 16'h008C; #100;
A = 16'h004B; B = 16'h008D; #100;
A = 16'h004B; B = 16'h008E; #100;
A = 16'h004B; B = 16'h008F; #100;
A = 16'h004B; B = 16'h0090; #100;
A = 16'h004B; B = 16'h0091; #100;
A = 16'h004B; B = 16'h0092; #100;
A = 16'h004B; B = 16'h0093; #100;
A = 16'h004B; B = 16'h0094; #100;
A = 16'h004B; B = 16'h0095; #100;
A = 16'h004B; B = 16'h0096; #100;
A = 16'h004B; B = 16'h0097; #100;
A = 16'h004B; B = 16'h0098; #100;
A = 16'h004B; B = 16'h0099; #100;
A = 16'h004B; B = 16'h009A; #100;
A = 16'h004B; B = 16'h009B; #100;
A = 16'h004B; B = 16'h009C; #100;
A = 16'h004B; B = 16'h009D; #100;
A = 16'h004B; B = 16'h009E; #100;
A = 16'h004B; B = 16'h009F; #100;
A = 16'h004B; B = 16'h00A0; #100;
A = 16'h004B; B = 16'h00A1; #100;
A = 16'h004B; B = 16'h00A2; #100;
A = 16'h004B; B = 16'h00A3; #100;
A = 16'h004B; B = 16'h00A4; #100;
A = 16'h004B; B = 16'h00A5; #100;
A = 16'h004B; B = 16'h00A6; #100;
A = 16'h004B; B = 16'h00A7; #100;
A = 16'h004B; B = 16'h00A8; #100;
A = 16'h004B; B = 16'h00A9; #100;
A = 16'h004B; B = 16'h00AA; #100;
A = 16'h004B; B = 16'h00AB; #100;
A = 16'h004B; B = 16'h00AC; #100;
A = 16'h004B; B = 16'h00AD; #100;
A = 16'h004B; B = 16'h00AE; #100;
A = 16'h004B; B = 16'h00AF; #100;
A = 16'h004B; B = 16'h00B0; #100;
A = 16'h004B; B = 16'h00B1; #100;
A = 16'h004B; B = 16'h00B2; #100;
A = 16'h004B; B = 16'h00B3; #100;
A = 16'h004B; B = 16'h00B4; #100;
A = 16'h004B; B = 16'h00B5; #100;
A = 16'h004B; B = 16'h00B6; #100;
A = 16'h004B; B = 16'h00B7; #100;
A = 16'h004B; B = 16'h00B8; #100;
A = 16'h004B; B = 16'h00B9; #100;
A = 16'h004B; B = 16'h00BA; #100;
A = 16'h004B; B = 16'h00BB; #100;
A = 16'h004B; B = 16'h00BC; #100;
A = 16'h004B; B = 16'h00BD; #100;
A = 16'h004B; B = 16'h00BE; #100;
A = 16'h004B; B = 16'h00BF; #100;
A = 16'h004B; B = 16'h00C0; #100;
A = 16'h004B; B = 16'h00C1; #100;
A = 16'h004B; B = 16'h00C2; #100;
A = 16'h004B; B = 16'h00C3; #100;
A = 16'h004B; B = 16'h00C4; #100;
A = 16'h004B; B = 16'h00C5; #100;
A = 16'h004B; B = 16'h00C6; #100;
A = 16'h004B; B = 16'h00C7; #100;
A = 16'h004B; B = 16'h00C8; #100;
A = 16'h004B; B = 16'h00C9; #100;
A = 16'h004B; B = 16'h00CA; #100;
A = 16'h004B; B = 16'h00CB; #100;
A = 16'h004B; B = 16'h00CC; #100;
A = 16'h004B; B = 16'h00CD; #100;
A = 16'h004B; B = 16'h00CE; #100;
A = 16'h004B; B = 16'h00CF; #100;
A = 16'h004B; B = 16'h00D0; #100;
A = 16'h004B; B = 16'h00D1; #100;
A = 16'h004B; B = 16'h00D2; #100;
A = 16'h004B; B = 16'h00D3; #100;
A = 16'h004B; B = 16'h00D4; #100;
A = 16'h004B; B = 16'h00D5; #100;
A = 16'h004B; B = 16'h00D6; #100;
A = 16'h004B; B = 16'h00D7; #100;
A = 16'h004B; B = 16'h00D8; #100;
A = 16'h004B; B = 16'h00D9; #100;
A = 16'h004B; B = 16'h00DA; #100;
A = 16'h004B; B = 16'h00DB; #100;
A = 16'h004B; B = 16'h00DC; #100;
A = 16'h004B; B = 16'h00DD; #100;
A = 16'h004B; B = 16'h00DE; #100;
A = 16'h004B; B = 16'h00DF; #100;
A = 16'h004B; B = 16'h00E0; #100;
A = 16'h004B; B = 16'h00E1; #100;
A = 16'h004B; B = 16'h00E2; #100;
A = 16'h004B; B = 16'h00E3; #100;
A = 16'h004B; B = 16'h00E4; #100;
A = 16'h004B; B = 16'h00E5; #100;
A = 16'h004B; B = 16'h00E6; #100;
A = 16'h004B; B = 16'h00E7; #100;
A = 16'h004B; B = 16'h00E8; #100;
A = 16'h004B; B = 16'h00E9; #100;
A = 16'h004B; B = 16'h00EA; #100;
A = 16'h004B; B = 16'h00EB; #100;
A = 16'h004B; B = 16'h00EC; #100;
A = 16'h004B; B = 16'h00ED; #100;
A = 16'h004B; B = 16'h00EE; #100;
A = 16'h004B; B = 16'h00EF; #100;
A = 16'h004B; B = 16'h00F0; #100;
A = 16'h004B; B = 16'h00F1; #100;
A = 16'h004B; B = 16'h00F2; #100;
A = 16'h004B; B = 16'h00F3; #100;
A = 16'h004B; B = 16'h00F4; #100;
A = 16'h004B; B = 16'h00F5; #100;
A = 16'h004B; B = 16'h00F6; #100;
A = 16'h004B; B = 16'h00F7; #100;
A = 16'h004B; B = 16'h00F8; #100;
A = 16'h004B; B = 16'h00F9; #100;
A = 16'h004B; B = 16'h00FA; #100;
A = 16'h004B; B = 16'h00FB; #100;
A = 16'h004B; B = 16'h00FC; #100;
A = 16'h004B; B = 16'h00FD; #100;
A = 16'h004B; B = 16'h00FE; #100;
A = 16'h004B; B = 16'h00FF; #100;
A = 16'h004C; B = 16'h000; #100;
A = 16'h004C; B = 16'h001; #100;
A = 16'h004C; B = 16'h002; #100;
A = 16'h004C; B = 16'h003; #100;
A = 16'h004C; B = 16'h004; #100;
A = 16'h004C; B = 16'h005; #100;
A = 16'h004C; B = 16'h006; #100;
A = 16'h004C; B = 16'h007; #100;
A = 16'h004C; B = 16'h008; #100;
A = 16'h004C; B = 16'h009; #100;
A = 16'h004C; B = 16'h00A; #100;
A = 16'h004C; B = 16'h00B; #100;
A = 16'h004C; B = 16'h00C; #100;
A = 16'h004C; B = 16'h00D; #100;
A = 16'h004C; B = 16'h00E; #100;
A = 16'h004C; B = 16'h00F; #100;
A = 16'h004C; B = 16'h0010; #100;
A = 16'h004C; B = 16'h0011; #100;
A = 16'h004C; B = 16'h0012; #100;
A = 16'h004C; B = 16'h0013; #100;
A = 16'h004C; B = 16'h0014; #100;
A = 16'h004C; B = 16'h0015; #100;
A = 16'h004C; B = 16'h0016; #100;
A = 16'h004C; B = 16'h0017; #100;
A = 16'h004C; B = 16'h0018; #100;
A = 16'h004C; B = 16'h0019; #100;
A = 16'h004C; B = 16'h001A; #100;
A = 16'h004C; B = 16'h001B; #100;
A = 16'h004C; B = 16'h001C; #100;
A = 16'h004C; B = 16'h001D; #100;
A = 16'h004C; B = 16'h001E; #100;
A = 16'h004C; B = 16'h001F; #100;
A = 16'h004C; B = 16'h0020; #100;
A = 16'h004C; B = 16'h0021; #100;
A = 16'h004C; B = 16'h0022; #100;
A = 16'h004C; B = 16'h0023; #100;
A = 16'h004C; B = 16'h0024; #100;
A = 16'h004C; B = 16'h0025; #100;
A = 16'h004C; B = 16'h0026; #100;
A = 16'h004C; B = 16'h0027; #100;
A = 16'h004C; B = 16'h0028; #100;
A = 16'h004C; B = 16'h0029; #100;
A = 16'h004C; B = 16'h002A; #100;
A = 16'h004C; B = 16'h002B; #100;
A = 16'h004C; B = 16'h002C; #100;
A = 16'h004C; B = 16'h002D; #100;
A = 16'h004C; B = 16'h002E; #100;
A = 16'h004C; B = 16'h002F; #100;
A = 16'h004C; B = 16'h0030; #100;
A = 16'h004C; B = 16'h0031; #100;
A = 16'h004C; B = 16'h0032; #100;
A = 16'h004C; B = 16'h0033; #100;
A = 16'h004C; B = 16'h0034; #100;
A = 16'h004C; B = 16'h0035; #100;
A = 16'h004C; B = 16'h0036; #100;
A = 16'h004C; B = 16'h0037; #100;
A = 16'h004C; B = 16'h0038; #100;
A = 16'h004C; B = 16'h0039; #100;
A = 16'h004C; B = 16'h003A; #100;
A = 16'h004C; B = 16'h003B; #100;
A = 16'h004C; B = 16'h003C; #100;
A = 16'h004C; B = 16'h003D; #100;
A = 16'h004C; B = 16'h003E; #100;
A = 16'h004C; B = 16'h003F; #100;
A = 16'h004C; B = 16'h0040; #100;
A = 16'h004C; B = 16'h0041; #100;
A = 16'h004C; B = 16'h0042; #100;
A = 16'h004C; B = 16'h0043; #100;
A = 16'h004C; B = 16'h0044; #100;
A = 16'h004C; B = 16'h0045; #100;
A = 16'h004C; B = 16'h0046; #100;
A = 16'h004C; B = 16'h0047; #100;
A = 16'h004C; B = 16'h0048; #100;
A = 16'h004C; B = 16'h0049; #100;
A = 16'h004C; B = 16'h004A; #100;
A = 16'h004C; B = 16'h004B; #100;
A = 16'h004C; B = 16'h004C; #100;
A = 16'h004C; B = 16'h004D; #100;
A = 16'h004C; B = 16'h004E; #100;
A = 16'h004C; B = 16'h004F; #100;
A = 16'h004C; B = 16'h0050; #100;
A = 16'h004C; B = 16'h0051; #100;
A = 16'h004C; B = 16'h0052; #100;
A = 16'h004C; B = 16'h0053; #100;
A = 16'h004C; B = 16'h0054; #100;
A = 16'h004C; B = 16'h0055; #100;
A = 16'h004C; B = 16'h0056; #100;
A = 16'h004C; B = 16'h0057; #100;
A = 16'h004C; B = 16'h0058; #100;
A = 16'h004C; B = 16'h0059; #100;
A = 16'h004C; B = 16'h005A; #100;
A = 16'h004C; B = 16'h005B; #100;
A = 16'h004C; B = 16'h005C; #100;
A = 16'h004C; B = 16'h005D; #100;
A = 16'h004C; B = 16'h005E; #100;
A = 16'h004C; B = 16'h005F; #100;
A = 16'h004C; B = 16'h0060; #100;
A = 16'h004C; B = 16'h0061; #100;
A = 16'h004C; B = 16'h0062; #100;
A = 16'h004C; B = 16'h0063; #100;
A = 16'h004C; B = 16'h0064; #100;
A = 16'h004C; B = 16'h0065; #100;
A = 16'h004C; B = 16'h0066; #100;
A = 16'h004C; B = 16'h0067; #100;
A = 16'h004C; B = 16'h0068; #100;
A = 16'h004C; B = 16'h0069; #100;
A = 16'h004C; B = 16'h006A; #100;
A = 16'h004C; B = 16'h006B; #100;
A = 16'h004C; B = 16'h006C; #100;
A = 16'h004C; B = 16'h006D; #100;
A = 16'h004C; B = 16'h006E; #100;
A = 16'h004C; B = 16'h006F; #100;
A = 16'h004C; B = 16'h0070; #100;
A = 16'h004C; B = 16'h0071; #100;
A = 16'h004C; B = 16'h0072; #100;
A = 16'h004C; B = 16'h0073; #100;
A = 16'h004C; B = 16'h0074; #100;
A = 16'h004C; B = 16'h0075; #100;
A = 16'h004C; B = 16'h0076; #100;
A = 16'h004C; B = 16'h0077; #100;
A = 16'h004C; B = 16'h0078; #100;
A = 16'h004C; B = 16'h0079; #100;
A = 16'h004C; B = 16'h007A; #100;
A = 16'h004C; B = 16'h007B; #100;
A = 16'h004C; B = 16'h007C; #100;
A = 16'h004C; B = 16'h007D; #100;
A = 16'h004C; B = 16'h007E; #100;
A = 16'h004C; B = 16'h007F; #100;
A = 16'h004C; B = 16'h0080; #100;
A = 16'h004C; B = 16'h0081; #100;
A = 16'h004C; B = 16'h0082; #100;
A = 16'h004C; B = 16'h0083; #100;
A = 16'h004C; B = 16'h0084; #100;
A = 16'h004C; B = 16'h0085; #100;
A = 16'h004C; B = 16'h0086; #100;
A = 16'h004C; B = 16'h0087; #100;
A = 16'h004C; B = 16'h0088; #100;
A = 16'h004C; B = 16'h0089; #100;
A = 16'h004C; B = 16'h008A; #100;
A = 16'h004C; B = 16'h008B; #100;
A = 16'h004C; B = 16'h008C; #100;
A = 16'h004C; B = 16'h008D; #100;
A = 16'h004C; B = 16'h008E; #100;
A = 16'h004C; B = 16'h008F; #100;
A = 16'h004C; B = 16'h0090; #100;
A = 16'h004C; B = 16'h0091; #100;
A = 16'h004C; B = 16'h0092; #100;
A = 16'h004C; B = 16'h0093; #100;
A = 16'h004C; B = 16'h0094; #100;
A = 16'h004C; B = 16'h0095; #100;
A = 16'h004C; B = 16'h0096; #100;
A = 16'h004C; B = 16'h0097; #100;
A = 16'h004C; B = 16'h0098; #100;
A = 16'h004C; B = 16'h0099; #100;
A = 16'h004C; B = 16'h009A; #100;
A = 16'h004C; B = 16'h009B; #100;
A = 16'h004C; B = 16'h009C; #100;
A = 16'h004C; B = 16'h009D; #100;
A = 16'h004C; B = 16'h009E; #100;
A = 16'h004C; B = 16'h009F; #100;
A = 16'h004C; B = 16'h00A0; #100;
A = 16'h004C; B = 16'h00A1; #100;
A = 16'h004C; B = 16'h00A2; #100;
A = 16'h004C; B = 16'h00A3; #100;
A = 16'h004C; B = 16'h00A4; #100;
A = 16'h004C; B = 16'h00A5; #100;
A = 16'h004C; B = 16'h00A6; #100;
A = 16'h004C; B = 16'h00A7; #100;
A = 16'h004C; B = 16'h00A8; #100;
A = 16'h004C; B = 16'h00A9; #100;
A = 16'h004C; B = 16'h00AA; #100;
A = 16'h004C; B = 16'h00AB; #100;
A = 16'h004C; B = 16'h00AC; #100;
A = 16'h004C; B = 16'h00AD; #100;
A = 16'h004C; B = 16'h00AE; #100;
A = 16'h004C; B = 16'h00AF; #100;
A = 16'h004C; B = 16'h00B0; #100;
A = 16'h004C; B = 16'h00B1; #100;
A = 16'h004C; B = 16'h00B2; #100;
A = 16'h004C; B = 16'h00B3; #100;
A = 16'h004C; B = 16'h00B4; #100;
A = 16'h004C; B = 16'h00B5; #100;
A = 16'h004C; B = 16'h00B6; #100;
A = 16'h004C; B = 16'h00B7; #100;
A = 16'h004C; B = 16'h00B8; #100;
A = 16'h004C; B = 16'h00B9; #100;
A = 16'h004C; B = 16'h00BA; #100;
A = 16'h004C; B = 16'h00BB; #100;
A = 16'h004C; B = 16'h00BC; #100;
A = 16'h004C; B = 16'h00BD; #100;
A = 16'h004C; B = 16'h00BE; #100;
A = 16'h004C; B = 16'h00BF; #100;
A = 16'h004C; B = 16'h00C0; #100;
A = 16'h004C; B = 16'h00C1; #100;
A = 16'h004C; B = 16'h00C2; #100;
A = 16'h004C; B = 16'h00C3; #100;
A = 16'h004C; B = 16'h00C4; #100;
A = 16'h004C; B = 16'h00C5; #100;
A = 16'h004C; B = 16'h00C6; #100;
A = 16'h004C; B = 16'h00C7; #100;
A = 16'h004C; B = 16'h00C8; #100;
A = 16'h004C; B = 16'h00C9; #100;
A = 16'h004C; B = 16'h00CA; #100;
A = 16'h004C; B = 16'h00CB; #100;
A = 16'h004C; B = 16'h00CC; #100;
A = 16'h004C; B = 16'h00CD; #100;
A = 16'h004C; B = 16'h00CE; #100;
A = 16'h004C; B = 16'h00CF; #100;
A = 16'h004C; B = 16'h00D0; #100;
A = 16'h004C; B = 16'h00D1; #100;
A = 16'h004C; B = 16'h00D2; #100;
A = 16'h004C; B = 16'h00D3; #100;
A = 16'h004C; B = 16'h00D4; #100;
A = 16'h004C; B = 16'h00D5; #100;
A = 16'h004C; B = 16'h00D6; #100;
A = 16'h004C; B = 16'h00D7; #100;
A = 16'h004C; B = 16'h00D8; #100;
A = 16'h004C; B = 16'h00D9; #100;
A = 16'h004C; B = 16'h00DA; #100;
A = 16'h004C; B = 16'h00DB; #100;
A = 16'h004C; B = 16'h00DC; #100;
A = 16'h004C; B = 16'h00DD; #100;
A = 16'h004C; B = 16'h00DE; #100;
A = 16'h004C; B = 16'h00DF; #100;
A = 16'h004C; B = 16'h00E0; #100;
A = 16'h004C; B = 16'h00E1; #100;
A = 16'h004C; B = 16'h00E2; #100;
A = 16'h004C; B = 16'h00E3; #100;
A = 16'h004C; B = 16'h00E4; #100;
A = 16'h004C; B = 16'h00E5; #100;
A = 16'h004C; B = 16'h00E6; #100;
A = 16'h004C; B = 16'h00E7; #100;
A = 16'h004C; B = 16'h00E8; #100;
A = 16'h004C; B = 16'h00E9; #100;
A = 16'h004C; B = 16'h00EA; #100;
A = 16'h004C; B = 16'h00EB; #100;
A = 16'h004C; B = 16'h00EC; #100;
A = 16'h004C; B = 16'h00ED; #100;
A = 16'h004C; B = 16'h00EE; #100;
A = 16'h004C; B = 16'h00EF; #100;
A = 16'h004C; B = 16'h00F0; #100;
A = 16'h004C; B = 16'h00F1; #100;
A = 16'h004C; B = 16'h00F2; #100;
A = 16'h004C; B = 16'h00F3; #100;
A = 16'h004C; B = 16'h00F4; #100;
A = 16'h004C; B = 16'h00F5; #100;
A = 16'h004C; B = 16'h00F6; #100;
A = 16'h004C; B = 16'h00F7; #100;
A = 16'h004C; B = 16'h00F8; #100;
A = 16'h004C; B = 16'h00F9; #100;
A = 16'h004C; B = 16'h00FA; #100;
A = 16'h004C; B = 16'h00FB; #100;
A = 16'h004C; B = 16'h00FC; #100;
A = 16'h004C; B = 16'h00FD; #100;
A = 16'h004C; B = 16'h00FE; #100;
A = 16'h004C; B = 16'h00FF; #100;
A = 16'h004D; B = 16'h000; #100;
A = 16'h004D; B = 16'h001; #100;
A = 16'h004D; B = 16'h002; #100;
A = 16'h004D; B = 16'h003; #100;
A = 16'h004D; B = 16'h004; #100;
A = 16'h004D; B = 16'h005; #100;
A = 16'h004D; B = 16'h006; #100;
A = 16'h004D; B = 16'h007; #100;
A = 16'h004D; B = 16'h008; #100;
A = 16'h004D; B = 16'h009; #100;
A = 16'h004D; B = 16'h00A; #100;
A = 16'h004D; B = 16'h00B; #100;
A = 16'h004D; B = 16'h00C; #100;
A = 16'h004D; B = 16'h00D; #100;
A = 16'h004D; B = 16'h00E; #100;
A = 16'h004D; B = 16'h00F; #100;
A = 16'h004D; B = 16'h0010; #100;
A = 16'h004D; B = 16'h0011; #100;
A = 16'h004D; B = 16'h0012; #100;
A = 16'h004D; B = 16'h0013; #100;
A = 16'h004D; B = 16'h0014; #100;
A = 16'h004D; B = 16'h0015; #100;
A = 16'h004D; B = 16'h0016; #100;
A = 16'h004D; B = 16'h0017; #100;
A = 16'h004D; B = 16'h0018; #100;
A = 16'h004D; B = 16'h0019; #100;
A = 16'h004D; B = 16'h001A; #100;
A = 16'h004D; B = 16'h001B; #100;
A = 16'h004D; B = 16'h001C; #100;
A = 16'h004D; B = 16'h001D; #100;
A = 16'h004D; B = 16'h001E; #100;
A = 16'h004D; B = 16'h001F; #100;
A = 16'h004D; B = 16'h0020; #100;
A = 16'h004D; B = 16'h0021; #100;
A = 16'h004D; B = 16'h0022; #100;
A = 16'h004D; B = 16'h0023; #100;
A = 16'h004D; B = 16'h0024; #100;
A = 16'h004D; B = 16'h0025; #100;
A = 16'h004D; B = 16'h0026; #100;
A = 16'h004D; B = 16'h0027; #100;
A = 16'h004D; B = 16'h0028; #100;
A = 16'h004D; B = 16'h0029; #100;
A = 16'h004D; B = 16'h002A; #100;
A = 16'h004D; B = 16'h002B; #100;
A = 16'h004D; B = 16'h002C; #100;
A = 16'h004D; B = 16'h002D; #100;
A = 16'h004D; B = 16'h002E; #100;
A = 16'h004D; B = 16'h002F; #100;
A = 16'h004D; B = 16'h0030; #100;
A = 16'h004D; B = 16'h0031; #100;
A = 16'h004D; B = 16'h0032; #100;
A = 16'h004D; B = 16'h0033; #100;
A = 16'h004D; B = 16'h0034; #100;
A = 16'h004D; B = 16'h0035; #100;
A = 16'h004D; B = 16'h0036; #100;
A = 16'h004D; B = 16'h0037; #100;
A = 16'h004D; B = 16'h0038; #100;
A = 16'h004D; B = 16'h0039; #100;
A = 16'h004D; B = 16'h003A; #100;
A = 16'h004D; B = 16'h003B; #100;
A = 16'h004D; B = 16'h003C; #100;
A = 16'h004D; B = 16'h003D; #100;
A = 16'h004D; B = 16'h003E; #100;
A = 16'h004D; B = 16'h003F; #100;
A = 16'h004D; B = 16'h0040; #100;
A = 16'h004D; B = 16'h0041; #100;
A = 16'h004D; B = 16'h0042; #100;
A = 16'h004D; B = 16'h0043; #100;
A = 16'h004D; B = 16'h0044; #100;
A = 16'h004D; B = 16'h0045; #100;
A = 16'h004D; B = 16'h0046; #100;
A = 16'h004D; B = 16'h0047; #100;
A = 16'h004D; B = 16'h0048; #100;
A = 16'h004D; B = 16'h0049; #100;
A = 16'h004D; B = 16'h004A; #100;
A = 16'h004D; B = 16'h004B; #100;
A = 16'h004D; B = 16'h004C; #100;
A = 16'h004D; B = 16'h004D; #100;
A = 16'h004D; B = 16'h004E; #100;
A = 16'h004D; B = 16'h004F; #100;
A = 16'h004D; B = 16'h0050; #100;
A = 16'h004D; B = 16'h0051; #100;
A = 16'h004D; B = 16'h0052; #100;
A = 16'h004D; B = 16'h0053; #100;
A = 16'h004D; B = 16'h0054; #100;
A = 16'h004D; B = 16'h0055; #100;
A = 16'h004D; B = 16'h0056; #100;
A = 16'h004D; B = 16'h0057; #100;
A = 16'h004D; B = 16'h0058; #100;
A = 16'h004D; B = 16'h0059; #100;
A = 16'h004D; B = 16'h005A; #100;
A = 16'h004D; B = 16'h005B; #100;
A = 16'h004D; B = 16'h005C; #100;
A = 16'h004D; B = 16'h005D; #100;
A = 16'h004D; B = 16'h005E; #100;
A = 16'h004D; B = 16'h005F; #100;
A = 16'h004D; B = 16'h0060; #100;
A = 16'h004D; B = 16'h0061; #100;
A = 16'h004D; B = 16'h0062; #100;
A = 16'h004D; B = 16'h0063; #100;
A = 16'h004D; B = 16'h0064; #100;
A = 16'h004D; B = 16'h0065; #100;
A = 16'h004D; B = 16'h0066; #100;
A = 16'h004D; B = 16'h0067; #100;
A = 16'h004D; B = 16'h0068; #100;
A = 16'h004D; B = 16'h0069; #100;
A = 16'h004D; B = 16'h006A; #100;
A = 16'h004D; B = 16'h006B; #100;
A = 16'h004D; B = 16'h006C; #100;
A = 16'h004D; B = 16'h006D; #100;
A = 16'h004D; B = 16'h006E; #100;
A = 16'h004D; B = 16'h006F; #100;
A = 16'h004D; B = 16'h0070; #100;
A = 16'h004D; B = 16'h0071; #100;
A = 16'h004D; B = 16'h0072; #100;
A = 16'h004D; B = 16'h0073; #100;
A = 16'h004D; B = 16'h0074; #100;
A = 16'h004D; B = 16'h0075; #100;
A = 16'h004D; B = 16'h0076; #100;
A = 16'h004D; B = 16'h0077; #100;
A = 16'h004D; B = 16'h0078; #100;
A = 16'h004D; B = 16'h0079; #100;
A = 16'h004D; B = 16'h007A; #100;
A = 16'h004D; B = 16'h007B; #100;
A = 16'h004D; B = 16'h007C; #100;
A = 16'h004D; B = 16'h007D; #100;
A = 16'h004D; B = 16'h007E; #100;
A = 16'h004D; B = 16'h007F; #100;
A = 16'h004D; B = 16'h0080; #100;
A = 16'h004D; B = 16'h0081; #100;
A = 16'h004D; B = 16'h0082; #100;
A = 16'h004D; B = 16'h0083; #100;
A = 16'h004D; B = 16'h0084; #100;
A = 16'h004D; B = 16'h0085; #100;
A = 16'h004D; B = 16'h0086; #100;
A = 16'h004D; B = 16'h0087; #100;
A = 16'h004D; B = 16'h0088; #100;
A = 16'h004D; B = 16'h0089; #100;
A = 16'h004D; B = 16'h008A; #100;
A = 16'h004D; B = 16'h008B; #100;
A = 16'h004D; B = 16'h008C; #100;
A = 16'h004D; B = 16'h008D; #100;
A = 16'h004D; B = 16'h008E; #100;
A = 16'h004D; B = 16'h008F; #100;
A = 16'h004D; B = 16'h0090; #100;
A = 16'h004D; B = 16'h0091; #100;
A = 16'h004D; B = 16'h0092; #100;
A = 16'h004D; B = 16'h0093; #100;
A = 16'h004D; B = 16'h0094; #100;
A = 16'h004D; B = 16'h0095; #100;
A = 16'h004D; B = 16'h0096; #100;
A = 16'h004D; B = 16'h0097; #100;
A = 16'h004D; B = 16'h0098; #100;
A = 16'h004D; B = 16'h0099; #100;
A = 16'h004D; B = 16'h009A; #100;
A = 16'h004D; B = 16'h009B; #100;
A = 16'h004D; B = 16'h009C; #100;
A = 16'h004D; B = 16'h009D; #100;
A = 16'h004D; B = 16'h009E; #100;
A = 16'h004D; B = 16'h009F; #100;
A = 16'h004D; B = 16'h00A0; #100;
A = 16'h004D; B = 16'h00A1; #100;
A = 16'h004D; B = 16'h00A2; #100;
A = 16'h004D; B = 16'h00A3; #100;
A = 16'h004D; B = 16'h00A4; #100;
A = 16'h004D; B = 16'h00A5; #100;
A = 16'h004D; B = 16'h00A6; #100;
A = 16'h004D; B = 16'h00A7; #100;
A = 16'h004D; B = 16'h00A8; #100;
A = 16'h004D; B = 16'h00A9; #100;
A = 16'h004D; B = 16'h00AA; #100;
A = 16'h004D; B = 16'h00AB; #100;
A = 16'h004D; B = 16'h00AC; #100;
A = 16'h004D; B = 16'h00AD; #100;
A = 16'h004D; B = 16'h00AE; #100;
A = 16'h004D; B = 16'h00AF; #100;
A = 16'h004D; B = 16'h00B0; #100;
A = 16'h004D; B = 16'h00B1; #100;
A = 16'h004D; B = 16'h00B2; #100;
A = 16'h004D; B = 16'h00B3; #100;
A = 16'h004D; B = 16'h00B4; #100;
A = 16'h004D; B = 16'h00B5; #100;
A = 16'h004D; B = 16'h00B6; #100;
A = 16'h004D; B = 16'h00B7; #100;
A = 16'h004D; B = 16'h00B8; #100;
A = 16'h004D; B = 16'h00B9; #100;
A = 16'h004D; B = 16'h00BA; #100;
A = 16'h004D; B = 16'h00BB; #100;
A = 16'h004D; B = 16'h00BC; #100;
A = 16'h004D; B = 16'h00BD; #100;
A = 16'h004D; B = 16'h00BE; #100;
A = 16'h004D; B = 16'h00BF; #100;
A = 16'h004D; B = 16'h00C0; #100;
A = 16'h004D; B = 16'h00C1; #100;
A = 16'h004D; B = 16'h00C2; #100;
A = 16'h004D; B = 16'h00C3; #100;
A = 16'h004D; B = 16'h00C4; #100;
A = 16'h004D; B = 16'h00C5; #100;
A = 16'h004D; B = 16'h00C6; #100;
A = 16'h004D; B = 16'h00C7; #100;
A = 16'h004D; B = 16'h00C8; #100;
A = 16'h004D; B = 16'h00C9; #100;
A = 16'h004D; B = 16'h00CA; #100;
A = 16'h004D; B = 16'h00CB; #100;
A = 16'h004D; B = 16'h00CC; #100;
A = 16'h004D; B = 16'h00CD; #100;
A = 16'h004D; B = 16'h00CE; #100;
A = 16'h004D; B = 16'h00CF; #100;
A = 16'h004D; B = 16'h00D0; #100;
A = 16'h004D; B = 16'h00D1; #100;
A = 16'h004D; B = 16'h00D2; #100;
A = 16'h004D; B = 16'h00D3; #100;
A = 16'h004D; B = 16'h00D4; #100;
A = 16'h004D; B = 16'h00D5; #100;
A = 16'h004D; B = 16'h00D6; #100;
A = 16'h004D; B = 16'h00D7; #100;
A = 16'h004D; B = 16'h00D8; #100;
A = 16'h004D; B = 16'h00D9; #100;
A = 16'h004D; B = 16'h00DA; #100;
A = 16'h004D; B = 16'h00DB; #100;
A = 16'h004D; B = 16'h00DC; #100;
A = 16'h004D; B = 16'h00DD; #100;
A = 16'h004D; B = 16'h00DE; #100;
A = 16'h004D; B = 16'h00DF; #100;
A = 16'h004D; B = 16'h00E0; #100;
A = 16'h004D; B = 16'h00E1; #100;
A = 16'h004D; B = 16'h00E2; #100;
A = 16'h004D; B = 16'h00E3; #100;
A = 16'h004D; B = 16'h00E4; #100;
A = 16'h004D; B = 16'h00E5; #100;
A = 16'h004D; B = 16'h00E6; #100;
A = 16'h004D; B = 16'h00E7; #100;
A = 16'h004D; B = 16'h00E8; #100;
A = 16'h004D; B = 16'h00E9; #100;
A = 16'h004D; B = 16'h00EA; #100;
A = 16'h004D; B = 16'h00EB; #100;
A = 16'h004D; B = 16'h00EC; #100;
A = 16'h004D; B = 16'h00ED; #100;
A = 16'h004D; B = 16'h00EE; #100;
A = 16'h004D; B = 16'h00EF; #100;
A = 16'h004D; B = 16'h00F0; #100;
A = 16'h004D; B = 16'h00F1; #100;
A = 16'h004D; B = 16'h00F2; #100;
A = 16'h004D; B = 16'h00F3; #100;
A = 16'h004D; B = 16'h00F4; #100;
A = 16'h004D; B = 16'h00F5; #100;
A = 16'h004D; B = 16'h00F6; #100;
A = 16'h004D; B = 16'h00F7; #100;
A = 16'h004D; B = 16'h00F8; #100;
A = 16'h004D; B = 16'h00F9; #100;
A = 16'h004D; B = 16'h00FA; #100;
A = 16'h004D; B = 16'h00FB; #100;
A = 16'h004D; B = 16'h00FC; #100;
A = 16'h004D; B = 16'h00FD; #100;
A = 16'h004D; B = 16'h00FE; #100;
A = 16'h004D; B = 16'h00FF; #100;
A = 16'h004E; B = 16'h000; #100;
A = 16'h004E; B = 16'h001; #100;
A = 16'h004E; B = 16'h002; #100;
A = 16'h004E; B = 16'h003; #100;
A = 16'h004E; B = 16'h004; #100;
A = 16'h004E; B = 16'h005; #100;
A = 16'h004E; B = 16'h006; #100;
A = 16'h004E; B = 16'h007; #100;
A = 16'h004E; B = 16'h008; #100;
A = 16'h004E; B = 16'h009; #100;
A = 16'h004E; B = 16'h00A; #100;
A = 16'h004E; B = 16'h00B; #100;
A = 16'h004E; B = 16'h00C; #100;
A = 16'h004E; B = 16'h00D; #100;
A = 16'h004E; B = 16'h00E; #100;
A = 16'h004E; B = 16'h00F; #100;
A = 16'h004E; B = 16'h0010; #100;
A = 16'h004E; B = 16'h0011; #100;
A = 16'h004E; B = 16'h0012; #100;
A = 16'h004E; B = 16'h0013; #100;
A = 16'h004E; B = 16'h0014; #100;
A = 16'h004E; B = 16'h0015; #100;
A = 16'h004E; B = 16'h0016; #100;
A = 16'h004E; B = 16'h0017; #100;
A = 16'h004E; B = 16'h0018; #100;
A = 16'h004E; B = 16'h0019; #100;
A = 16'h004E; B = 16'h001A; #100;
A = 16'h004E; B = 16'h001B; #100;
A = 16'h004E; B = 16'h001C; #100;
A = 16'h004E; B = 16'h001D; #100;
A = 16'h004E; B = 16'h001E; #100;
A = 16'h004E; B = 16'h001F; #100;
A = 16'h004E; B = 16'h0020; #100;
A = 16'h004E; B = 16'h0021; #100;
A = 16'h004E; B = 16'h0022; #100;
A = 16'h004E; B = 16'h0023; #100;
A = 16'h004E; B = 16'h0024; #100;
A = 16'h004E; B = 16'h0025; #100;
A = 16'h004E; B = 16'h0026; #100;
A = 16'h004E; B = 16'h0027; #100;
A = 16'h004E; B = 16'h0028; #100;
A = 16'h004E; B = 16'h0029; #100;
A = 16'h004E; B = 16'h002A; #100;
A = 16'h004E; B = 16'h002B; #100;
A = 16'h004E; B = 16'h002C; #100;
A = 16'h004E; B = 16'h002D; #100;
A = 16'h004E; B = 16'h002E; #100;
A = 16'h004E; B = 16'h002F; #100;
A = 16'h004E; B = 16'h0030; #100;
A = 16'h004E; B = 16'h0031; #100;
A = 16'h004E; B = 16'h0032; #100;
A = 16'h004E; B = 16'h0033; #100;
A = 16'h004E; B = 16'h0034; #100;
A = 16'h004E; B = 16'h0035; #100;
A = 16'h004E; B = 16'h0036; #100;
A = 16'h004E; B = 16'h0037; #100;
A = 16'h004E; B = 16'h0038; #100;
A = 16'h004E; B = 16'h0039; #100;
A = 16'h004E; B = 16'h003A; #100;
A = 16'h004E; B = 16'h003B; #100;
A = 16'h004E; B = 16'h003C; #100;
A = 16'h004E; B = 16'h003D; #100;
A = 16'h004E; B = 16'h003E; #100;
A = 16'h004E; B = 16'h003F; #100;
A = 16'h004E; B = 16'h0040; #100;
A = 16'h004E; B = 16'h0041; #100;
A = 16'h004E; B = 16'h0042; #100;
A = 16'h004E; B = 16'h0043; #100;
A = 16'h004E; B = 16'h0044; #100;
A = 16'h004E; B = 16'h0045; #100;
A = 16'h004E; B = 16'h0046; #100;
A = 16'h004E; B = 16'h0047; #100;
A = 16'h004E; B = 16'h0048; #100;
A = 16'h004E; B = 16'h0049; #100;
A = 16'h004E; B = 16'h004A; #100;
A = 16'h004E; B = 16'h004B; #100;
A = 16'h004E; B = 16'h004C; #100;
A = 16'h004E; B = 16'h004D; #100;
A = 16'h004E; B = 16'h004E; #100;
A = 16'h004E; B = 16'h004F; #100;
A = 16'h004E; B = 16'h0050; #100;
A = 16'h004E; B = 16'h0051; #100;
A = 16'h004E; B = 16'h0052; #100;
A = 16'h004E; B = 16'h0053; #100;
A = 16'h004E; B = 16'h0054; #100;
A = 16'h004E; B = 16'h0055; #100;
A = 16'h004E; B = 16'h0056; #100;
A = 16'h004E; B = 16'h0057; #100;
A = 16'h004E; B = 16'h0058; #100;
A = 16'h004E; B = 16'h0059; #100;
A = 16'h004E; B = 16'h005A; #100;
A = 16'h004E; B = 16'h005B; #100;
A = 16'h004E; B = 16'h005C; #100;
A = 16'h004E; B = 16'h005D; #100;
A = 16'h004E; B = 16'h005E; #100;
A = 16'h004E; B = 16'h005F; #100;
A = 16'h004E; B = 16'h0060; #100;
A = 16'h004E; B = 16'h0061; #100;
A = 16'h004E; B = 16'h0062; #100;
A = 16'h004E; B = 16'h0063; #100;
A = 16'h004E; B = 16'h0064; #100;
A = 16'h004E; B = 16'h0065; #100;
A = 16'h004E; B = 16'h0066; #100;
A = 16'h004E; B = 16'h0067; #100;
A = 16'h004E; B = 16'h0068; #100;
A = 16'h004E; B = 16'h0069; #100;
A = 16'h004E; B = 16'h006A; #100;
A = 16'h004E; B = 16'h006B; #100;
A = 16'h004E; B = 16'h006C; #100;
A = 16'h004E; B = 16'h006D; #100;
A = 16'h004E; B = 16'h006E; #100;
A = 16'h004E; B = 16'h006F; #100;
A = 16'h004E; B = 16'h0070; #100;
A = 16'h004E; B = 16'h0071; #100;
A = 16'h004E; B = 16'h0072; #100;
A = 16'h004E; B = 16'h0073; #100;
A = 16'h004E; B = 16'h0074; #100;
A = 16'h004E; B = 16'h0075; #100;
A = 16'h004E; B = 16'h0076; #100;
A = 16'h004E; B = 16'h0077; #100;
A = 16'h004E; B = 16'h0078; #100;
A = 16'h004E; B = 16'h0079; #100;
A = 16'h004E; B = 16'h007A; #100;
A = 16'h004E; B = 16'h007B; #100;
A = 16'h004E; B = 16'h007C; #100;
A = 16'h004E; B = 16'h007D; #100;
A = 16'h004E; B = 16'h007E; #100;
A = 16'h004E; B = 16'h007F; #100;
A = 16'h004E; B = 16'h0080; #100;
A = 16'h004E; B = 16'h0081; #100;
A = 16'h004E; B = 16'h0082; #100;
A = 16'h004E; B = 16'h0083; #100;
A = 16'h004E; B = 16'h0084; #100;
A = 16'h004E; B = 16'h0085; #100;
A = 16'h004E; B = 16'h0086; #100;
A = 16'h004E; B = 16'h0087; #100;
A = 16'h004E; B = 16'h0088; #100;
A = 16'h004E; B = 16'h0089; #100;
A = 16'h004E; B = 16'h008A; #100;
A = 16'h004E; B = 16'h008B; #100;
A = 16'h004E; B = 16'h008C; #100;
A = 16'h004E; B = 16'h008D; #100;
A = 16'h004E; B = 16'h008E; #100;
A = 16'h004E; B = 16'h008F; #100;
A = 16'h004E; B = 16'h0090; #100;
A = 16'h004E; B = 16'h0091; #100;
A = 16'h004E; B = 16'h0092; #100;
A = 16'h004E; B = 16'h0093; #100;
A = 16'h004E; B = 16'h0094; #100;
A = 16'h004E; B = 16'h0095; #100;
A = 16'h004E; B = 16'h0096; #100;
A = 16'h004E; B = 16'h0097; #100;
A = 16'h004E; B = 16'h0098; #100;
A = 16'h004E; B = 16'h0099; #100;
A = 16'h004E; B = 16'h009A; #100;
A = 16'h004E; B = 16'h009B; #100;
A = 16'h004E; B = 16'h009C; #100;
A = 16'h004E; B = 16'h009D; #100;
A = 16'h004E; B = 16'h009E; #100;
A = 16'h004E; B = 16'h009F; #100;
A = 16'h004E; B = 16'h00A0; #100;
A = 16'h004E; B = 16'h00A1; #100;
A = 16'h004E; B = 16'h00A2; #100;
A = 16'h004E; B = 16'h00A3; #100;
A = 16'h004E; B = 16'h00A4; #100;
A = 16'h004E; B = 16'h00A5; #100;
A = 16'h004E; B = 16'h00A6; #100;
A = 16'h004E; B = 16'h00A7; #100;
A = 16'h004E; B = 16'h00A8; #100;
A = 16'h004E; B = 16'h00A9; #100;
A = 16'h004E; B = 16'h00AA; #100;
A = 16'h004E; B = 16'h00AB; #100;
A = 16'h004E; B = 16'h00AC; #100;
A = 16'h004E; B = 16'h00AD; #100;
A = 16'h004E; B = 16'h00AE; #100;
A = 16'h004E; B = 16'h00AF; #100;
A = 16'h004E; B = 16'h00B0; #100;
A = 16'h004E; B = 16'h00B1; #100;
A = 16'h004E; B = 16'h00B2; #100;
A = 16'h004E; B = 16'h00B3; #100;
A = 16'h004E; B = 16'h00B4; #100;
A = 16'h004E; B = 16'h00B5; #100;
A = 16'h004E; B = 16'h00B6; #100;
A = 16'h004E; B = 16'h00B7; #100;
A = 16'h004E; B = 16'h00B8; #100;
A = 16'h004E; B = 16'h00B9; #100;
A = 16'h004E; B = 16'h00BA; #100;
A = 16'h004E; B = 16'h00BB; #100;
A = 16'h004E; B = 16'h00BC; #100;
A = 16'h004E; B = 16'h00BD; #100;
A = 16'h004E; B = 16'h00BE; #100;
A = 16'h004E; B = 16'h00BF; #100;
A = 16'h004E; B = 16'h00C0; #100;
A = 16'h004E; B = 16'h00C1; #100;
A = 16'h004E; B = 16'h00C2; #100;
A = 16'h004E; B = 16'h00C3; #100;
A = 16'h004E; B = 16'h00C4; #100;
A = 16'h004E; B = 16'h00C5; #100;
A = 16'h004E; B = 16'h00C6; #100;
A = 16'h004E; B = 16'h00C7; #100;
A = 16'h004E; B = 16'h00C8; #100;
A = 16'h004E; B = 16'h00C9; #100;
A = 16'h004E; B = 16'h00CA; #100;
A = 16'h004E; B = 16'h00CB; #100;
A = 16'h004E; B = 16'h00CC; #100;
A = 16'h004E; B = 16'h00CD; #100;
A = 16'h004E; B = 16'h00CE; #100;
A = 16'h004E; B = 16'h00CF; #100;
A = 16'h004E; B = 16'h00D0; #100;
A = 16'h004E; B = 16'h00D1; #100;
A = 16'h004E; B = 16'h00D2; #100;
A = 16'h004E; B = 16'h00D3; #100;
A = 16'h004E; B = 16'h00D4; #100;
A = 16'h004E; B = 16'h00D5; #100;
A = 16'h004E; B = 16'h00D6; #100;
A = 16'h004E; B = 16'h00D7; #100;
A = 16'h004E; B = 16'h00D8; #100;
A = 16'h004E; B = 16'h00D9; #100;
A = 16'h004E; B = 16'h00DA; #100;
A = 16'h004E; B = 16'h00DB; #100;
A = 16'h004E; B = 16'h00DC; #100;
A = 16'h004E; B = 16'h00DD; #100;
A = 16'h004E; B = 16'h00DE; #100;
A = 16'h004E; B = 16'h00DF; #100;
A = 16'h004E; B = 16'h00E0; #100;
A = 16'h004E; B = 16'h00E1; #100;
A = 16'h004E; B = 16'h00E2; #100;
A = 16'h004E; B = 16'h00E3; #100;
A = 16'h004E; B = 16'h00E4; #100;
A = 16'h004E; B = 16'h00E5; #100;
A = 16'h004E; B = 16'h00E6; #100;
A = 16'h004E; B = 16'h00E7; #100;
A = 16'h004E; B = 16'h00E8; #100;
A = 16'h004E; B = 16'h00E9; #100;
A = 16'h004E; B = 16'h00EA; #100;
A = 16'h004E; B = 16'h00EB; #100;
A = 16'h004E; B = 16'h00EC; #100;
A = 16'h004E; B = 16'h00ED; #100;
A = 16'h004E; B = 16'h00EE; #100;
A = 16'h004E; B = 16'h00EF; #100;
A = 16'h004E; B = 16'h00F0; #100;
A = 16'h004E; B = 16'h00F1; #100;
A = 16'h004E; B = 16'h00F2; #100;
A = 16'h004E; B = 16'h00F3; #100;
A = 16'h004E; B = 16'h00F4; #100;
A = 16'h004E; B = 16'h00F5; #100;
A = 16'h004E; B = 16'h00F6; #100;
A = 16'h004E; B = 16'h00F7; #100;
A = 16'h004E; B = 16'h00F8; #100;
A = 16'h004E; B = 16'h00F9; #100;
A = 16'h004E; B = 16'h00FA; #100;
A = 16'h004E; B = 16'h00FB; #100;
A = 16'h004E; B = 16'h00FC; #100;
A = 16'h004E; B = 16'h00FD; #100;
A = 16'h004E; B = 16'h00FE; #100;
A = 16'h004E; B = 16'h00FF; #100;
A = 16'h004F; B = 16'h000; #100;
A = 16'h004F; B = 16'h001; #100;
A = 16'h004F; B = 16'h002; #100;
A = 16'h004F; B = 16'h003; #100;
A = 16'h004F; B = 16'h004; #100;
A = 16'h004F; B = 16'h005; #100;
A = 16'h004F; B = 16'h006; #100;
A = 16'h004F; B = 16'h007; #100;
A = 16'h004F; B = 16'h008; #100;
A = 16'h004F; B = 16'h009; #100;
A = 16'h004F; B = 16'h00A; #100;
A = 16'h004F; B = 16'h00B; #100;
A = 16'h004F; B = 16'h00C; #100;
A = 16'h004F; B = 16'h00D; #100;
A = 16'h004F; B = 16'h00E; #100;
A = 16'h004F; B = 16'h00F; #100;
A = 16'h004F; B = 16'h0010; #100;
A = 16'h004F; B = 16'h0011; #100;
A = 16'h004F; B = 16'h0012; #100;
A = 16'h004F; B = 16'h0013; #100;
A = 16'h004F; B = 16'h0014; #100;
A = 16'h004F; B = 16'h0015; #100;
A = 16'h004F; B = 16'h0016; #100;
A = 16'h004F; B = 16'h0017; #100;
A = 16'h004F; B = 16'h0018; #100;
A = 16'h004F; B = 16'h0019; #100;
A = 16'h004F; B = 16'h001A; #100;
A = 16'h004F; B = 16'h001B; #100;
A = 16'h004F; B = 16'h001C; #100;
A = 16'h004F; B = 16'h001D; #100;
A = 16'h004F; B = 16'h001E; #100;
A = 16'h004F; B = 16'h001F; #100;
A = 16'h004F; B = 16'h0020; #100;
A = 16'h004F; B = 16'h0021; #100;
A = 16'h004F; B = 16'h0022; #100;
A = 16'h004F; B = 16'h0023; #100;
A = 16'h004F; B = 16'h0024; #100;
A = 16'h004F; B = 16'h0025; #100;
A = 16'h004F; B = 16'h0026; #100;
A = 16'h004F; B = 16'h0027; #100;
A = 16'h004F; B = 16'h0028; #100;
A = 16'h004F; B = 16'h0029; #100;
A = 16'h004F; B = 16'h002A; #100;
A = 16'h004F; B = 16'h002B; #100;
A = 16'h004F; B = 16'h002C; #100;
A = 16'h004F; B = 16'h002D; #100;
A = 16'h004F; B = 16'h002E; #100;
A = 16'h004F; B = 16'h002F; #100;
A = 16'h004F; B = 16'h0030; #100;
A = 16'h004F; B = 16'h0031; #100;
A = 16'h004F; B = 16'h0032; #100;
A = 16'h004F; B = 16'h0033; #100;
A = 16'h004F; B = 16'h0034; #100;
A = 16'h004F; B = 16'h0035; #100;
A = 16'h004F; B = 16'h0036; #100;
A = 16'h004F; B = 16'h0037; #100;
A = 16'h004F; B = 16'h0038; #100;
A = 16'h004F; B = 16'h0039; #100;
A = 16'h004F; B = 16'h003A; #100;
A = 16'h004F; B = 16'h003B; #100;
A = 16'h004F; B = 16'h003C; #100;
A = 16'h004F; B = 16'h003D; #100;
A = 16'h004F; B = 16'h003E; #100;
A = 16'h004F; B = 16'h003F; #100;
A = 16'h004F; B = 16'h0040; #100;
A = 16'h004F; B = 16'h0041; #100;
A = 16'h004F; B = 16'h0042; #100;
A = 16'h004F; B = 16'h0043; #100;
A = 16'h004F; B = 16'h0044; #100;
A = 16'h004F; B = 16'h0045; #100;
A = 16'h004F; B = 16'h0046; #100;
A = 16'h004F; B = 16'h0047; #100;
A = 16'h004F; B = 16'h0048; #100;
A = 16'h004F; B = 16'h0049; #100;
A = 16'h004F; B = 16'h004A; #100;
A = 16'h004F; B = 16'h004B; #100;
A = 16'h004F; B = 16'h004C; #100;
A = 16'h004F; B = 16'h004D; #100;
A = 16'h004F; B = 16'h004E; #100;
A = 16'h004F; B = 16'h004F; #100;
A = 16'h004F; B = 16'h0050; #100;
A = 16'h004F; B = 16'h0051; #100;
A = 16'h004F; B = 16'h0052; #100;
A = 16'h004F; B = 16'h0053; #100;
A = 16'h004F; B = 16'h0054; #100;
A = 16'h004F; B = 16'h0055; #100;
A = 16'h004F; B = 16'h0056; #100;
A = 16'h004F; B = 16'h0057; #100;
A = 16'h004F; B = 16'h0058; #100;
A = 16'h004F; B = 16'h0059; #100;
A = 16'h004F; B = 16'h005A; #100;
A = 16'h004F; B = 16'h005B; #100;
A = 16'h004F; B = 16'h005C; #100;
A = 16'h004F; B = 16'h005D; #100;
A = 16'h004F; B = 16'h005E; #100;
A = 16'h004F; B = 16'h005F; #100;
A = 16'h004F; B = 16'h0060; #100;
A = 16'h004F; B = 16'h0061; #100;
A = 16'h004F; B = 16'h0062; #100;
A = 16'h004F; B = 16'h0063; #100;
A = 16'h004F; B = 16'h0064; #100;
A = 16'h004F; B = 16'h0065; #100;
A = 16'h004F; B = 16'h0066; #100;
A = 16'h004F; B = 16'h0067; #100;
A = 16'h004F; B = 16'h0068; #100;
A = 16'h004F; B = 16'h0069; #100;
A = 16'h004F; B = 16'h006A; #100;
A = 16'h004F; B = 16'h006B; #100;
A = 16'h004F; B = 16'h006C; #100;
A = 16'h004F; B = 16'h006D; #100;
A = 16'h004F; B = 16'h006E; #100;
A = 16'h004F; B = 16'h006F; #100;
A = 16'h004F; B = 16'h0070; #100;
A = 16'h004F; B = 16'h0071; #100;
A = 16'h004F; B = 16'h0072; #100;
A = 16'h004F; B = 16'h0073; #100;
A = 16'h004F; B = 16'h0074; #100;
A = 16'h004F; B = 16'h0075; #100;
A = 16'h004F; B = 16'h0076; #100;
A = 16'h004F; B = 16'h0077; #100;
A = 16'h004F; B = 16'h0078; #100;
A = 16'h004F; B = 16'h0079; #100;
A = 16'h004F; B = 16'h007A; #100;
A = 16'h004F; B = 16'h007B; #100;
A = 16'h004F; B = 16'h007C; #100;
A = 16'h004F; B = 16'h007D; #100;
A = 16'h004F; B = 16'h007E; #100;
A = 16'h004F; B = 16'h007F; #100;
A = 16'h004F; B = 16'h0080; #100;
A = 16'h004F; B = 16'h0081; #100;
A = 16'h004F; B = 16'h0082; #100;
A = 16'h004F; B = 16'h0083; #100;
A = 16'h004F; B = 16'h0084; #100;
A = 16'h004F; B = 16'h0085; #100;
A = 16'h004F; B = 16'h0086; #100;
A = 16'h004F; B = 16'h0087; #100;
A = 16'h004F; B = 16'h0088; #100;
A = 16'h004F; B = 16'h0089; #100;
A = 16'h004F; B = 16'h008A; #100;
A = 16'h004F; B = 16'h008B; #100;
A = 16'h004F; B = 16'h008C; #100;
A = 16'h004F; B = 16'h008D; #100;
A = 16'h004F; B = 16'h008E; #100;
A = 16'h004F; B = 16'h008F; #100;
A = 16'h004F; B = 16'h0090; #100;
A = 16'h004F; B = 16'h0091; #100;
A = 16'h004F; B = 16'h0092; #100;
A = 16'h004F; B = 16'h0093; #100;
A = 16'h004F; B = 16'h0094; #100;
A = 16'h004F; B = 16'h0095; #100;
A = 16'h004F; B = 16'h0096; #100;
A = 16'h004F; B = 16'h0097; #100;
A = 16'h004F; B = 16'h0098; #100;
A = 16'h004F; B = 16'h0099; #100;
A = 16'h004F; B = 16'h009A; #100;
A = 16'h004F; B = 16'h009B; #100;
A = 16'h004F; B = 16'h009C; #100;
A = 16'h004F; B = 16'h009D; #100;
A = 16'h004F; B = 16'h009E; #100;
A = 16'h004F; B = 16'h009F; #100;
A = 16'h004F; B = 16'h00A0; #100;
A = 16'h004F; B = 16'h00A1; #100;
A = 16'h004F; B = 16'h00A2; #100;
A = 16'h004F; B = 16'h00A3; #100;
A = 16'h004F; B = 16'h00A4; #100;
A = 16'h004F; B = 16'h00A5; #100;
A = 16'h004F; B = 16'h00A6; #100;
A = 16'h004F; B = 16'h00A7; #100;
A = 16'h004F; B = 16'h00A8; #100;
A = 16'h004F; B = 16'h00A9; #100;
A = 16'h004F; B = 16'h00AA; #100;
A = 16'h004F; B = 16'h00AB; #100;
A = 16'h004F; B = 16'h00AC; #100;
A = 16'h004F; B = 16'h00AD; #100;
A = 16'h004F; B = 16'h00AE; #100;
A = 16'h004F; B = 16'h00AF; #100;
A = 16'h004F; B = 16'h00B0; #100;
A = 16'h004F; B = 16'h00B1; #100;
A = 16'h004F; B = 16'h00B2; #100;
A = 16'h004F; B = 16'h00B3; #100;
A = 16'h004F; B = 16'h00B4; #100;
A = 16'h004F; B = 16'h00B5; #100;
A = 16'h004F; B = 16'h00B6; #100;
A = 16'h004F; B = 16'h00B7; #100;
A = 16'h004F; B = 16'h00B8; #100;
A = 16'h004F; B = 16'h00B9; #100;
A = 16'h004F; B = 16'h00BA; #100;
A = 16'h004F; B = 16'h00BB; #100;
A = 16'h004F; B = 16'h00BC; #100;
A = 16'h004F; B = 16'h00BD; #100;
A = 16'h004F; B = 16'h00BE; #100;
A = 16'h004F; B = 16'h00BF; #100;
A = 16'h004F; B = 16'h00C0; #100;
A = 16'h004F; B = 16'h00C1; #100;
A = 16'h004F; B = 16'h00C2; #100;
A = 16'h004F; B = 16'h00C3; #100;
A = 16'h004F; B = 16'h00C4; #100;
A = 16'h004F; B = 16'h00C5; #100;
A = 16'h004F; B = 16'h00C6; #100;
A = 16'h004F; B = 16'h00C7; #100;
A = 16'h004F; B = 16'h00C8; #100;
A = 16'h004F; B = 16'h00C9; #100;
A = 16'h004F; B = 16'h00CA; #100;
A = 16'h004F; B = 16'h00CB; #100;
A = 16'h004F; B = 16'h00CC; #100;
A = 16'h004F; B = 16'h00CD; #100;
A = 16'h004F; B = 16'h00CE; #100;
A = 16'h004F; B = 16'h00CF; #100;
A = 16'h004F; B = 16'h00D0; #100;
A = 16'h004F; B = 16'h00D1; #100;
A = 16'h004F; B = 16'h00D2; #100;
A = 16'h004F; B = 16'h00D3; #100;
A = 16'h004F; B = 16'h00D4; #100;
A = 16'h004F; B = 16'h00D5; #100;
A = 16'h004F; B = 16'h00D6; #100;
A = 16'h004F; B = 16'h00D7; #100;
A = 16'h004F; B = 16'h00D8; #100;
A = 16'h004F; B = 16'h00D9; #100;
A = 16'h004F; B = 16'h00DA; #100;
A = 16'h004F; B = 16'h00DB; #100;
A = 16'h004F; B = 16'h00DC; #100;
A = 16'h004F; B = 16'h00DD; #100;
A = 16'h004F; B = 16'h00DE; #100;
A = 16'h004F; B = 16'h00DF; #100;
A = 16'h004F; B = 16'h00E0; #100;
A = 16'h004F; B = 16'h00E1; #100;
A = 16'h004F; B = 16'h00E2; #100;
A = 16'h004F; B = 16'h00E3; #100;
A = 16'h004F; B = 16'h00E4; #100;
A = 16'h004F; B = 16'h00E5; #100;
A = 16'h004F; B = 16'h00E6; #100;
A = 16'h004F; B = 16'h00E7; #100;
A = 16'h004F; B = 16'h00E8; #100;
A = 16'h004F; B = 16'h00E9; #100;
A = 16'h004F; B = 16'h00EA; #100;
A = 16'h004F; B = 16'h00EB; #100;
A = 16'h004F; B = 16'h00EC; #100;
A = 16'h004F; B = 16'h00ED; #100;
A = 16'h004F; B = 16'h00EE; #100;
A = 16'h004F; B = 16'h00EF; #100;
A = 16'h004F; B = 16'h00F0; #100;
A = 16'h004F; B = 16'h00F1; #100;
A = 16'h004F; B = 16'h00F2; #100;
A = 16'h004F; B = 16'h00F3; #100;
A = 16'h004F; B = 16'h00F4; #100;
A = 16'h004F; B = 16'h00F5; #100;
A = 16'h004F; B = 16'h00F6; #100;
A = 16'h004F; B = 16'h00F7; #100;
A = 16'h004F; B = 16'h00F8; #100;
A = 16'h004F; B = 16'h00F9; #100;
A = 16'h004F; B = 16'h00FA; #100;
A = 16'h004F; B = 16'h00FB; #100;
A = 16'h004F; B = 16'h00FC; #100;
A = 16'h004F; B = 16'h00FD; #100;
A = 16'h004F; B = 16'h00FE; #100;
A = 16'h004F; B = 16'h00FF; #100;
A = 16'h0050; B = 16'h000; #100;
A = 16'h0050; B = 16'h001; #100;
A = 16'h0050; B = 16'h002; #100;
A = 16'h0050; B = 16'h003; #100;
A = 16'h0050; B = 16'h004; #100;
A = 16'h0050; B = 16'h005; #100;
A = 16'h0050; B = 16'h006; #100;
A = 16'h0050; B = 16'h007; #100;
A = 16'h0050; B = 16'h008; #100;
A = 16'h0050; B = 16'h009; #100;
A = 16'h0050; B = 16'h00A; #100;
A = 16'h0050; B = 16'h00B; #100;
A = 16'h0050; B = 16'h00C; #100;
A = 16'h0050; B = 16'h00D; #100;
A = 16'h0050; B = 16'h00E; #100;
A = 16'h0050; B = 16'h00F; #100;
A = 16'h0050; B = 16'h0010; #100;
A = 16'h0050; B = 16'h0011; #100;
A = 16'h0050; B = 16'h0012; #100;
A = 16'h0050; B = 16'h0013; #100;
A = 16'h0050; B = 16'h0014; #100;
A = 16'h0050; B = 16'h0015; #100;
A = 16'h0050; B = 16'h0016; #100;
A = 16'h0050; B = 16'h0017; #100;
A = 16'h0050; B = 16'h0018; #100;
A = 16'h0050; B = 16'h0019; #100;
A = 16'h0050; B = 16'h001A; #100;
A = 16'h0050; B = 16'h001B; #100;
A = 16'h0050; B = 16'h001C; #100;
A = 16'h0050; B = 16'h001D; #100;
A = 16'h0050; B = 16'h001E; #100;
A = 16'h0050; B = 16'h001F; #100;
A = 16'h0050; B = 16'h0020; #100;
A = 16'h0050; B = 16'h0021; #100;
A = 16'h0050; B = 16'h0022; #100;
A = 16'h0050; B = 16'h0023; #100;
A = 16'h0050; B = 16'h0024; #100;
A = 16'h0050; B = 16'h0025; #100;
A = 16'h0050; B = 16'h0026; #100;
A = 16'h0050; B = 16'h0027; #100;
A = 16'h0050; B = 16'h0028; #100;
A = 16'h0050; B = 16'h0029; #100;
A = 16'h0050; B = 16'h002A; #100;
A = 16'h0050; B = 16'h002B; #100;
A = 16'h0050; B = 16'h002C; #100;
A = 16'h0050; B = 16'h002D; #100;
A = 16'h0050; B = 16'h002E; #100;
A = 16'h0050; B = 16'h002F; #100;
A = 16'h0050; B = 16'h0030; #100;
A = 16'h0050; B = 16'h0031; #100;
A = 16'h0050; B = 16'h0032; #100;
A = 16'h0050; B = 16'h0033; #100;
A = 16'h0050; B = 16'h0034; #100;
A = 16'h0050; B = 16'h0035; #100;
A = 16'h0050; B = 16'h0036; #100;
A = 16'h0050; B = 16'h0037; #100;
A = 16'h0050; B = 16'h0038; #100;
A = 16'h0050; B = 16'h0039; #100;
A = 16'h0050; B = 16'h003A; #100;
A = 16'h0050; B = 16'h003B; #100;
A = 16'h0050; B = 16'h003C; #100;
A = 16'h0050; B = 16'h003D; #100;
A = 16'h0050; B = 16'h003E; #100;
A = 16'h0050; B = 16'h003F; #100;
A = 16'h0050; B = 16'h0040; #100;
A = 16'h0050; B = 16'h0041; #100;
A = 16'h0050; B = 16'h0042; #100;
A = 16'h0050; B = 16'h0043; #100;
A = 16'h0050; B = 16'h0044; #100;
A = 16'h0050; B = 16'h0045; #100;
A = 16'h0050; B = 16'h0046; #100;
A = 16'h0050; B = 16'h0047; #100;
A = 16'h0050; B = 16'h0048; #100;
A = 16'h0050; B = 16'h0049; #100;
A = 16'h0050; B = 16'h004A; #100;
A = 16'h0050; B = 16'h004B; #100;
A = 16'h0050; B = 16'h004C; #100;
A = 16'h0050; B = 16'h004D; #100;
A = 16'h0050; B = 16'h004E; #100;
A = 16'h0050; B = 16'h004F; #100;
A = 16'h0050; B = 16'h0050; #100;
A = 16'h0050; B = 16'h0051; #100;
A = 16'h0050; B = 16'h0052; #100;
A = 16'h0050; B = 16'h0053; #100;
A = 16'h0050; B = 16'h0054; #100;
A = 16'h0050; B = 16'h0055; #100;
A = 16'h0050; B = 16'h0056; #100;
A = 16'h0050; B = 16'h0057; #100;
A = 16'h0050; B = 16'h0058; #100;
A = 16'h0050; B = 16'h0059; #100;
A = 16'h0050; B = 16'h005A; #100;
A = 16'h0050; B = 16'h005B; #100;
A = 16'h0050; B = 16'h005C; #100;
A = 16'h0050; B = 16'h005D; #100;
A = 16'h0050; B = 16'h005E; #100;
A = 16'h0050; B = 16'h005F; #100;
A = 16'h0050; B = 16'h0060; #100;
A = 16'h0050; B = 16'h0061; #100;
A = 16'h0050; B = 16'h0062; #100;
A = 16'h0050; B = 16'h0063; #100;
A = 16'h0050; B = 16'h0064; #100;
A = 16'h0050; B = 16'h0065; #100;
A = 16'h0050; B = 16'h0066; #100;
A = 16'h0050; B = 16'h0067; #100;
A = 16'h0050; B = 16'h0068; #100;
A = 16'h0050; B = 16'h0069; #100;
A = 16'h0050; B = 16'h006A; #100;
A = 16'h0050; B = 16'h006B; #100;
A = 16'h0050; B = 16'h006C; #100;
A = 16'h0050; B = 16'h006D; #100;
A = 16'h0050; B = 16'h006E; #100;
A = 16'h0050; B = 16'h006F; #100;
A = 16'h0050; B = 16'h0070; #100;
A = 16'h0050; B = 16'h0071; #100;
A = 16'h0050; B = 16'h0072; #100;
A = 16'h0050; B = 16'h0073; #100;
A = 16'h0050; B = 16'h0074; #100;
A = 16'h0050; B = 16'h0075; #100;
A = 16'h0050; B = 16'h0076; #100;
A = 16'h0050; B = 16'h0077; #100;
A = 16'h0050; B = 16'h0078; #100;
A = 16'h0050; B = 16'h0079; #100;
A = 16'h0050; B = 16'h007A; #100;
A = 16'h0050; B = 16'h007B; #100;
A = 16'h0050; B = 16'h007C; #100;
A = 16'h0050; B = 16'h007D; #100;
A = 16'h0050; B = 16'h007E; #100;
A = 16'h0050; B = 16'h007F; #100;
A = 16'h0050; B = 16'h0080; #100;
A = 16'h0050; B = 16'h0081; #100;
A = 16'h0050; B = 16'h0082; #100;
A = 16'h0050; B = 16'h0083; #100;
A = 16'h0050; B = 16'h0084; #100;
A = 16'h0050; B = 16'h0085; #100;
A = 16'h0050; B = 16'h0086; #100;
A = 16'h0050; B = 16'h0087; #100;
A = 16'h0050; B = 16'h0088; #100;
A = 16'h0050; B = 16'h0089; #100;
A = 16'h0050; B = 16'h008A; #100;
A = 16'h0050; B = 16'h008B; #100;
A = 16'h0050; B = 16'h008C; #100;
A = 16'h0050; B = 16'h008D; #100;
A = 16'h0050; B = 16'h008E; #100;
A = 16'h0050; B = 16'h008F; #100;
A = 16'h0050; B = 16'h0090; #100;
A = 16'h0050; B = 16'h0091; #100;
A = 16'h0050; B = 16'h0092; #100;
A = 16'h0050; B = 16'h0093; #100;
A = 16'h0050; B = 16'h0094; #100;
A = 16'h0050; B = 16'h0095; #100;
A = 16'h0050; B = 16'h0096; #100;
A = 16'h0050; B = 16'h0097; #100;
A = 16'h0050; B = 16'h0098; #100;
A = 16'h0050; B = 16'h0099; #100;
A = 16'h0050; B = 16'h009A; #100;
A = 16'h0050; B = 16'h009B; #100;
A = 16'h0050; B = 16'h009C; #100;
A = 16'h0050; B = 16'h009D; #100;
A = 16'h0050; B = 16'h009E; #100;
A = 16'h0050; B = 16'h009F; #100;
A = 16'h0050; B = 16'h00A0; #100;
A = 16'h0050; B = 16'h00A1; #100;
A = 16'h0050; B = 16'h00A2; #100;
A = 16'h0050; B = 16'h00A3; #100;
A = 16'h0050; B = 16'h00A4; #100;
A = 16'h0050; B = 16'h00A5; #100;
A = 16'h0050; B = 16'h00A6; #100;
A = 16'h0050; B = 16'h00A7; #100;
A = 16'h0050; B = 16'h00A8; #100;
A = 16'h0050; B = 16'h00A9; #100;
A = 16'h0050; B = 16'h00AA; #100;
A = 16'h0050; B = 16'h00AB; #100;
A = 16'h0050; B = 16'h00AC; #100;
A = 16'h0050; B = 16'h00AD; #100;
A = 16'h0050; B = 16'h00AE; #100;
A = 16'h0050; B = 16'h00AF; #100;
A = 16'h0050; B = 16'h00B0; #100;
A = 16'h0050; B = 16'h00B1; #100;
A = 16'h0050; B = 16'h00B2; #100;
A = 16'h0050; B = 16'h00B3; #100;
A = 16'h0050; B = 16'h00B4; #100;
A = 16'h0050; B = 16'h00B5; #100;
A = 16'h0050; B = 16'h00B6; #100;
A = 16'h0050; B = 16'h00B7; #100;
A = 16'h0050; B = 16'h00B8; #100;
A = 16'h0050; B = 16'h00B9; #100;
A = 16'h0050; B = 16'h00BA; #100;
A = 16'h0050; B = 16'h00BB; #100;
A = 16'h0050; B = 16'h00BC; #100;
A = 16'h0050; B = 16'h00BD; #100;
A = 16'h0050; B = 16'h00BE; #100;
A = 16'h0050; B = 16'h00BF; #100;
A = 16'h0050; B = 16'h00C0; #100;
A = 16'h0050; B = 16'h00C1; #100;
A = 16'h0050; B = 16'h00C2; #100;
A = 16'h0050; B = 16'h00C3; #100;
A = 16'h0050; B = 16'h00C4; #100;
A = 16'h0050; B = 16'h00C5; #100;
A = 16'h0050; B = 16'h00C6; #100;
A = 16'h0050; B = 16'h00C7; #100;
A = 16'h0050; B = 16'h00C8; #100;
A = 16'h0050; B = 16'h00C9; #100;
A = 16'h0050; B = 16'h00CA; #100;
A = 16'h0050; B = 16'h00CB; #100;
A = 16'h0050; B = 16'h00CC; #100;
A = 16'h0050; B = 16'h00CD; #100;
A = 16'h0050; B = 16'h00CE; #100;
A = 16'h0050; B = 16'h00CF; #100;
A = 16'h0050; B = 16'h00D0; #100;
A = 16'h0050; B = 16'h00D1; #100;
A = 16'h0050; B = 16'h00D2; #100;
A = 16'h0050; B = 16'h00D3; #100;
A = 16'h0050; B = 16'h00D4; #100;
A = 16'h0050; B = 16'h00D5; #100;
A = 16'h0050; B = 16'h00D6; #100;
A = 16'h0050; B = 16'h00D7; #100;
A = 16'h0050; B = 16'h00D8; #100;
A = 16'h0050; B = 16'h00D9; #100;
A = 16'h0050; B = 16'h00DA; #100;
A = 16'h0050; B = 16'h00DB; #100;
A = 16'h0050; B = 16'h00DC; #100;
A = 16'h0050; B = 16'h00DD; #100;
A = 16'h0050; B = 16'h00DE; #100;
A = 16'h0050; B = 16'h00DF; #100;
A = 16'h0050; B = 16'h00E0; #100;
A = 16'h0050; B = 16'h00E1; #100;
A = 16'h0050; B = 16'h00E2; #100;
A = 16'h0050; B = 16'h00E3; #100;
A = 16'h0050; B = 16'h00E4; #100;
A = 16'h0050; B = 16'h00E5; #100;
A = 16'h0050; B = 16'h00E6; #100;
A = 16'h0050; B = 16'h00E7; #100;
A = 16'h0050; B = 16'h00E8; #100;
A = 16'h0050; B = 16'h00E9; #100;
A = 16'h0050; B = 16'h00EA; #100;
A = 16'h0050; B = 16'h00EB; #100;
A = 16'h0050; B = 16'h00EC; #100;
A = 16'h0050; B = 16'h00ED; #100;
A = 16'h0050; B = 16'h00EE; #100;
A = 16'h0050; B = 16'h00EF; #100;
A = 16'h0050; B = 16'h00F0; #100;
A = 16'h0050; B = 16'h00F1; #100;
A = 16'h0050; B = 16'h00F2; #100;
A = 16'h0050; B = 16'h00F3; #100;
A = 16'h0050; B = 16'h00F4; #100;
A = 16'h0050; B = 16'h00F5; #100;
A = 16'h0050; B = 16'h00F6; #100;
A = 16'h0050; B = 16'h00F7; #100;
A = 16'h0050; B = 16'h00F8; #100;
A = 16'h0050; B = 16'h00F9; #100;
A = 16'h0050; B = 16'h00FA; #100;
A = 16'h0050; B = 16'h00FB; #100;
A = 16'h0050; B = 16'h00FC; #100;
A = 16'h0050; B = 16'h00FD; #100;
A = 16'h0050; B = 16'h00FE; #100;
A = 16'h0050; B = 16'h00FF; #100;
A = 16'h0051; B = 16'h000; #100;
A = 16'h0051; B = 16'h001; #100;
A = 16'h0051; B = 16'h002; #100;
A = 16'h0051; B = 16'h003; #100;
A = 16'h0051; B = 16'h004; #100;
A = 16'h0051; B = 16'h005; #100;
A = 16'h0051; B = 16'h006; #100;
A = 16'h0051; B = 16'h007; #100;
A = 16'h0051; B = 16'h008; #100;
A = 16'h0051; B = 16'h009; #100;
A = 16'h0051; B = 16'h00A; #100;
A = 16'h0051; B = 16'h00B; #100;
A = 16'h0051; B = 16'h00C; #100;
A = 16'h0051; B = 16'h00D; #100;
A = 16'h0051; B = 16'h00E; #100;
A = 16'h0051; B = 16'h00F; #100;
A = 16'h0051; B = 16'h0010; #100;
A = 16'h0051; B = 16'h0011; #100;
A = 16'h0051; B = 16'h0012; #100;
A = 16'h0051; B = 16'h0013; #100;
A = 16'h0051; B = 16'h0014; #100;
A = 16'h0051; B = 16'h0015; #100;
A = 16'h0051; B = 16'h0016; #100;
A = 16'h0051; B = 16'h0017; #100;
A = 16'h0051; B = 16'h0018; #100;
A = 16'h0051; B = 16'h0019; #100;
A = 16'h0051; B = 16'h001A; #100;
A = 16'h0051; B = 16'h001B; #100;
A = 16'h0051; B = 16'h001C; #100;
A = 16'h0051; B = 16'h001D; #100;
A = 16'h0051; B = 16'h001E; #100;
A = 16'h0051; B = 16'h001F; #100;
A = 16'h0051; B = 16'h0020; #100;
A = 16'h0051; B = 16'h0021; #100;
A = 16'h0051; B = 16'h0022; #100;
A = 16'h0051; B = 16'h0023; #100;
A = 16'h0051; B = 16'h0024; #100;
A = 16'h0051; B = 16'h0025; #100;
A = 16'h0051; B = 16'h0026; #100;
A = 16'h0051; B = 16'h0027; #100;
A = 16'h0051; B = 16'h0028; #100;
A = 16'h0051; B = 16'h0029; #100;
A = 16'h0051; B = 16'h002A; #100;
A = 16'h0051; B = 16'h002B; #100;
A = 16'h0051; B = 16'h002C; #100;
A = 16'h0051; B = 16'h002D; #100;
A = 16'h0051; B = 16'h002E; #100;
A = 16'h0051; B = 16'h002F; #100;
A = 16'h0051; B = 16'h0030; #100;
A = 16'h0051; B = 16'h0031; #100;
A = 16'h0051; B = 16'h0032; #100;
A = 16'h0051; B = 16'h0033; #100;
A = 16'h0051; B = 16'h0034; #100;
A = 16'h0051; B = 16'h0035; #100;
A = 16'h0051; B = 16'h0036; #100;
A = 16'h0051; B = 16'h0037; #100;
A = 16'h0051; B = 16'h0038; #100;
A = 16'h0051; B = 16'h0039; #100;
A = 16'h0051; B = 16'h003A; #100;
A = 16'h0051; B = 16'h003B; #100;
A = 16'h0051; B = 16'h003C; #100;
A = 16'h0051; B = 16'h003D; #100;
A = 16'h0051; B = 16'h003E; #100;
A = 16'h0051; B = 16'h003F; #100;
A = 16'h0051; B = 16'h0040; #100;
A = 16'h0051; B = 16'h0041; #100;
A = 16'h0051; B = 16'h0042; #100;
A = 16'h0051; B = 16'h0043; #100;
A = 16'h0051; B = 16'h0044; #100;
A = 16'h0051; B = 16'h0045; #100;
A = 16'h0051; B = 16'h0046; #100;
A = 16'h0051; B = 16'h0047; #100;
A = 16'h0051; B = 16'h0048; #100;
A = 16'h0051; B = 16'h0049; #100;
A = 16'h0051; B = 16'h004A; #100;
A = 16'h0051; B = 16'h004B; #100;
A = 16'h0051; B = 16'h004C; #100;
A = 16'h0051; B = 16'h004D; #100;
A = 16'h0051; B = 16'h004E; #100;
A = 16'h0051; B = 16'h004F; #100;
A = 16'h0051; B = 16'h0050; #100;
A = 16'h0051; B = 16'h0051; #100;
A = 16'h0051; B = 16'h0052; #100;
A = 16'h0051; B = 16'h0053; #100;
A = 16'h0051; B = 16'h0054; #100;
A = 16'h0051; B = 16'h0055; #100;
A = 16'h0051; B = 16'h0056; #100;
A = 16'h0051; B = 16'h0057; #100;
A = 16'h0051; B = 16'h0058; #100;
A = 16'h0051; B = 16'h0059; #100;
A = 16'h0051; B = 16'h005A; #100;
A = 16'h0051; B = 16'h005B; #100;
A = 16'h0051; B = 16'h005C; #100;
A = 16'h0051; B = 16'h005D; #100;
A = 16'h0051; B = 16'h005E; #100;
A = 16'h0051; B = 16'h005F; #100;
A = 16'h0051; B = 16'h0060; #100;
A = 16'h0051; B = 16'h0061; #100;
A = 16'h0051; B = 16'h0062; #100;
A = 16'h0051; B = 16'h0063; #100;
A = 16'h0051; B = 16'h0064; #100;
A = 16'h0051; B = 16'h0065; #100;
A = 16'h0051; B = 16'h0066; #100;
A = 16'h0051; B = 16'h0067; #100;
A = 16'h0051; B = 16'h0068; #100;
A = 16'h0051; B = 16'h0069; #100;
A = 16'h0051; B = 16'h006A; #100;
A = 16'h0051; B = 16'h006B; #100;
A = 16'h0051; B = 16'h006C; #100;
A = 16'h0051; B = 16'h006D; #100;
A = 16'h0051; B = 16'h006E; #100;
A = 16'h0051; B = 16'h006F; #100;
A = 16'h0051; B = 16'h0070; #100;
A = 16'h0051; B = 16'h0071; #100;
A = 16'h0051; B = 16'h0072; #100;
A = 16'h0051; B = 16'h0073; #100;
A = 16'h0051; B = 16'h0074; #100;
A = 16'h0051; B = 16'h0075; #100;
A = 16'h0051; B = 16'h0076; #100;
A = 16'h0051; B = 16'h0077; #100;
A = 16'h0051; B = 16'h0078; #100;
A = 16'h0051; B = 16'h0079; #100;
A = 16'h0051; B = 16'h007A; #100;
A = 16'h0051; B = 16'h007B; #100;
A = 16'h0051; B = 16'h007C; #100;
A = 16'h0051; B = 16'h007D; #100;
A = 16'h0051; B = 16'h007E; #100;
A = 16'h0051; B = 16'h007F; #100;
A = 16'h0051; B = 16'h0080; #100;
A = 16'h0051; B = 16'h0081; #100;
A = 16'h0051; B = 16'h0082; #100;
A = 16'h0051; B = 16'h0083; #100;
A = 16'h0051; B = 16'h0084; #100;
A = 16'h0051; B = 16'h0085; #100;
A = 16'h0051; B = 16'h0086; #100;
A = 16'h0051; B = 16'h0087; #100;
A = 16'h0051; B = 16'h0088; #100;
A = 16'h0051; B = 16'h0089; #100;
A = 16'h0051; B = 16'h008A; #100;
A = 16'h0051; B = 16'h008B; #100;
A = 16'h0051; B = 16'h008C; #100;
A = 16'h0051; B = 16'h008D; #100;
A = 16'h0051; B = 16'h008E; #100;
A = 16'h0051; B = 16'h008F; #100;
A = 16'h0051; B = 16'h0090; #100;
A = 16'h0051; B = 16'h0091; #100;
A = 16'h0051; B = 16'h0092; #100;
A = 16'h0051; B = 16'h0093; #100;
A = 16'h0051; B = 16'h0094; #100;
A = 16'h0051; B = 16'h0095; #100;
A = 16'h0051; B = 16'h0096; #100;
A = 16'h0051; B = 16'h0097; #100;
A = 16'h0051; B = 16'h0098; #100;
A = 16'h0051; B = 16'h0099; #100;
A = 16'h0051; B = 16'h009A; #100;
A = 16'h0051; B = 16'h009B; #100;
A = 16'h0051; B = 16'h009C; #100;
A = 16'h0051; B = 16'h009D; #100;
A = 16'h0051; B = 16'h009E; #100;
A = 16'h0051; B = 16'h009F; #100;
A = 16'h0051; B = 16'h00A0; #100;
A = 16'h0051; B = 16'h00A1; #100;
A = 16'h0051; B = 16'h00A2; #100;
A = 16'h0051; B = 16'h00A3; #100;
A = 16'h0051; B = 16'h00A4; #100;
A = 16'h0051; B = 16'h00A5; #100;
A = 16'h0051; B = 16'h00A6; #100;
A = 16'h0051; B = 16'h00A7; #100;
A = 16'h0051; B = 16'h00A8; #100;
A = 16'h0051; B = 16'h00A9; #100;
A = 16'h0051; B = 16'h00AA; #100;
A = 16'h0051; B = 16'h00AB; #100;
A = 16'h0051; B = 16'h00AC; #100;
A = 16'h0051; B = 16'h00AD; #100;
A = 16'h0051; B = 16'h00AE; #100;
A = 16'h0051; B = 16'h00AF; #100;
A = 16'h0051; B = 16'h00B0; #100;
A = 16'h0051; B = 16'h00B1; #100;
A = 16'h0051; B = 16'h00B2; #100;
A = 16'h0051; B = 16'h00B3; #100;
A = 16'h0051; B = 16'h00B4; #100;
A = 16'h0051; B = 16'h00B5; #100;
A = 16'h0051; B = 16'h00B6; #100;
A = 16'h0051; B = 16'h00B7; #100;
A = 16'h0051; B = 16'h00B8; #100;
A = 16'h0051; B = 16'h00B9; #100;
A = 16'h0051; B = 16'h00BA; #100;
A = 16'h0051; B = 16'h00BB; #100;
A = 16'h0051; B = 16'h00BC; #100;
A = 16'h0051; B = 16'h00BD; #100;
A = 16'h0051; B = 16'h00BE; #100;
A = 16'h0051; B = 16'h00BF; #100;
A = 16'h0051; B = 16'h00C0; #100;
A = 16'h0051; B = 16'h00C1; #100;
A = 16'h0051; B = 16'h00C2; #100;
A = 16'h0051; B = 16'h00C3; #100;
A = 16'h0051; B = 16'h00C4; #100;
A = 16'h0051; B = 16'h00C5; #100;
A = 16'h0051; B = 16'h00C6; #100;
A = 16'h0051; B = 16'h00C7; #100;
A = 16'h0051; B = 16'h00C8; #100;
A = 16'h0051; B = 16'h00C9; #100;
A = 16'h0051; B = 16'h00CA; #100;
A = 16'h0051; B = 16'h00CB; #100;
A = 16'h0051; B = 16'h00CC; #100;
A = 16'h0051; B = 16'h00CD; #100;
A = 16'h0051; B = 16'h00CE; #100;
A = 16'h0051; B = 16'h00CF; #100;
A = 16'h0051; B = 16'h00D0; #100;
A = 16'h0051; B = 16'h00D1; #100;
A = 16'h0051; B = 16'h00D2; #100;
A = 16'h0051; B = 16'h00D3; #100;
A = 16'h0051; B = 16'h00D4; #100;
A = 16'h0051; B = 16'h00D5; #100;
A = 16'h0051; B = 16'h00D6; #100;
A = 16'h0051; B = 16'h00D7; #100;
A = 16'h0051; B = 16'h00D8; #100;
A = 16'h0051; B = 16'h00D9; #100;
A = 16'h0051; B = 16'h00DA; #100;
A = 16'h0051; B = 16'h00DB; #100;
A = 16'h0051; B = 16'h00DC; #100;
A = 16'h0051; B = 16'h00DD; #100;
A = 16'h0051; B = 16'h00DE; #100;
A = 16'h0051; B = 16'h00DF; #100;
A = 16'h0051; B = 16'h00E0; #100;
A = 16'h0051; B = 16'h00E1; #100;
A = 16'h0051; B = 16'h00E2; #100;
A = 16'h0051; B = 16'h00E3; #100;
A = 16'h0051; B = 16'h00E4; #100;
A = 16'h0051; B = 16'h00E5; #100;
A = 16'h0051; B = 16'h00E6; #100;
A = 16'h0051; B = 16'h00E7; #100;
A = 16'h0051; B = 16'h00E8; #100;
A = 16'h0051; B = 16'h00E9; #100;
A = 16'h0051; B = 16'h00EA; #100;
A = 16'h0051; B = 16'h00EB; #100;
A = 16'h0051; B = 16'h00EC; #100;
A = 16'h0051; B = 16'h00ED; #100;
A = 16'h0051; B = 16'h00EE; #100;
A = 16'h0051; B = 16'h00EF; #100;
A = 16'h0051; B = 16'h00F0; #100;
A = 16'h0051; B = 16'h00F1; #100;
A = 16'h0051; B = 16'h00F2; #100;
A = 16'h0051; B = 16'h00F3; #100;
A = 16'h0051; B = 16'h00F4; #100;
A = 16'h0051; B = 16'h00F5; #100;
A = 16'h0051; B = 16'h00F6; #100;
A = 16'h0051; B = 16'h00F7; #100;
A = 16'h0051; B = 16'h00F8; #100;
A = 16'h0051; B = 16'h00F9; #100;
A = 16'h0051; B = 16'h00FA; #100;
A = 16'h0051; B = 16'h00FB; #100;
A = 16'h0051; B = 16'h00FC; #100;
A = 16'h0051; B = 16'h00FD; #100;
A = 16'h0051; B = 16'h00FE; #100;
A = 16'h0051; B = 16'h00FF; #100;
A = 16'h0052; B = 16'h000; #100;
A = 16'h0052; B = 16'h001; #100;
A = 16'h0052; B = 16'h002; #100;
A = 16'h0052; B = 16'h003; #100;
A = 16'h0052; B = 16'h004; #100;
A = 16'h0052; B = 16'h005; #100;
A = 16'h0052; B = 16'h006; #100;
A = 16'h0052; B = 16'h007; #100;
A = 16'h0052; B = 16'h008; #100;
A = 16'h0052; B = 16'h009; #100;
A = 16'h0052; B = 16'h00A; #100;
A = 16'h0052; B = 16'h00B; #100;
A = 16'h0052; B = 16'h00C; #100;
A = 16'h0052; B = 16'h00D; #100;
A = 16'h0052; B = 16'h00E; #100;
A = 16'h0052; B = 16'h00F; #100;
A = 16'h0052; B = 16'h0010; #100;
A = 16'h0052; B = 16'h0011; #100;
A = 16'h0052; B = 16'h0012; #100;
A = 16'h0052; B = 16'h0013; #100;
A = 16'h0052; B = 16'h0014; #100;
A = 16'h0052; B = 16'h0015; #100;
A = 16'h0052; B = 16'h0016; #100;
A = 16'h0052; B = 16'h0017; #100;
A = 16'h0052; B = 16'h0018; #100;
A = 16'h0052; B = 16'h0019; #100;
A = 16'h0052; B = 16'h001A; #100;
A = 16'h0052; B = 16'h001B; #100;
A = 16'h0052; B = 16'h001C; #100;
A = 16'h0052; B = 16'h001D; #100;
A = 16'h0052; B = 16'h001E; #100;
A = 16'h0052; B = 16'h001F; #100;
A = 16'h0052; B = 16'h0020; #100;
A = 16'h0052; B = 16'h0021; #100;
A = 16'h0052; B = 16'h0022; #100;
A = 16'h0052; B = 16'h0023; #100;
A = 16'h0052; B = 16'h0024; #100;
A = 16'h0052; B = 16'h0025; #100;
A = 16'h0052; B = 16'h0026; #100;
A = 16'h0052; B = 16'h0027; #100;
A = 16'h0052; B = 16'h0028; #100;
A = 16'h0052; B = 16'h0029; #100;
A = 16'h0052; B = 16'h002A; #100;
A = 16'h0052; B = 16'h002B; #100;
A = 16'h0052; B = 16'h002C; #100;
A = 16'h0052; B = 16'h002D; #100;
A = 16'h0052; B = 16'h002E; #100;
A = 16'h0052; B = 16'h002F; #100;
A = 16'h0052; B = 16'h0030; #100;
A = 16'h0052; B = 16'h0031; #100;
A = 16'h0052; B = 16'h0032; #100;
A = 16'h0052; B = 16'h0033; #100;
A = 16'h0052; B = 16'h0034; #100;
A = 16'h0052; B = 16'h0035; #100;
A = 16'h0052; B = 16'h0036; #100;
A = 16'h0052; B = 16'h0037; #100;
A = 16'h0052; B = 16'h0038; #100;
A = 16'h0052; B = 16'h0039; #100;
A = 16'h0052; B = 16'h003A; #100;
A = 16'h0052; B = 16'h003B; #100;
A = 16'h0052; B = 16'h003C; #100;
A = 16'h0052; B = 16'h003D; #100;
A = 16'h0052; B = 16'h003E; #100;
A = 16'h0052; B = 16'h003F; #100;
A = 16'h0052; B = 16'h0040; #100;
A = 16'h0052; B = 16'h0041; #100;
A = 16'h0052; B = 16'h0042; #100;
A = 16'h0052; B = 16'h0043; #100;
A = 16'h0052; B = 16'h0044; #100;
A = 16'h0052; B = 16'h0045; #100;
A = 16'h0052; B = 16'h0046; #100;
A = 16'h0052; B = 16'h0047; #100;
A = 16'h0052; B = 16'h0048; #100;
A = 16'h0052; B = 16'h0049; #100;
A = 16'h0052; B = 16'h004A; #100;
A = 16'h0052; B = 16'h004B; #100;
A = 16'h0052; B = 16'h004C; #100;
A = 16'h0052; B = 16'h004D; #100;
A = 16'h0052; B = 16'h004E; #100;
A = 16'h0052; B = 16'h004F; #100;
A = 16'h0052; B = 16'h0050; #100;
A = 16'h0052; B = 16'h0051; #100;
A = 16'h0052; B = 16'h0052; #100;
A = 16'h0052; B = 16'h0053; #100;
A = 16'h0052; B = 16'h0054; #100;
A = 16'h0052; B = 16'h0055; #100;
A = 16'h0052; B = 16'h0056; #100;
A = 16'h0052; B = 16'h0057; #100;
A = 16'h0052; B = 16'h0058; #100;
A = 16'h0052; B = 16'h0059; #100;
A = 16'h0052; B = 16'h005A; #100;
A = 16'h0052; B = 16'h005B; #100;
A = 16'h0052; B = 16'h005C; #100;
A = 16'h0052; B = 16'h005D; #100;
A = 16'h0052; B = 16'h005E; #100;
A = 16'h0052; B = 16'h005F; #100;
A = 16'h0052; B = 16'h0060; #100;
A = 16'h0052; B = 16'h0061; #100;
A = 16'h0052; B = 16'h0062; #100;
A = 16'h0052; B = 16'h0063; #100;
A = 16'h0052; B = 16'h0064; #100;
A = 16'h0052; B = 16'h0065; #100;
A = 16'h0052; B = 16'h0066; #100;
A = 16'h0052; B = 16'h0067; #100;
A = 16'h0052; B = 16'h0068; #100;
A = 16'h0052; B = 16'h0069; #100;
A = 16'h0052; B = 16'h006A; #100;
A = 16'h0052; B = 16'h006B; #100;
A = 16'h0052; B = 16'h006C; #100;
A = 16'h0052; B = 16'h006D; #100;
A = 16'h0052; B = 16'h006E; #100;
A = 16'h0052; B = 16'h006F; #100;
A = 16'h0052; B = 16'h0070; #100;
A = 16'h0052; B = 16'h0071; #100;
A = 16'h0052; B = 16'h0072; #100;
A = 16'h0052; B = 16'h0073; #100;
A = 16'h0052; B = 16'h0074; #100;
A = 16'h0052; B = 16'h0075; #100;
A = 16'h0052; B = 16'h0076; #100;
A = 16'h0052; B = 16'h0077; #100;
A = 16'h0052; B = 16'h0078; #100;
A = 16'h0052; B = 16'h0079; #100;
A = 16'h0052; B = 16'h007A; #100;
A = 16'h0052; B = 16'h007B; #100;
A = 16'h0052; B = 16'h007C; #100;
A = 16'h0052; B = 16'h007D; #100;
A = 16'h0052; B = 16'h007E; #100;
A = 16'h0052; B = 16'h007F; #100;
A = 16'h0052; B = 16'h0080; #100;
A = 16'h0052; B = 16'h0081; #100;
A = 16'h0052; B = 16'h0082; #100;
A = 16'h0052; B = 16'h0083; #100;
A = 16'h0052; B = 16'h0084; #100;
A = 16'h0052; B = 16'h0085; #100;
A = 16'h0052; B = 16'h0086; #100;
A = 16'h0052; B = 16'h0087; #100;
A = 16'h0052; B = 16'h0088; #100;
A = 16'h0052; B = 16'h0089; #100;
A = 16'h0052; B = 16'h008A; #100;
A = 16'h0052; B = 16'h008B; #100;
A = 16'h0052; B = 16'h008C; #100;
A = 16'h0052; B = 16'h008D; #100;
A = 16'h0052; B = 16'h008E; #100;
A = 16'h0052; B = 16'h008F; #100;
A = 16'h0052; B = 16'h0090; #100;
A = 16'h0052; B = 16'h0091; #100;
A = 16'h0052; B = 16'h0092; #100;
A = 16'h0052; B = 16'h0093; #100;
A = 16'h0052; B = 16'h0094; #100;
A = 16'h0052; B = 16'h0095; #100;
A = 16'h0052; B = 16'h0096; #100;
A = 16'h0052; B = 16'h0097; #100;
A = 16'h0052; B = 16'h0098; #100;
A = 16'h0052; B = 16'h0099; #100;
A = 16'h0052; B = 16'h009A; #100;
A = 16'h0052; B = 16'h009B; #100;
A = 16'h0052; B = 16'h009C; #100;
A = 16'h0052; B = 16'h009D; #100;
A = 16'h0052; B = 16'h009E; #100;
A = 16'h0052; B = 16'h009F; #100;
A = 16'h0052; B = 16'h00A0; #100;
A = 16'h0052; B = 16'h00A1; #100;
A = 16'h0052; B = 16'h00A2; #100;
A = 16'h0052; B = 16'h00A3; #100;
A = 16'h0052; B = 16'h00A4; #100;
A = 16'h0052; B = 16'h00A5; #100;
A = 16'h0052; B = 16'h00A6; #100;
A = 16'h0052; B = 16'h00A7; #100;
A = 16'h0052; B = 16'h00A8; #100;
A = 16'h0052; B = 16'h00A9; #100;
A = 16'h0052; B = 16'h00AA; #100;
A = 16'h0052; B = 16'h00AB; #100;
A = 16'h0052; B = 16'h00AC; #100;
A = 16'h0052; B = 16'h00AD; #100;
A = 16'h0052; B = 16'h00AE; #100;
A = 16'h0052; B = 16'h00AF; #100;
A = 16'h0052; B = 16'h00B0; #100;
A = 16'h0052; B = 16'h00B1; #100;
A = 16'h0052; B = 16'h00B2; #100;
A = 16'h0052; B = 16'h00B3; #100;
A = 16'h0052; B = 16'h00B4; #100;
A = 16'h0052; B = 16'h00B5; #100;
A = 16'h0052; B = 16'h00B6; #100;
A = 16'h0052; B = 16'h00B7; #100;
A = 16'h0052; B = 16'h00B8; #100;
A = 16'h0052; B = 16'h00B9; #100;
A = 16'h0052; B = 16'h00BA; #100;
A = 16'h0052; B = 16'h00BB; #100;
A = 16'h0052; B = 16'h00BC; #100;
A = 16'h0052; B = 16'h00BD; #100;
A = 16'h0052; B = 16'h00BE; #100;
A = 16'h0052; B = 16'h00BF; #100;
A = 16'h0052; B = 16'h00C0; #100;
A = 16'h0052; B = 16'h00C1; #100;
A = 16'h0052; B = 16'h00C2; #100;
A = 16'h0052; B = 16'h00C3; #100;
A = 16'h0052; B = 16'h00C4; #100;
A = 16'h0052; B = 16'h00C5; #100;
A = 16'h0052; B = 16'h00C6; #100;
A = 16'h0052; B = 16'h00C7; #100;
A = 16'h0052; B = 16'h00C8; #100;
A = 16'h0052; B = 16'h00C9; #100;
A = 16'h0052; B = 16'h00CA; #100;
A = 16'h0052; B = 16'h00CB; #100;
A = 16'h0052; B = 16'h00CC; #100;
A = 16'h0052; B = 16'h00CD; #100;
A = 16'h0052; B = 16'h00CE; #100;
A = 16'h0052; B = 16'h00CF; #100;
A = 16'h0052; B = 16'h00D0; #100;
A = 16'h0052; B = 16'h00D1; #100;
A = 16'h0052; B = 16'h00D2; #100;
A = 16'h0052; B = 16'h00D3; #100;
A = 16'h0052; B = 16'h00D4; #100;
A = 16'h0052; B = 16'h00D5; #100;
A = 16'h0052; B = 16'h00D6; #100;
A = 16'h0052; B = 16'h00D7; #100;
A = 16'h0052; B = 16'h00D8; #100;
A = 16'h0052; B = 16'h00D9; #100;
A = 16'h0052; B = 16'h00DA; #100;
A = 16'h0052; B = 16'h00DB; #100;
A = 16'h0052; B = 16'h00DC; #100;
A = 16'h0052; B = 16'h00DD; #100;
A = 16'h0052; B = 16'h00DE; #100;
A = 16'h0052; B = 16'h00DF; #100;
A = 16'h0052; B = 16'h00E0; #100;
A = 16'h0052; B = 16'h00E1; #100;
A = 16'h0052; B = 16'h00E2; #100;
A = 16'h0052; B = 16'h00E3; #100;
A = 16'h0052; B = 16'h00E4; #100;
A = 16'h0052; B = 16'h00E5; #100;
A = 16'h0052; B = 16'h00E6; #100;
A = 16'h0052; B = 16'h00E7; #100;
A = 16'h0052; B = 16'h00E8; #100;
A = 16'h0052; B = 16'h00E9; #100;
A = 16'h0052; B = 16'h00EA; #100;
A = 16'h0052; B = 16'h00EB; #100;
A = 16'h0052; B = 16'h00EC; #100;
A = 16'h0052; B = 16'h00ED; #100;
A = 16'h0052; B = 16'h00EE; #100;
A = 16'h0052; B = 16'h00EF; #100;
A = 16'h0052; B = 16'h00F0; #100;
A = 16'h0052; B = 16'h00F1; #100;
A = 16'h0052; B = 16'h00F2; #100;
A = 16'h0052; B = 16'h00F3; #100;
A = 16'h0052; B = 16'h00F4; #100;
A = 16'h0052; B = 16'h00F5; #100;
A = 16'h0052; B = 16'h00F6; #100;
A = 16'h0052; B = 16'h00F7; #100;
A = 16'h0052; B = 16'h00F8; #100;
A = 16'h0052; B = 16'h00F9; #100;
A = 16'h0052; B = 16'h00FA; #100;
A = 16'h0052; B = 16'h00FB; #100;
A = 16'h0052; B = 16'h00FC; #100;
A = 16'h0052; B = 16'h00FD; #100;
A = 16'h0052; B = 16'h00FE; #100;
A = 16'h0052; B = 16'h00FF; #100;
A = 16'h0053; B = 16'h000; #100;
A = 16'h0053; B = 16'h001; #100;
A = 16'h0053; B = 16'h002; #100;
A = 16'h0053; B = 16'h003; #100;
A = 16'h0053; B = 16'h004; #100;
A = 16'h0053; B = 16'h005; #100;
A = 16'h0053; B = 16'h006; #100;
A = 16'h0053; B = 16'h007; #100;
A = 16'h0053; B = 16'h008; #100;
A = 16'h0053; B = 16'h009; #100;
A = 16'h0053; B = 16'h00A; #100;
A = 16'h0053; B = 16'h00B; #100;
A = 16'h0053; B = 16'h00C; #100;
A = 16'h0053; B = 16'h00D; #100;
A = 16'h0053; B = 16'h00E; #100;
A = 16'h0053; B = 16'h00F; #100;
A = 16'h0053; B = 16'h0010; #100;
A = 16'h0053; B = 16'h0011; #100;
A = 16'h0053; B = 16'h0012; #100;
A = 16'h0053; B = 16'h0013; #100;
A = 16'h0053; B = 16'h0014; #100;
A = 16'h0053; B = 16'h0015; #100;
A = 16'h0053; B = 16'h0016; #100;
A = 16'h0053; B = 16'h0017; #100;
A = 16'h0053; B = 16'h0018; #100;
A = 16'h0053; B = 16'h0019; #100;
A = 16'h0053; B = 16'h001A; #100;
A = 16'h0053; B = 16'h001B; #100;
A = 16'h0053; B = 16'h001C; #100;
A = 16'h0053; B = 16'h001D; #100;
A = 16'h0053; B = 16'h001E; #100;
A = 16'h0053; B = 16'h001F; #100;
A = 16'h0053; B = 16'h0020; #100;
A = 16'h0053; B = 16'h0021; #100;
A = 16'h0053; B = 16'h0022; #100;
A = 16'h0053; B = 16'h0023; #100;
A = 16'h0053; B = 16'h0024; #100;
A = 16'h0053; B = 16'h0025; #100;
A = 16'h0053; B = 16'h0026; #100;
A = 16'h0053; B = 16'h0027; #100;
A = 16'h0053; B = 16'h0028; #100;
A = 16'h0053; B = 16'h0029; #100;
A = 16'h0053; B = 16'h002A; #100;
A = 16'h0053; B = 16'h002B; #100;
A = 16'h0053; B = 16'h002C; #100;
A = 16'h0053; B = 16'h002D; #100;
A = 16'h0053; B = 16'h002E; #100;
A = 16'h0053; B = 16'h002F; #100;
A = 16'h0053; B = 16'h0030; #100;
A = 16'h0053; B = 16'h0031; #100;
A = 16'h0053; B = 16'h0032; #100;
A = 16'h0053; B = 16'h0033; #100;
A = 16'h0053; B = 16'h0034; #100;
A = 16'h0053; B = 16'h0035; #100;
A = 16'h0053; B = 16'h0036; #100;
A = 16'h0053; B = 16'h0037; #100;
A = 16'h0053; B = 16'h0038; #100;
A = 16'h0053; B = 16'h0039; #100;
A = 16'h0053; B = 16'h003A; #100;
A = 16'h0053; B = 16'h003B; #100;
A = 16'h0053; B = 16'h003C; #100;
A = 16'h0053; B = 16'h003D; #100;
A = 16'h0053; B = 16'h003E; #100;
A = 16'h0053; B = 16'h003F; #100;
A = 16'h0053; B = 16'h0040; #100;
A = 16'h0053; B = 16'h0041; #100;
A = 16'h0053; B = 16'h0042; #100;
A = 16'h0053; B = 16'h0043; #100;
A = 16'h0053; B = 16'h0044; #100;
A = 16'h0053; B = 16'h0045; #100;
A = 16'h0053; B = 16'h0046; #100;
A = 16'h0053; B = 16'h0047; #100;
A = 16'h0053; B = 16'h0048; #100;
A = 16'h0053; B = 16'h0049; #100;
A = 16'h0053; B = 16'h004A; #100;
A = 16'h0053; B = 16'h004B; #100;
A = 16'h0053; B = 16'h004C; #100;
A = 16'h0053; B = 16'h004D; #100;
A = 16'h0053; B = 16'h004E; #100;
A = 16'h0053; B = 16'h004F; #100;
A = 16'h0053; B = 16'h0050; #100;
A = 16'h0053; B = 16'h0051; #100;
A = 16'h0053; B = 16'h0052; #100;
A = 16'h0053; B = 16'h0053; #100;
A = 16'h0053; B = 16'h0054; #100;
A = 16'h0053; B = 16'h0055; #100;
A = 16'h0053; B = 16'h0056; #100;
A = 16'h0053; B = 16'h0057; #100;
A = 16'h0053; B = 16'h0058; #100;
A = 16'h0053; B = 16'h0059; #100;
A = 16'h0053; B = 16'h005A; #100;
A = 16'h0053; B = 16'h005B; #100;
A = 16'h0053; B = 16'h005C; #100;
A = 16'h0053; B = 16'h005D; #100;
A = 16'h0053; B = 16'h005E; #100;
A = 16'h0053; B = 16'h005F; #100;
A = 16'h0053; B = 16'h0060; #100;
A = 16'h0053; B = 16'h0061; #100;
A = 16'h0053; B = 16'h0062; #100;
A = 16'h0053; B = 16'h0063; #100;
A = 16'h0053; B = 16'h0064; #100;
A = 16'h0053; B = 16'h0065; #100;
A = 16'h0053; B = 16'h0066; #100;
A = 16'h0053; B = 16'h0067; #100;
A = 16'h0053; B = 16'h0068; #100;
A = 16'h0053; B = 16'h0069; #100;
A = 16'h0053; B = 16'h006A; #100;
A = 16'h0053; B = 16'h006B; #100;
A = 16'h0053; B = 16'h006C; #100;
A = 16'h0053; B = 16'h006D; #100;
A = 16'h0053; B = 16'h006E; #100;
A = 16'h0053; B = 16'h006F; #100;
A = 16'h0053; B = 16'h0070; #100;
A = 16'h0053; B = 16'h0071; #100;
A = 16'h0053; B = 16'h0072; #100;
A = 16'h0053; B = 16'h0073; #100;
A = 16'h0053; B = 16'h0074; #100;
A = 16'h0053; B = 16'h0075; #100;
A = 16'h0053; B = 16'h0076; #100;
A = 16'h0053; B = 16'h0077; #100;
A = 16'h0053; B = 16'h0078; #100;
A = 16'h0053; B = 16'h0079; #100;
A = 16'h0053; B = 16'h007A; #100;
A = 16'h0053; B = 16'h007B; #100;
A = 16'h0053; B = 16'h007C; #100;
A = 16'h0053; B = 16'h007D; #100;
A = 16'h0053; B = 16'h007E; #100;
A = 16'h0053; B = 16'h007F; #100;
A = 16'h0053; B = 16'h0080; #100;
A = 16'h0053; B = 16'h0081; #100;
A = 16'h0053; B = 16'h0082; #100;
A = 16'h0053; B = 16'h0083; #100;
A = 16'h0053; B = 16'h0084; #100;
A = 16'h0053; B = 16'h0085; #100;
A = 16'h0053; B = 16'h0086; #100;
A = 16'h0053; B = 16'h0087; #100;
A = 16'h0053; B = 16'h0088; #100;
A = 16'h0053; B = 16'h0089; #100;
A = 16'h0053; B = 16'h008A; #100;
A = 16'h0053; B = 16'h008B; #100;
A = 16'h0053; B = 16'h008C; #100;
A = 16'h0053; B = 16'h008D; #100;
A = 16'h0053; B = 16'h008E; #100;
A = 16'h0053; B = 16'h008F; #100;
A = 16'h0053; B = 16'h0090; #100;
A = 16'h0053; B = 16'h0091; #100;
A = 16'h0053; B = 16'h0092; #100;
A = 16'h0053; B = 16'h0093; #100;
A = 16'h0053; B = 16'h0094; #100;
A = 16'h0053; B = 16'h0095; #100;
A = 16'h0053; B = 16'h0096; #100;
A = 16'h0053; B = 16'h0097; #100;
A = 16'h0053; B = 16'h0098; #100;
A = 16'h0053; B = 16'h0099; #100;
A = 16'h0053; B = 16'h009A; #100;
A = 16'h0053; B = 16'h009B; #100;
A = 16'h0053; B = 16'h009C; #100;
A = 16'h0053; B = 16'h009D; #100;
A = 16'h0053; B = 16'h009E; #100;
A = 16'h0053; B = 16'h009F; #100;
A = 16'h0053; B = 16'h00A0; #100;
A = 16'h0053; B = 16'h00A1; #100;
A = 16'h0053; B = 16'h00A2; #100;
A = 16'h0053; B = 16'h00A3; #100;
A = 16'h0053; B = 16'h00A4; #100;
A = 16'h0053; B = 16'h00A5; #100;
A = 16'h0053; B = 16'h00A6; #100;
A = 16'h0053; B = 16'h00A7; #100;
A = 16'h0053; B = 16'h00A8; #100;
A = 16'h0053; B = 16'h00A9; #100;
A = 16'h0053; B = 16'h00AA; #100;
A = 16'h0053; B = 16'h00AB; #100;
A = 16'h0053; B = 16'h00AC; #100;
A = 16'h0053; B = 16'h00AD; #100;
A = 16'h0053; B = 16'h00AE; #100;
A = 16'h0053; B = 16'h00AF; #100;
A = 16'h0053; B = 16'h00B0; #100;
A = 16'h0053; B = 16'h00B1; #100;
A = 16'h0053; B = 16'h00B2; #100;
A = 16'h0053; B = 16'h00B3; #100;
A = 16'h0053; B = 16'h00B4; #100;
A = 16'h0053; B = 16'h00B5; #100;
A = 16'h0053; B = 16'h00B6; #100;
A = 16'h0053; B = 16'h00B7; #100;
A = 16'h0053; B = 16'h00B8; #100;
A = 16'h0053; B = 16'h00B9; #100;
A = 16'h0053; B = 16'h00BA; #100;
A = 16'h0053; B = 16'h00BB; #100;
A = 16'h0053; B = 16'h00BC; #100;
A = 16'h0053; B = 16'h00BD; #100;
A = 16'h0053; B = 16'h00BE; #100;
A = 16'h0053; B = 16'h00BF; #100;
A = 16'h0053; B = 16'h00C0; #100;
A = 16'h0053; B = 16'h00C1; #100;
A = 16'h0053; B = 16'h00C2; #100;
A = 16'h0053; B = 16'h00C3; #100;
A = 16'h0053; B = 16'h00C4; #100;
A = 16'h0053; B = 16'h00C5; #100;
A = 16'h0053; B = 16'h00C6; #100;
A = 16'h0053; B = 16'h00C7; #100;
A = 16'h0053; B = 16'h00C8; #100;
A = 16'h0053; B = 16'h00C9; #100;
A = 16'h0053; B = 16'h00CA; #100;
A = 16'h0053; B = 16'h00CB; #100;
A = 16'h0053; B = 16'h00CC; #100;
A = 16'h0053; B = 16'h00CD; #100;
A = 16'h0053; B = 16'h00CE; #100;
A = 16'h0053; B = 16'h00CF; #100;
A = 16'h0053; B = 16'h00D0; #100;
A = 16'h0053; B = 16'h00D1; #100;
A = 16'h0053; B = 16'h00D2; #100;
A = 16'h0053; B = 16'h00D3; #100;
A = 16'h0053; B = 16'h00D4; #100;
A = 16'h0053; B = 16'h00D5; #100;
A = 16'h0053; B = 16'h00D6; #100;
A = 16'h0053; B = 16'h00D7; #100;
A = 16'h0053; B = 16'h00D8; #100;
A = 16'h0053; B = 16'h00D9; #100;
A = 16'h0053; B = 16'h00DA; #100;
A = 16'h0053; B = 16'h00DB; #100;
A = 16'h0053; B = 16'h00DC; #100;
A = 16'h0053; B = 16'h00DD; #100;
A = 16'h0053; B = 16'h00DE; #100;
A = 16'h0053; B = 16'h00DF; #100;
A = 16'h0053; B = 16'h00E0; #100;
A = 16'h0053; B = 16'h00E1; #100;
A = 16'h0053; B = 16'h00E2; #100;
A = 16'h0053; B = 16'h00E3; #100;
A = 16'h0053; B = 16'h00E4; #100;
A = 16'h0053; B = 16'h00E5; #100;
A = 16'h0053; B = 16'h00E6; #100;
A = 16'h0053; B = 16'h00E7; #100;
A = 16'h0053; B = 16'h00E8; #100;
A = 16'h0053; B = 16'h00E9; #100;
A = 16'h0053; B = 16'h00EA; #100;
A = 16'h0053; B = 16'h00EB; #100;
A = 16'h0053; B = 16'h00EC; #100;
A = 16'h0053; B = 16'h00ED; #100;
A = 16'h0053; B = 16'h00EE; #100;
A = 16'h0053; B = 16'h00EF; #100;
A = 16'h0053; B = 16'h00F0; #100;
A = 16'h0053; B = 16'h00F1; #100;
A = 16'h0053; B = 16'h00F2; #100;
A = 16'h0053; B = 16'h00F3; #100;
A = 16'h0053; B = 16'h00F4; #100;
A = 16'h0053; B = 16'h00F5; #100;
A = 16'h0053; B = 16'h00F6; #100;
A = 16'h0053; B = 16'h00F7; #100;
A = 16'h0053; B = 16'h00F8; #100;
A = 16'h0053; B = 16'h00F9; #100;
A = 16'h0053; B = 16'h00FA; #100;
A = 16'h0053; B = 16'h00FB; #100;
A = 16'h0053; B = 16'h00FC; #100;
A = 16'h0053; B = 16'h00FD; #100;
A = 16'h0053; B = 16'h00FE; #100;
A = 16'h0053; B = 16'h00FF; #100;
A = 16'h0054; B = 16'h000; #100;
A = 16'h0054; B = 16'h001; #100;
A = 16'h0054; B = 16'h002; #100;
A = 16'h0054; B = 16'h003; #100;
A = 16'h0054; B = 16'h004; #100;
A = 16'h0054; B = 16'h005; #100;
A = 16'h0054; B = 16'h006; #100;
A = 16'h0054; B = 16'h007; #100;
A = 16'h0054; B = 16'h008; #100;
A = 16'h0054; B = 16'h009; #100;
A = 16'h0054; B = 16'h00A; #100;
A = 16'h0054; B = 16'h00B; #100;
A = 16'h0054; B = 16'h00C; #100;
A = 16'h0054; B = 16'h00D; #100;
A = 16'h0054; B = 16'h00E; #100;
A = 16'h0054; B = 16'h00F; #100;
A = 16'h0054; B = 16'h0010; #100;
A = 16'h0054; B = 16'h0011; #100;
A = 16'h0054; B = 16'h0012; #100;
A = 16'h0054; B = 16'h0013; #100;
A = 16'h0054; B = 16'h0014; #100;
A = 16'h0054; B = 16'h0015; #100;
A = 16'h0054; B = 16'h0016; #100;
A = 16'h0054; B = 16'h0017; #100;
A = 16'h0054; B = 16'h0018; #100;
A = 16'h0054; B = 16'h0019; #100;
A = 16'h0054; B = 16'h001A; #100;
A = 16'h0054; B = 16'h001B; #100;
A = 16'h0054; B = 16'h001C; #100;
A = 16'h0054; B = 16'h001D; #100;
A = 16'h0054; B = 16'h001E; #100;
A = 16'h0054; B = 16'h001F; #100;
A = 16'h0054; B = 16'h0020; #100;
A = 16'h0054; B = 16'h0021; #100;
A = 16'h0054; B = 16'h0022; #100;
A = 16'h0054; B = 16'h0023; #100;
A = 16'h0054; B = 16'h0024; #100;
A = 16'h0054; B = 16'h0025; #100;
A = 16'h0054; B = 16'h0026; #100;
A = 16'h0054; B = 16'h0027; #100;
A = 16'h0054; B = 16'h0028; #100;
A = 16'h0054; B = 16'h0029; #100;
A = 16'h0054; B = 16'h002A; #100;
A = 16'h0054; B = 16'h002B; #100;
A = 16'h0054; B = 16'h002C; #100;
A = 16'h0054; B = 16'h002D; #100;
A = 16'h0054; B = 16'h002E; #100;
A = 16'h0054; B = 16'h002F; #100;
A = 16'h0054; B = 16'h0030; #100;
A = 16'h0054; B = 16'h0031; #100;
A = 16'h0054; B = 16'h0032; #100;
A = 16'h0054; B = 16'h0033; #100;
A = 16'h0054; B = 16'h0034; #100;
A = 16'h0054; B = 16'h0035; #100;
A = 16'h0054; B = 16'h0036; #100;
A = 16'h0054; B = 16'h0037; #100;
A = 16'h0054; B = 16'h0038; #100;
A = 16'h0054; B = 16'h0039; #100;
A = 16'h0054; B = 16'h003A; #100;
A = 16'h0054; B = 16'h003B; #100;
A = 16'h0054; B = 16'h003C; #100;
A = 16'h0054; B = 16'h003D; #100;
A = 16'h0054; B = 16'h003E; #100;
A = 16'h0054; B = 16'h003F; #100;
A = 16'h0054; B = 16'h0040; #100;
A = 16'h0054; B = 16'h0041; #100;
A = 16'h0054; B = 16'h0042; #100;
A = 16'h0054; B = 16'h0043; #100;
A = 16'h0054; B = 16'h0044; #100;
A = 16'h0054; B = 16'h0045; #100;
A = 16'h0054; B = 16'h0046; #100;
A = 16'h0054; B = 16'h0047; #100;
A = 16'h0054; B = 16'h0048; #100;
A = 16'h0054; B = 16'h0049; #100;
A = 16'h0054; B = 16'h004A; #100;
A = 16'h0054; B = 16'h004B; #100;
A = 16'h0054; B = 16'h004C; #100;
A = 16'h0054; B = 16'h004D; #100;
A = 16'h0054; B = 16'h004E; #100;
A = 16'h0054; B = 16'h004F; #100;
A = 16'h0054; B = 16'h0050; #100;
A = 16'h0054; B = 16'h0051; #100;
A = 16'h0054; B = 16'h0052; #100;
A = 16'h0054; B = 16'h0053; #100;
A = 16'h0054; B = 16'h0054; #100;
A = 16'h0054; B = 16'h0055; #100;
A = 16'h0054; B = 16'h0056; #100;
A = 16'h0054; B = 16'h0057; #100;
A = 16'h0054; B = 16'h0058; #100;
A = 16'h0054; B = 16'h0059; #100;
A = 16'h0054; B = 16'h005A; #100;
A = 16'h0054; B = 16'h005B; #100;
A = 16'h0054; B = 16'h005C; #100;
A = 16'h0054; B = 16'h005D; #100;
A = 16'h0054; B = 16'h005E; #100;
A = 16'h0054; B = 16'h005F; #100;
A = 16'h0054; B = 16'h0060; #100;
A = 16'h0054; B = 16'h0061; #100;
A = 16'h0054; B = 16'h0062; #100;
A = 16'h0054; B = 16'h0063; #100;
A = 16'h0054; B = 16'h0064; #100;
A = 16'h0054; B = 16'h0065; #100;
A = 16'h0054; B = 16'h0066; #100;
A = 16'h0054; B = 16'h0067; #100;
A = 16'h0054; B = 16'h0068; #100;
A = 16'h0054; B = 16'h0069; #100;
A = 16'h0054; B = 16'h006A; #100;
A = 16'h0054; B = 16'h006B; #100;
A = 16'h0054; B = 16'h006C; #100;
A = 16'h0054; B = 16'h006D; #100;
A = 16'h0054; B = 16'h006E; #100;
A = 16'h0054; B = 16'h006F; #100;
A = 16'h0054; B = 16'h0070; #100;
A = 16'h0054; B = 16'h0071; #100;
A = 16'h0054; B = 16'h0072; #100;
A = 16'h0054; B = 16'h0073; #100;
A = 16'h0054; B = 16'h0074; #100;
A = 16'h0054; B = 16'h0075; #100;
A = 16'h0054; B = 16'h0076; #100;
A = 16'h0054; B = 16'h0077; #100;
A = 16'h0054; B = 16'h0078; #100;
A = 16'h0054; B = 16'h0079; #100;
A = 16'h0054; B = 16'h007A; #100;
A = 16'h0054; B = 16'h007B; #100;
A = 16'h0054; B = 16'h007C; #100;
A = 16'h0054; B = 16'h007D; #100;
A = 16'h0054; B = 16'h007E; #100;
A = 16'h0054; B = 16'h007F; #100;
A = 16'h0054; B = 16'h0080; #100;
A = 16'h0054; B = 16'h0081; #100;
A = 16'h0054; B = 16'h0082; #100;
A = 16'h0054; B = 16'h0083; #100;
A = 16'h0054; B = 16'h0084; #100;
A = 16'h0054; B = 16'h0085; #100;
A = 16'h0054; B = 16'h0086; #100;
A = 16'h0054; B = 16'h0087; #100;
A = 16'h0054; B = 16'h0088; #100;
A = 16'h0054; B = 16'h0089; #100;
A = 16'h0054; B = 16'h008A; #100;
A = 16'h0054; B = 16'h008B; #100;
A = 16'h0054; B = 16'h008C; #100;
A = 16'h0054; B = 16'h008D; #100;
A = 16'h0054; B = 16'h008E; #100;
A = 16'h0054; B = 16'h008F; #100;
A = 16'h0054; B = 16'h0090; #100;
A = 16'h0054; B = 16'h0091; #100;
A = 16'h0054; B = 16'h0092; #100;
A = 16'h0054; B = 16'h0093; #100;
A = 16'h0054; B = 16'h0094; #100;
A = 16'h0054; B = 16'h0095; #100;
A = 16'h0054; B = 16'h0096; #100;
A = 16'h0054; B = 16'h0097; #100;
A = 16'h0054; B = 16'h0098; #100;
A = 16'h0054; B = 16'h0099; #100;
A = 16'h0054; B = 16'h009A; #100;
A = 16'h0054; B = 16'h009B; #100;
A = 16'h0054; B = 16'h009C; #100;
A = 16'h0054; B = 16'h009D; #100;
A = 16'h0054; B = 16'h009E; #100;
A = 16'h0054; B = 16'h009F; #100;
A = 16'h0054; B = 16'h00A0; #100;
A = 16'h0054; B = 16'h00A1; #100;
A = 16'h0054; B = 16'h00A2; #100;
A = 16'h0054; B = 16'h00A3; #100;
A = 16'h0054; B = 16'h00A4; #100;
A = 16'h0054; B = 16'h00A5; #100;
A = 16'h0054; B = 16'h00A6; #100;
A = 16'h0054; B = 16'h00A7; #100;
A = 16'h0054; B = 16'h00A8; #100;
A = 16'h0054; B = 16'h00A9; #100;
A = 16'h0054; B = 16'h00AA; #100;
A = 16'h0054; B = 16'h00AB; #100;
A = 16'h0054; B = 16'h00AC; #100;
A = 16'h0054; B = 16'h00AD; #100;
A = 16'h0054; B = 16'h00AE; #100;
A = 16'h0054; B = 16'h00AF; #100;
A = 16'h0054; B = 16'h00B0; #100;
A = 16'h0054; B = 16'h00B1; #100;
A = 16'h0054; B = 16'h00B2; #100;
A = 16'h0054; B = 16'h00B3; #100;
A = 16'h0054; B = 16'h00B4; #100;
A = 16'h0054; B = 16'h00B5; #100;
A = 16'h0054; B = 16'h00B6; #100;
A = 16'h0054; B = 16'h00B7; #100;
A = 16'h0054; B = 16'h00B8; #100;
A = 16'h0054; B = 16'h00B9; #100;
A = 16'h0054; B = 16'h00BA; #100;
A = 16'h0054; B = 16'h00BB; #100;
A = 16'h0054; B = 16'h00BC; #100;
A = 16'h0054; B = 16'h00BD; #100;
A = 16'h0054; B = 16'h00BE; #100;
A = 16'h0054; B = 16'h00BF; #100;
A = 16'h0054; B = 16'h00C0; #100;
A = 16'h0054; B = 16'h00C1; #100;
A = 16'h0054; B = 16'h00C2; #100;
A = 16'h0054; B = 16'h00C3; #100;
A = 16'h0054; B = 16'h00C4; #100;
A = 16'h0054; B = 16'h00C5; #100;
A = 16'h0054; B = 16'h00C6; #100;
A = 16'h0054; B = 16'h00C7; #100;
A = 16'h0054; B = 16'h00C8; #100;
A = 16'h0054; B = 16'h00C9; #100;
A = 16'h0054; B = 16'h00CA; #100;
A = 16'h0054; B = 16'h00CB; #100;
A = 16'h0054; B = 16'h00CC; #100;
A = 16'h0054; B = 16'h00CD; #100;
A = 16'h0054; B = 16'h00CE; #100;
A = 16'h0054; B = 16'h00CF; #100;
A = 16'h0054; B = 16'h00D0; #100;
A = 16'h0054; B = 16'h00D1; #100;
A = 16'h0054; B = 16'h00D2; #100;
A = 16'h0054; B = 16'h00D3; #100;
A = 16'h0054; B = 16'h00D4; #100;
A = 16'h0054; B = 16'h00D5; #100;
A = 16'h0054; B = 16'h00D6; #100;
A = 16'h0054; B = 16'h00D7; #100;
A = 16'h0054; B = 16'h00D8; #100;
A = 16'h0054; B = 16'h00D9; #100;
A = 16'h0054; B = 16'h00DA; #100;
A = 16'h0054; B = 16'h00DB; #100;
A = 16'h0054; B = 16'h00DC; #100;
A = 16'h0054; B = 16'h00DD; #100;
A = 16'h0054; B = 16'h00DE; #100;
A = 16'h0054; B = 16'h00DF; #100;
A = 16'h0054; B = 16'h00E0; #100;
A = 16'h0054; B = 16'h00E1; #100;
A = 16'h0054; B = 16'h00E2; #100;
A = 16'h0054; B = 16'h00E3; #100;
A = 16'h0054; B = 16'h00E4; #100;
A = 16'h0054; B = 16'h00E5; #100;
A = 16'h0054; B = 16'h00E6; #100;
A = 16'h0054; B = 16'h00E7; #100;
A = 16'h0054; B = 16'h00E8; #100;
A = 16'h0054; B = 16'h00E9; #100;
A = 16'h0054; B = 16'h00EA; #100;
A = 16'h0054; B = 16'h00EB; #100;
A = 16'h0054; B = 16'h00EC; #100;
A = 16'h0054; B = 16'h00ED; #100;
A = 16'h0054; B = 16'h00EE; #100;
A = 16'h0054; B = 16'h00EF; #100;
A = 16'h0054; B = 16'h00F0; #100;
A = 16'h0054; B = 16'h00F1; #100;
A = 16'h0054; B = 16'h00F2; #100;
A = 16'h0054; B = 16'h00F3; #100;
A = 16'h0054; B = 16'h00F4; #100;
A = 16'h0054; B = 16'h00F5; #100;
A = 16'h0054; B = 16'h00F6; #100;
A = 16'h0054; B = 16'h00F7; #100;
A = 16'h0054; B = 16'h00F8; #100;
A = 16'h0054; B = 16'h00F9; #100;
A = 16'h0054; B = 16'h00FA; #100;
A = 16'h0054; B = 16'h00FB; #100;
A = 16'h0054; B = 16'h00FC; #100;
A = 16'h0054; B = 16'h00FD; #100;
A = 16'h0054; B = 16'h00FE; #100;
A = 16'h0054; B = 16'h00FF; #100;
A = 16'h0055; B = 16'h000; #100;
A = 16'h0055; B = 16'h001; #100;
A = 16'h0055; B = 16'h002; #100;
A = 16'h0055; B = 16'h003; #100;
A = 16'h0055; B = 16'h004; #100;
A = 16'h0055; B = 16'h005; #100;
A = 16'h0055; B = 16'h006; #100;
A = 16'h0055; B = 16'h007; #100;
A = 16'h0055; B = 16'h008; #100;
A = 16'h0055; B = 16'h009; #100;
A = 16'h0055; B = 16'h00A; #100;
A = 16'h0055; B = 16'h00B; #100;
A = 16'h0055; B = 16'h00C; #100;
A = 16'h0055; B = 16'h00D; #100;
A = 16'h0055; B = 16'h00E; #100;
A = 16'h0055; B = 16'h00F; #100;
A = 16'h0055; B = 16'h0010; #100;
A = 16'h0055; B = 16'h0011; #100;
A = 16'h0055; B = 16'h0012; #100;
A = 16'h0055; B = 16'h0013; #100;
A = 16'h0055; B = 16'h0014; #100;
A = 16'h0055; B = 16'h0015; #100;
A = 16'h0055; B = 16'h0016; #100;
A = 16'h0055; B = 16'h0017; #100;
A = 16'h0055; B = 16'h0018; #100;
A = 16'h0055; B = 16'h0019; #100;
A = 16'h0055; B = 16'h001A; #100;
A = 16'h0055; B = 16'h001B; #100;
A = 16'h0055; B = 16'h001C; #100;
A = 16'h0055; B = 16'h001D; #100;
A = 16'h0055; B = 16'h001E; #100;
A = 16'h0055; B = 16'h001F; #100;
A = 16'h0055; B = 16'h0020; #100;
A = 16'h0055; B = 16'h0021; #100;
A = 16'h0055; B = 16'h0022; #100;
A = 16'h0055; B = 16'h0023; #100;
A = 16'h0055; B = 16'h0024; #100;
A = 16'h0055; B = 16'h0025; #100;
A = 16'h0055; B = 16'h0026; #100;
A = 16'h0055; B = 16'h0027; #100;
A = 16'h0055; B = 16'h0028; #100;
A = 16'h0055; B = 16'h0029; #100;
A = 16'h0055; B = 16'h002A; #100;
A = 16'h0055; B = 16'h002B; #100;
A = 16'h0055; B = 16'h002C; #100;
A = 16'h0055; B = 16'h002D; #100;
A = 16'h0055; B = 16'h002E; #100;
A = 16'h0055; B = 16'h002F; #100;
A = 16'h0055; B = 16'h0030; #100;
A = 16'h0055; B = 16'h0031; #100;
A = 16'h0055; B = 16'h0032; #100;
A = 16'h0055; B = 16'h0033; #100;
A = 16'h0055; B = 16'h0034; #100;
A = 16'h0055; B = 16'h0035; #100;
A = 16'h0055; B = 16'h0036; #100;
A = 16'h0055; B = 16'h0037; #100;
A = 16'h0055; B = 16'h0038; #100;
A = 16'h0055; B = 16'h0039; #100;
A = 16'h0055; B = 16'h003A; #100;
A = 16'h0055; B = 16'h003B; #100;
A = 16'h0055; B = 16'h003C; #100;
A = 16'h0055; B = 16'h003D; #100;
A = 16'h0055; B = 16'h003E; #100;
A = 16'h0055; B = 16'h003F; #100;
A = 16'h0055; B = 16'h0040; #100;
A = 16'h0055; B = 16'h0041; #100;
A = 16'h0055; B = 16'h0042; #100;
A = 16'h0055; B = 16'h0043; #100;
A = 16'h0055; B = 16'h0044; #100;
A = 16'h0055; B = 16'h0045; #100;
A = 16'h0055; B = 16'h0046; #100;
A = 16'h0055; B = 16'h0047; #100;
A = 16'h0055; B = 16'h0048; #100;
A = 16'h0055; B = 16'h0049; #100;
A = 16'h0055; B = 16'h004A; #100;
A = 16'h0055; B = 16'h004B; #100;
A = 16'h0055; B = 16'h004C; #100;
A = 16'h0055; B = 16'h004D; #100;
A = 16'h0055; B = 16'h004E; #100;
A = 16'h0055; B = 16'h004F; #100;
A = 16'h0055; B = 16'h0050; #100;
A = 16'h0055; B = 16'h0051; #100;
A = 16'h0055; B = 16'h0052; #100;
A = 16'h0055; B = 16'h0053; #100;
A = 16'h0055; B = 16'h0054; #100;
A = 16'h0055; B = 16'h0055; #100;
A = 16'h0055; B = 16'h0056; #100;
A = 16'h0055; B = 16'h0057; #100;
A = 16'h0055; B = 16'h0058; #100;
A = 16'h0055; B = 16'h0059; #100;
A = 16'h0055; B = 16'h005A; #100;
A = 16'h0055; B = 16'h005B; #100;
A = 16'h0055; B = 16'h005C; #100;
A = 16'h0055; B = 16'h005D; #100;
A = 16'h0055; B = 16'h005E; #100;
A = 16'h0055; B = 16'h005F; #100;
A = 16'h0055; B = 16'h0060; #100;
A = 16'h0055; B = 16'h0061; #100;
A = 16'h0055; B = 16'h0062; #100;
A = 16'h0055; B = 16'h0063; #100;
A = 16'h0055; B = 16'h0064; #100;
A = 16'h0055; B = 16'h0065; #100;
A = 16'h0055; B = 16'h0066; #100;
A = 16'h0055; B = 16'h0067; #100;
A = 16'h0055; B = 16'h0068; #100;
A = 16'h0055; B = 16'h0069; #100;
A = 16'h0055; B = 16'h006A; #100;
A = 16'h0055; B = 16'h006B; #100;
A = 16'h0055; B = 16'h006C; #100;
A = 16'h0055; B = 16'h006D; #100;
A = 16'h0055; B = 16'h006E; #100;
A = 16'h0055; B = 16'h006F; #100;
A = 16'h0055; B = 16'h0070; #100;
A = 16'h0055; B = 16'h0071; #100;
A = 16'h0055; B = 16'h0072; #100;
A = 16'h0055; B = 16'h0073; #100;
A = 16'h0055; B = 16'h0074; #100;
A = 16'h0055; B = 16'h0075; #100;
A = 16'h0055; B = 16'h0076; #100;
A = 16'h0055; B = 16'h0077; #100;
A = 16'h0055; B = 16'h0078; #100;
A = 16'h0055; B = 16'h0079; #100;
A = 16'h0055; B = 16'h007A; #100;
A = 16'h0055; B = 16'h007B; #100;
A = 16'h0055; B = 16'h007C; #100;
A = 16'h0055; B = 16'h007D; #100;
A = 16'h0055; B = 16'h007E; #100;
A = 16'h0055; B = 16'h007F; #100;
A = 16'h0055; B = 16'h0080; #100;
A = 16'h0055; B = 16'h0081; #100;
A = 16'h0055; B = 16'h0082; #100;
A = 16'h0055; B = 16'h0083; #100;
A = 16'h0055; B = 16'h0084; #100;
A = 16'h0055; B = 16'h0085; #100;
A = 16'h0055; B = 16'h0086; #100;
A = 16'h0055; B = 16'h0087; #100;
A = 16'h0055; B = 16'h0088; #100;
A = 16'h0055; B = 16'h0089; #100;
A = 16'h0055; B = 16'h008A; #100;
A = 16'h0055; B = 16'h008B; #100;
A = 16'h0055; B = 16'h008C; #100;
A = 16'h0055; B = 16'h008D; #100;
A = 16'h0055; B = 16'h008E; #100;
A = 16'h0055; B = 16'h008F; #100;
A = 16'h0055; B = 16'h0090; #100;
A = 16'h0055; B = 16'h0091; #100;
A = 16'h0055; B = 16'h0092; #100;
A = 16'h0055; B = 16'h0093; #100;
A = 16'h0055; B = 16'h0094; #100;
A = 16'h0055; B = 16'h0095; #100;
A = 16'h0055; B = 16'h0096; #100;
A = 16'h0055; B = 16'h0097; #100;
A = 16'h0055; B = 16'h0098; #100;
A = 16'h0055; B = 16'h0099; #100;
A = 16'h0055; B = 16'h009A; #100;
A = 16'h0055; B = 16'h009B; #100;
A = 16'h0055; B = 16'h009C; #100;
A = 16'h0055; B = 16'h009D; #100;
A = 16'h0055; B = 16'h009E; #100;
A = 16'h0055; B = 16'h009F; #100;
A = 16'h0055; B = 16'h00A0; #100;
A = 16'h0055; B = 16'h00A1; #100;
A = 16'h0055; B = 16'h00A2; #100;
A = 16'h0055; B = 16'h00A3; #100;
A = 16'h0055; B = 16'h00A4; #100;
A = 16'h0055; B = 16'h00A5; #100;
A = 16'h0055; B = 16'h00A6; #100;
A = 16'h0055; B = 16'h00A7; #100;
A = 16'h0055; B = 16'h00A8; #100;
A = 16'h0055; B = 16'h00A9; #100;
A = 16'h0055; B = 16'h00AA; #100;
A = 16'h0055; B = 16'h00AB; #100;
A = 16'h0055; B = 16'h00AC; #100;
A = 16'h0055; B = 16'h00AD; #100;
A = 16'h0055; B = 16'h00AE; #100;
A = 16'h0055; B = 16'h00AF; #100;
A = 16'h0055; B = 16'h00B0; #100;
A = 16'h0055; B = 16'h00B1; #100;
A = 16'h0055; B = 16'h00B2; #100;
A = 16'h0055; B = 16'h00B3; #100;
A = 16'h0055; B = 16'h00B4; #100;
A = 16'h0055; B = 16'h00B5; #100;
A = 16'h0055; B = 16'h00B6; #100;
A = 16'h0055; B = 16'h00B7; #100;
A = 16'h0055; B = 16'h00B8; #100;
A = 16'h0055; B = 16'h00B9; #100;
A = 16'h0055; B = 16'h00BA; #100;
A = 16'h0055; B = 16'h00BB; #100;
A = 16'h0055; B = 16'h00BC; #100;
A = 16'h0055; B = 16'h00BD; #100;
A = 16'h0055; B = 16'h00BE; #100;
A = 16'h0055; B = 16'h00BF; #100;
A = 16'h0055; B = 16'h00C0; #100;
A = 16'h0055; B = 16'h00C1; #100;
A = 16'h0055; B = 16'h00C2; #100;
A = 16'h0055; B = 16'h00C3; #100;
A = 16'h0055; B = 16'h00C4; #100;
A = 16'h0055; B = 16'h00C5; #100;
A = 16'h0055; B = 16'h00C6; #100;
A = 16'h0055; B = 16'h00C7; #100;
A = 16'h0055; B = 16'h00C8; #100;
A = 16'h0055; B = 16'h00C9; #100;
A = 16'h0055; B = 16'h00CA; #100;
A = 16'h0055; B = 16'h00CB; #100;
A = 16'h0055; B = 16'h00CC; #100;
A = 16'h0055; B = 16'h00CD; #100;
A = 16'h0055; B = 16'h00CE; #100;
A = 16'h0055; B = 16'h00CF; #100;
A = 16'h0055; B = 16'h00D0; #100;
A = 16'h0055; B = 16'h00D1; #100;
A = 16'h0055; B = 16'h00D2; #100;
A = 16'h0055; B = 16'h00D3; #100;
A = 16'h0055; B = 16'h00D4; #100;
A = 16'h0055; B = 16'h00D5; #100;
A = 16'h0055; B = 16'h00D6; #100;
A = 16'h0055; B = 16'h00D7; #100;
A = 16'h0055; B = 16'h00D8; #100;
A = 16'h0055; B = 16'h00D9; #100;
A = 16'h0055; B = 16'h00DA; #100;
A = 16'h0055; B = 16'h00DB; #100;
A = 16'h0055; B = 16'h00DC; #100;
A = 16'h0055; B = 16'h00DD; #100;
A = 16'h0055; B = 16'h00DE; #100;
A = 16'h0055; B = 16'h00DF; #100;
A = 16'h0055; B = 16'h00E0; #100;
A = 16'h0055; B = 16'h00E1; #100;
A = 16'h0055; B = 16'h00E2; #100;
A = 16'h0055; B = 16'h00E3; #100;
A = 16'h0055; B = 16'h00E4; #100;
A = 16'h0055; B = 16'h00E5; #100;
A = 16'h0055; B = 16'h00E6; #100;
A = 16'h0055; B = 16'h00E7; #100;
A = 16'h0055; B = 16'h00E8; #100;
A = 16'h0055; B = 16'h00E9; #100;
A = 16'h0055; B = 16'h00EA; #100;
A = 16'h0055; B = 16'h00EB; #100;
A = 16'h0055; B = 16'h00EC; #100;
A = 16'h0055; B = 16'h00ED; #100;
A = 16'h0055; B = 16'h00EE; #100;
A = 16'h0055; B = 16'h00EF; #100;
A = 16'h0055; B = 16'h00F0; #100;
A = 16'h0055; B = 16'h00F1; #100;
A = 16'h0055; B = 16'h00F2; #100;
A = 16'h0055; B = 16'h00F3; #100;
A = 16'h0055; B = 16'h00F4; #100;
A = 16'h0055; B = 16'h00F5; #100;
A = 16'h0055; B = 16'h00F6; #100;
A = 16'h0055; B = 16'h00F7; #100;
A = 16'h0055; B = 16'h00F8; #100;
A = 16'h0055; B = 16'h00F9; #100;
A = 16'h0055; B = 16'h00FA; #100;
A = 16'h0055; B = 16'h00FB; #100;
A = 16'h0055; B = 16'h00FC; #100;
A = 16'h0055; B = 16'h00FD; #100;
A = 16'h0055; B = 16'h00FE; #100;
A = 16'h0055; B = 16'h00FF; #100;
A = 16'h0056; B = 16'h000; #100;
A = 16'h0056; B = 16'h001; #100;
A = 16'h0056; B = 16'h002; #100;
A = 16'h0056; B = 16'h003; #100;
A = 16'h0056; B = 16'h004; #100;
A = 16'h0056; B = 16'h005; #100;
A = 16'h0056; B = 16'h006; #100;
A = 16'h0056; B = 16'h007; #100;
A = 16'h0056; B = 16'h008; #100;
A = 16'h0056; B = 16'h009; #100;
A = 16'h0056; B = 16'h00A; #100;
A = 16'h0056; B = 16'h00B; #100;
A = 16'h0056; B = 16'h00C; #100;
A = 16'h0056; B = 16'h00D; #100;
A = 16'h0056; B = 16'h00E; #100;
A = 16'h0056; B = 16'h00F; #100;
A = 16'h0056; B = 16'h0010; #100;
A = 16'h0056; B = 16'h0011; #100;
A = 16'h0056; B = 16'h0012; #100;
A = 16'h0056; B = 16'h0013; #100;
A = 16'h0056; B = 16'h0014; #100;
A = 16'h0056; B = 16'h0015; #100;
A = 16'h0056; B = 16'h0016; #100;
A = 16'h0056; B = 16'h0017; #100;
A = 16'h0056; B = 16'h0018; #100;
A = 16'h0056; B = 16'h0019; #100;
A = 16'h0056; B = 16'h001A; #100;
A = 16'h0056; B = 16'h001B; #100;
A = 16'h0056; B = 16'h001C; #100;
A = 16'h0056; B = 16'h001D; #100;
A = 16'h0056; B = 16'h001E; #100;
A = 16'h0056; B = 16'h001F; #100;
A = 16'h0056; B = 16'h0020; #100;
A = 16'h0056; B = 16'h0021; #100;
A = 16'h0056; B = 16'h0022; #100;
A = 16'h0056; B = 16'h0023; #100;
A = 16'h0056; B = 16'h0024; #100;
A = 16'h0056; B = 16'h0025; #100;
A = 16'h0056; B = 16'h0026; #100;
A = 16'h0056; B = 16'h0027; #100;
A = 16'h0056; B = 16'h0028; #100;
A = 16'h0056; B = 16'h0029; #100;
A = 16'h0056; B = 16'h002A; #100;
A = 16'h0056; B = 16'h002B; #100;
A = 16'h0056; B = 16'h002C; #100;
A = 16'h0056; B = 16'h002D; #100;
A = 16'h0056; B = 16'h002E; #100;
A = 16'h0056; B = 16'h002F; #100;
A = 16'h0056; B = 16'h0030; #100;
A = 16'h0056; B = 16'h0031; #100;
A = 16'h0056; B = 16'h0032; #100;
A = 16'h0056; B = 16'h0033; #100;
A = 16'h0056; B = 16'h0034; #100;
A = 16'h0056; B = 16'h0035; #100;
A = 16'h0056; B = 16'h0036; #100;
A = 16'h0056; B = 16'h0037; #100;
A = 16'h0056; B = 16'h0038; #100;
A = 16'h0056; B = 16'h0039; #100;
A = 16'h0056; B = 16'h003A; #100;
A = 16'h0056; B = 16'h003B; #100;
A = 16'h0056; B = 16'h003C; #100;
A = 16'h0056; B = 16'h003D; #100;
A = 16'h0056; B = 16'h003E; #100;
A = 16'h0056; B = 16'h003F; #100;
A = 16'h0056; B = 16'h0040; #100;
A = 16'h0056; B = 16'h0041; #100;
A = 16'h0056; B = 16'h0042; #100;
A = 16'h0056; B = 16'h0043; #100;
A = 16'h0056; B = 16'h0044; #100;
A = 16'h0056; B = 16'h0045; #100;
A = 16'h0056; B = 16'h0046; #100;
A = 16'h0056; B = 16'h0047; #100;
A = 16'h0056; B = 16'h0048; #100;
A = 16'h0056; B = 16'h0049; #100;
A = 16'h0056; B = 16'h004A; #100;
A = 16'h0056; B = 16'h004B; #100;
A = 16'h0056; B = 16'h004C; #100;
A = 16'h0056; B = 16'h004D; #100;
A = 16'h0056; B = 16'h004E; #100;
A = 16'h0056; B = 16'h004F; #100;
A = 16'h0056; B = 16'h0050; #100;
A = 16'h0056; B = 16'h0051; #100;
A = 16'h0056; B = 16'h0052; #100;
A = 16'h0056; B = 16'h0053; #100;
A = 16'h0056; B = 16'h0054; #100;
A = 16'h0056; B = 16'h0055; #100;
A = 16'h0056; B = 16'h0056; #100;
A = 16'h0056; B = 16'h0057; #100;
A = 16'h0056; B = 16'h0058; #100;
A = 16'h0056; B = 16'h0059; #100;
A = 16'h0056; B = 16'h005A; #100;
A = 16'h0056; B = 16'h005B; #100;
A = 16'h0056; B = 16'h005C; #100;
A = 16'h0056; B = 16'h005D; #100;
A = 16'h0056; B = 16'h005E; #100;
A = 16'h0056; B = 16'h005F; #100;
A = 16'h0056; B = 16'h0060; #100;
A = 16'h0056; B = 16'h0061; #100;
A = 16'h0056; B = 16'h0062; #100;
A = 16'h0056; B = 16'h0063; #100;
A = 16'h0056; B = 16'h0064; #100;
A = 16'h0056; B = 16'h0065; #100;
A = 16'h0056; B = 16'h0066; #100;
A = 16'h0056; B = 16'h0067; #100;
A = 16'h0056; B = 16'h0068; #100;
A = 16'h0056; B = 16'h0069; #100;
A = 16'h0056; B = 16'h006A; #100;
A = 16'h0056; B = 16'h006B; #100;
A = 16'h0056; B = 16'h006C; #100;
A = 16'h0056; B = 16'h006D; #100;
A = 16'h0056; B = 16'h006E; #100;
A = 16'h0056; B = 16'h006F; #100;
A = 16'h0056; B = 16'h0070; #100;
A = 16'h0056; B = 16'h0071; #100;
A = 16'h0056; B = 16'h0072; #100;
A = 16'h0056; B = 16'h0073; #100;
A = 16'h0056; B = 16'h0074; #100;
A = 16'h0056; B = 16'h0075; #100;
A = 16'h0056; B = 16'h0076; #100;
A = 16'h0056; B = 16'h0077; #100;
A = 16'h0056; B = 16'h0078; #100;
A = 16'h0056; B = 16'h0079; #100;
A = 16'h0056; B = 16'h007A; #100;
A = 16'h0056; B = 16'h007B; #100;
A = 16'h0056; B = 16'h007C; #100;
A = 16'h0056; B = 16'h007D; #100;
A = 16'h0056; B = 16'h007E; #100;
A = 16'h0056; B = 16'h007F; #100;
A = 16'h0056; B = 16'h0080; #100;
A = 16'h0056; B = 16'h0081; #100;
A = 16'h0056; B = 16'h0082; #100;
A = 16'h0056; B = 16'h0083; #100;
A = 16'h0056; B = 16'h0084; #100;
A = 16'h0056; B = 16'h0085; #100;
A = 16'h0056; B = 16'h0086; #100;
A = 16'h0056; B = 16'h0087; #100;
A = 16'h0056; B = 16'h0088; #100;
A = 16'h0056; B = 16'h0089; #100;
A = 16'h0056; B = 16'h008A; #100;
A = 16'h0056; B = 16'h008B; #100;
A = 16'h0056; B = 16'h008C; #100;
A = 16'h0056; B = 16'h008D; #100;
A = 16'h0056; B = 16'h008E; #100;
A = 16'h0056; B = 16'h008F; #100;
A = 16'h0056; B = 16'h0090; #100;
A = 16'h0056; B = 16'h0091; #100;
A = 16'h0056; B = 16'h0092; #100;
A = 16'h0056; B = 16'h0093; #100;
A = 16'h0056; B = 16'h0094; #100;
A = 16'h0056; B = 16'h0095; #100;
A = 16'h0056; B = 16'h0096; #100;
A = 16'h0056; B = 16'h0097; #100;
A = 16'h0056; B = 16'h0098; #100;
A = 16'h0056; B = 16'h0099; #100;
A = 16'h0056; B = 16'h009A; #100;
A = 16'h0056; B = 16'h009B; #100;
A = 16'h0056; B = 16'h009C; #100;
A = 16'h0056; B = 16'h009D; #100;
A = 16'h0056; B = 16'h009E; #100;
A = 16'h0056; B = 16'h009F; #100;
A = 16'h0056; B = 16'h00A0; #100;
A = 16'h0056; B = 16'h00A1; #100;
A = 16'h0056; B = 16'h00A2; #100;
A = 16'h0056; B = 16'h00A3; #100;
A = 16'h0056; B = 16'h00A4; #100;
A = 16'h0056; B = 16'h00A5; #100;
A = 16'h0056; B = 16'h00A6; #100;
A = 16'h0056; B = 16'h00A7; #100;
A = 16'h0056; B = 16'h00A8; #100;
A = 16'h0056; B = 16'h00A9; #100;
A = 16'h0056; B = 16'h00AA; #100;
A = 16'h0056; B = 16'h00AB; #100;
A = 16'h0056; B = 16'h00AC; #100;
A = 16'h0056; B = 16'h00AD; #100;
A = 16'h0056; B = 16'h00AE; #100;
A = 16'h0056; B = 16'h00AF; #100;
A = 16'h0056; B = 16'h00B0; #100;
A = 16'h0056; B = 16'h00B1; #100;
A = 16'h0056; B = 16'h00B2; #100;
A = 16'h0056; B = 16'h00B3; #100;
A = 16'h0056; B = 16'h00B4; #100;
A = 16'h0056; B = 16'h00B5; #100;
A = 16'h0056; B = 16'h00B6; #100;
A = 16'h0056; B = 16'h00B7; #100;
A = 16'h0056; B = 16'h00B8; #100;
A = 16'h0056; B = 16'h00B9; #100;
A = 16'h0056; B = 16'h00BA; #100;
A = 16'h0056; B = 16'h00BB; #100;
A = 16'h0056; B = 16'h00BC; #100;
A = 16'h0056; B = 16'h00BD; #100;
A = 16'h0056; B = 16'h00BE; #100;
A = 16'h0056; B = 16'h00BF; #100;
A = 16'h0056; B = 16'h00C0; #100;
A = 16'h0056; B = 16'h00C1; #100;
A = 16'h0056; B = 16'h00C2; #100;
A = 16'h0056; B = 16'h00C3; #100;
A = 16'h0056; B = 16'h00C4; #100;
A = 16'h0056; B = 16'h00C5; #100;
A = 16'h0056; B = 16'h00C6; #100;
A = 16'h0056; B = 16'h00C7; #100;
A = 16'h0056; B = 16'h00C8; #100;
A = 16'h0056; B = 16'h00C9; #100;
A = 16'h0056; B = 16'h00CA; #100;
A = 16'h0056; B = 16'h00CB; #100;
A = 16'h0056; B = 16'h00CC; #100;
A = 16'h0056; B = 16'h00CD; #100;
A = 16'h0056; B = 16'h00CE; #100;
A = 16'h0056; B = 16'h00CF; #100;
A = 16'h0056; B = 16'h00D0; #100;
A = 16'h0056; B = 16'h00D1; #100;
A = 16'h0056; B = 16'h00D2; #100;
A = 16'h0056; B = 16'h00D3; #100;
A = 16'h0056; B = 16'h00D4; #100;
A = 16'h0056; B = 16'h00D5; #100;
A = 16'h0056; B = 16'h00D6; #100;
A = 16'h0056; B = 16'h00D7; #100;
A = 16'h0056; B = 16'h00D8; #100;
A = 16'h0056; B = 16'h00D9; #100;
A = 16'h0056; B = 16'h00DA; #100;
A = 16'h0056; B = 16'h00DB; #100;
A = 16'h0056; B = 16'h00DC; #100;
A = 16'h0056; B = 16'h00DD; #100;
A = 16'h0056; B = 16'h00DE; #100;
A = 16'h0056; B = 16'h00DF; #100;
A = 16'h0056; B = 16'h00E0; #100;
A = 16'h0056; B = 16'h00E1; #100;
A = 16'h0056; B = 16'h00E2; #100;
A = 16'h0056; B = 16'h00E3; #100;
A = 16'h0056; B = 16'h00E4; #100;
A = 16'h0056; B = 16'h00E5; #100;
A = 16'h0056; B = 16'h00E6; #100;
A = 16'h0056; B = 16'h00E7; #100;
A = 16'h0056; B = 16'h00E8; #100;
A = 16'h0056; B = 16'h00E9; #100;
A = 16'h0056; B = 16'h00EA; #100;
A = 16'h0056; B = 16'h00EB; #100;
A = 16'h0056; B = 16'h00EC; #100;
A = 16'h0056; B = 16'h00ED; #100;
A = 16'h0056; B = 16'h00EE; #100;
A = 16'h0056; B = 16'h00EF; #100;
A = 16'h0056; B = 16'h00F0; #100;
A = 16'h0056; B = 16'h00F1; #100;
A = 16'h0056; B = 16'h00F2; #100;
A = 16'h0056; B = 16'h00F3; #100;
A = 16'h0056; B = 16'h00F4; #100;
A = 16'h0056; B = 16'h00F5; #100;
A = 16'h0056; B = 16'h00F6; #100;
A = 16'h0056; B = 16'h00F7; #100;
A = 16'h0056; B = 16'h00F8; #100;
A = 16'h0056; B = 16'h00F9; #100;
A = 16'h0056; B = 16'h00FA; #100;
A = 16'h0056; B = 16'h00FB; #100;
A = 16'h0056; B = 16'h00FC; #100;
A = 16'h0056; B = 16'h00FD; #100;
A = 16'h0056; B = 16'h00FE; #100;
A = 16'h0056; B = 16'h00FF; #100;
A = 16'h0057; B = 16'h000; #100;
A = 16'h0057; B = 16'h001; #100;
A = 16'h0057; B = 16'h002; #100;
A = 16'h0057; B = 16'h003; #100;
A = 16'h0057; B = 16'h004; #100;
A = 16'h0057; B = 16'h005; #100;
A = 16'h0057; B = 16'h006; #100;
A = 16'h0057; B = 16'h007; #100;
A = 16'h0057; B = 16'h008; #100;
A = 16'h0057; B = 16'h009; #100;
A = 16'h0057; B = 16'h00A; #100;
A = 16'h0057; B = 16'h00B; #100;
A = 16'h0057; B = 16'h00C; #100;
A = 16'h0057; B = 16'h00D; #100;
A = 16'h0057; B = 16'h00E; #100;
A = 16'h0057; B = 16'h00F; #100;
A = 16'h0057; B = 16'h0010; #100;
A = 16'h0057; B = 16'h0011; #100;
A = 16'h0057; B = 16'h0012; #100;
A = 16'h0057; B = 16'h0013; #100;
A = 16'h0057; B = 16'h0014; #100;
A = 16'h0057; B = 16'h0015; #100;
A = 16'h0057; B = 16'h0016; #100;
A = 16'h0057; B = 16'h0017; #100;
A = 16'h0057; B = 16'h0018; #100;
A = 16'h0057; B = 16'h0019; #100;
A = 16'h0057; B = 16'h001A; #100;
A = 16'h0057; B = 16'h001B; #100;
A = 16'h0057; B = 16'h001C; #100;
A = 16'h0057; B = 16'h001D; #100;
A = 16'h0057; B = 16'h001E; #100;
A = 16'h0057; B = 16'h001F; #100;
A = 16'h0057; B = 16'h0020; #100;
A = 16'h0057; B = 16'h0021; #100;
A = 16'h0057; B = 16'h0022; #100;
A = 16'h0057; B = 16'h0023; #100;
A = 16'h0057; B = 16'h0024; #100;
A = 16'h0057; B = 16'h0025; #100;
A = 16'h0057; B = 16'h0026; #100;
A = 16'h0057; B = 16'h0027; #100;
A = 16'h0057; B = 16'h0028; #100;
A = 16'h0057; B = 16'h0029; #100;
A = 16'h0057; B = 16'h002A; #100;
A = 16'h0057; B = 16'h002B; #100;
A = 16'h0057; B = 16'h002C; #100;
A = 16'h0057; B = 16'h002D; #100;
A = 16'h0057; B = 16'h002E; #100;
A = 16'h0057; B = 16'h002F; #100;
A = 16'h0057; B = 16'h0030; #100;
A = 16'h0057; B = 16'h0031; #100;
A = 16'h0057; B = 16'h0032; #100;
A = 16'h0057; B = 16'h0033; #100;
A = 16'h0057; B = 16'h0034; #100;
A = 16'h0057; B = 16'h0035; #100;
A = 16'h0057; B = 16'h0036; #100;
A = 16'h0057; B = 16'h0037; #100;
A = 16'h0057; B = 16'h0038; #100;
A = 16'h0057; B = 16'h0039; #100;
A = 16'h0057; B = 16'h003A; #100;
A = 16'h0057; B = 16'h003B; #100;
A = 16'h0057; B = 16'h003C; #100;
A = 16'h0057; B = 16'h003D; #100;
A = 16'h0057; B = 16'h003E; #100;
A = 16'h0057; B = 16'h003F; #100;
A = 16'h0057; B = 16'h0040; #100;
A = 16'h0057; B = 16'h0041; #100;
A = 16'h0057; B = 16'h0042; #100;
A = 16'h0057; B = 16'h0043; #100;
A = 16'h0057; B = 16'h0044; #100;
A = 16'h0057; B = 16'h0045; #100;
A = 16'h0057; B = 16'h0046; #100;
A = 16'h0057; B = 16'h0047; #100;
A = 16'h0057; B = 16'h0048; #100;
A = 16'h0057; B = 16'h0049; #100;
A = 16'h0057; B = 16'h004A; #100;
A = 16'h0057; B = 16'h004B; #100;
A = 16'h0057; B = 16'h004C; #100;
A = 16'h0057; B = 16'h004D; #100;
A = 16'h0057; B = 16'h004E; #100;
A = 16'h0057; B = 16'h004F; #100;
A = 16'h0057; B = 16'h0050; #100;
A = 16'h0057; B = 16'h0051; #100;
A = 16'h0057; B = 16'h0052; #100;
A = 16'h0057; B = 16'h0053; #100;
A = 16'h0057; B = 16'h0054; #100;
A = 16'h0057; B = 16'h0055; #100;
A = 16'h0057; B = 16'h0056; #100;
A = 16'h0057; B = 16'h0057; #100;
A = 16'h0057; B = 16'h0058; #100;
A = 16'h0057; B = 16'h0059; #100;
A = 16'h0057; B = 16'h005A; #100;
A = 16'h0057; B = 16'h005B; #100;
A = 16'h0057; B = 16'h005C; #100;
A = 16'h0057; B = 16'h005D; #100;
A = 16'h0057; B = 16'h005E; #100;
A = 16'h0057; B = 16'h005F; #100;
A = 16'h0057; B = 16'h0060; #100;
A = 16'h0057; B = 16'h0061; #100;
A = 16'h0057; B = 16'h0062; #100;
A = 16'h0057; B = 16'h0063; #100;
A = 16'h0057; B = 16'h0064; #100;
A = 16'h0057; B = 16'h0065; #100;
A = 16'h0057; B = 16'h0066; #100;
A = 16'h0057; B = 16'h0067; #100;
A = 16'h0057; B = 16'h0068; #100;
A = 16'h0057; B = 16'h0069; #100;
A = 16'h0057; B = 16'h006A; #100;
A = 16'h0057; B = 16'h006B; #100;
A = 16'h0057; B = 16'h006C; #100;
A = 16'h0057; B = 16'h006D; #100;
A = 16'h0057; B = 16'h006E; #100;
A = 16'h0057; B = 16'h006F; #100;
A = 16'h0057; B = 16'h0070; #100;
A = 16'h0057; B = 16'h0071; #100;
A = 16'h0057; B = 16'h0072; #100;
A = 16'h0057; B = 16'h0073; #100;
A = 16'h0057; B = 16'h0074; #100;
A = 16'h0057; B = 16'h0075; #100;
A = 16'h0057; B = 16'h0076; #100;
A = 16'h0057; B = 16'h0077; #100;
A = 16'h0057; B = 16'h0078; #100;
A = 16'h0057; B = 16'h0079; #100;
A = 16'h0057; B = 16'h007A; #100;
A = 16'h0057; B = 16'h007B; #100;
A = 16'h0057; B = 16'h007C; #100;
A = 16'h0057; B = 16'h007D; #100;
A = 16'h0057; B = 16'h007E; #100;
A = 16'h0057; B = 16'h007F; #100;
A = 16'h0057; B = 16'h0080; #100;
A = 16'h0057; B = 16'h0081; #100;
A = 16'h0057; B = 16'h0082; #100;
A = 16'h0057; B = 16'h0083; #100;
A = 16'h0057; B = 16'h0084; #100;
A = 16'h0057; B = 16'h0085; #100;
A = 16'h0057; B = 16'h0086; #100;
A = 16'h0057; B = 16'h0087; #100;
A = 16'h0057; B = 16'h0088; #100;
A = 16'h0057; B = 16'h0089; #100;
A = 16'h0057; B = 16'h008A; #100;
A = 16'h0057; B = 16'h008B; #100;
A = 16'h0057; B = 16'h008C; #100;
A = 16'h0057; B = 16'h008D; #100;
A = 16'h0057; B = 16'h008E; #100;
A = 16'h0057; B = 16'h008F; #100;
A = 16'h0057; B = 16'h0090; #100;
A = 16'h0057; B = 16'h0091; #100;
A = 16'h0057; B = 16'h0092; #100;
A = 16'h0057; B = 16'h0093; #100;
A = 16'h0057; B = 16'h0094; #100;
A = 16'h0057; B = 16'h0095; #100;
A = 16'h0057; B = 16'h0096; #100;
A = 16'h0057; B = 16'h0097; #100;
A = 16'h0057; B = 16'h0098; #100;
A = 16'h0057; B = 16'h0099; #100;
A = 16'h0057; B = 16'h009A; #100;
A = 16'h0057; B = 16'h009B; #100;
A = 16'h0057; B = 16'h009C; #100;
A = 16'h0057; B = 16'h009D; #100;
A = 16'h0057; B = 16'h009E; #100;
A = 16'h0057; B = 16'h009F; #100;
A = 16'h0057; B = 16'h00A0; #100;
A = 16'h0057; B = 16'h00A1; #100;
A = 16'h0057; B = 16'h00A2; #100;
A = 16'h0057; B = 16'h00A3; #100;
A = 16'h0057; B = 16'h00A4; #100;
A = 16'h0057; B = 16'h00A5; #100;
A = 16'h0057; B = 16'h00A6; #100;
A = 16'h0057; B = 16'h00A7; #100;
A = 16'h0057; B = 16'h00A8; #100;
A = 16'h0057; B = 16'h00A9; #100;
A = 16'h0057; B = 16'h00AA; #100;
A = 16'h0057; B = 16'h00AB; #100;
A = 16'h0057; B = 16'h00AC; #100;
A = 16'h0057; B = 16'h00AD; #100;
A = 16'h0057; B = 16'h00AE; #100;
A = 16'h0057; B = 16'h00AF; #100;
A = 16'h0057; B = 16'h00B0; #100;
A = 16'h0057; B = 16'h00B1; #100;
A = 16'h0057; B = 16'h00B2; #100;
A = 16'h0057; B = 16'h00B3; #100;
A = 16'h0057; B = 16'h00B4; #100;
A = 16'h0057; B = 16'h00B5; #100;
A = 16'h0057; B = 16'h00B6; #100;
A = 16'h0057; B = 16'h00B7; #100;
A = 16'h0057; B = 16'h00B8; #100;
A = 16'h0057; B = 16'h00B9; #100;
A = 16'h0057; B = 16'h00BA; #100;
A = 16'h0057; B = 16'h00BB; #100;
A = 16'h0057; B = 16'h00BC; #100;
A = 16'h0057; B = 16'h00BD; #100;
A = 16'h0057; B = 16'h00BE; #100;
A = 16'h0057; B = 16'h00BF; #100;
A = 16'h0057; B = 16'h00C0; #100;
A = 16'h0057; B = 16'h00C1; #100;
A = 16'h0057; B = 16'h00C2; #100;
A = 16'h0057; B = 16'h00C3; #100;
A = 16'h0057; B = 16'h00C4; #100;
A = 16'h0057; B = 16'h00C5; #100;
A = 16'h0057; B = 16'h00C6; #100;
A = 16'h0057; B = 16'h00C7; #100;
A = 16'h0057; B = 16'h00C8; #100;
A = 16'h0057; B = 16'h00C9; #100;
A = 16'h0057; B = 16'h00CA; #100;
A = 16'h0057; B = 16'h00CB; #100;
A = 16'h0057; B = 16'h00CC; #100;
A = 16'h0057; B = 16'h00CD; #100;
A = 16'h0057; B = 16'h00CE; #100;
A = 16'h0057; B = 16'h00CF; #100;
A = 16'h0057; B = 16'h00D0; #100;
A = 16'h0057; B = 16'h00D1; #100;
A = 16'h0057; B = 16'h00D2; #100;
A = 16'h0057; B = 16'h00D3; #100;
A = 16'h0057; B = 16'h00D4; #100;
A = 16'h0057; B = 16'h00D5; #100;
A = 16'h0057; B = 16'h00D6; #100;
A = 16'h0057; B = 16'h00D7; #100;
A = 16'h0057; B = 16'h00D8; #100;
A = 16'h0057; B = 16'h00D9; #100;
A = 16'h0057; B = 16'h00DA; #100;
A = 16'h0057; B = 16'h00DB; #100;
A = 16'h0057; B = 16'h00DC; #100;
A = 16'h0057; B = 16'h00DD; #100;
A = 16'h0057; B = 16'h00DE; #100;
A = 16'h0057; B = 16'h00DF; #100;
A = 16'h0057; B = 16'h00E0; #100;
A = 16'h0057; B = 16'h00E1; #100;
A = 16'h0057; B = 16'h00E2; #100;
A = 16'h0057; B = 16'h00E3; #100;
A = 16'h0057; B = 16'h00E4; #100;
A = 16'h0057; B = 16'h00E5; #100;
A = 16'h0057; B = 16'h00E6; #100;
A = 16'h0057; B = 16'h00E7; #100;
A = 16'h0057; B = 16'h00E8; #100;
A = 16'h0057; B = 16'h00E9; #100;
A = 16'h0057; B = 16'h00EA; #100;
A = 16'h0057; B = 16'h00EB; #100;
A = 16'h0057; B = 16'h00EC; #100;
A = 16'h0057; B = 16'h00ED; #100;
A = 16'h0057; B = 16'h00EE; #100;
A = 16'h0057; B = 16'h00EF; #100;
A = 16'h0057; B = 16'h00F0; #100;
A = 16'h0057; B = 16'h00F1; #100;
A = 16'h0057; B = 16'h00F2; #100;
A = 16'h0057; B = 16'h00F3; #100;
A = 16'h0057; B = 16'h00F4; #100;
A = 16'h0057; B = 16'h00F5; #100;
A = 16'h0057; B = 16'h00F6; #100;
A = 16'h0057; B = 16'h00F7; #100;
A = 16'h0057; B = 16'h00F8; #100;
A = 16'h0057; B = 16'h00F9; #100;
A = 16'h0057; B = 16'h00FA; #100;
A = 16'h0057; B = 16'h00FB; #100;
A = 16'h0057; B = 16'h00FC; #100;
A = 16'h0057; B = 16'h00FD; #100;
A = 16'h0057; B = 16'h00FE; #100;
A = 16'h0057; B = 16'h00FF; #100;
A = 16'h0058; B = 16'h000; #100;
A = 16'h0058; B = 16'h001; #100;
A = 16'h0058; B = 16'h002; #100;
A = 16'h0058; B = 16'h003; #100;
A = 16'h0058; B = 16'h004; #100;
A = 16'h0058; B = 16'h005; #100;
A = 16'h0058; B = 16'h006; #100;
A = 16'h0058; B = 16'h007; #100;
A = 16'h0058; B = 16'h008; #100;
A = 16'h0058; B = 16'h009; #100;
A = 16'h0058; B = 16'h00A; #100;
A = 16'h0058; B = 16'h00B; #100;
A = 16'h0058; B = 16'h00C; #100;
A = 16'h0058; B = 16'h00D; #100;
A = 16'h0058; B = 16'h00E; #100;
A = 16'h0058; B = 16'h00F; #100;
A = 16'h0058; B = 16'h0010; #100;
A = 16'h0058; B = 16'h0011; #100;
A = 16'h0058; B = 16'h0012; #100;
A = 16'h0058; B = 16'h0013; #100;
A = 16'h0058; B = 16'h0014; #100;
A = 16'h0058; B = 16'h0015; #100;
A = 16'h0058; B = 16'h0016; #100;
A = 16'h0058; B = 16'h0017; #100;
A = 16'h0058; B = 16'h0018; #100;
A = 16'h0058; B = 16'h0019; #100;
A = 16'h0058; B = 16'h001A; #100;
A = 16'h0058; B = 16'h001B; #100;
A = 16'h0058; B = 16'h001C; #100;
A = 16'h0058; B = 16'h001D; #100;
A = 16'h0058; B = 16'h001E; #100;
A = 16'h0058; B = 16'h001F; #100;
A = 16'h0058; B = 16'h0020; #100;
A = 16'h0058; B = 16'h0021; #100;
A = 16'h0058; B = 16'h0022; #100;
A = 16'h0058; B = 16'h0023; #100;
A = 16'h0058; B = 16'h0024; #100;
A = 16'h0058; B = 16'h0025; #100;
A = 16'h0058; B = 16'h0026; #100;
A = 16'h0058; B = 16'h0027; #100;
A = 16'h0058; B = 16'h0028; #100;
A = 16'h0058; B = 16'h0029; #100;
A = 16'h0058; B = 16'h002A; #100;
A = 16'h0058; B = 16'h002B; #100;
A = 16'h0058; B = 16'h002C; #100;
A = 16'h0058; B = 16'h002D; #100;
A = 16'h0058; B = 16'h002E; #100;
A = 16'h0058; B = 16'h002F; #100;
A = 16'h0058; B = 16'h0030; #100;
A = 16'h0058; B = 16'h0031; #100;
A = 16'h0058; B = 16'h0032; #100;
A = 16'h0058; B = 16'h0033; #100;
A = 16'h0058; B = 16'h0034; #100;
A = 16'h0058; B = 16'h0035; #100;
A = 16'h0058; B = 16'h0036; #100;
A = 16'h0058; B = 16'h0037; #100;
A = 16'h0058; B = 16'h0038; #100;
A = 16'h0058; B = 16'h0039; #100;
A = 16'h0058; B = 16'h003A; #100;
A = 16'h0058; B = 16'h003B; #100;
A = 16'h0058; B = 16'h003C; #100;
A = 16'h0058; B = 16'h003D; #100;
A = 16'h0058; B = 16'h003E; #100;
A = 16'h0058; B = 16'h003F; #100;
A = 16'h0058; B = 16'h0040; #100;
A = 16'h0058; B = 16'h0041; #100;
A = 16'h0058; B = 16'h0042; #100;
A = 16'h0058; B = 16'h0043; #100;
A = 16'h0058; B = 16'h0044; #100;
A = 16'h0058; B = 16'h0045; #100;
A = 16'h0058; B = 16'h0046; #100;
A = 16'h0058; B = 16'h0047; #100;
A = 16'h0058; B = 16'h0048; #100;
A = 16'h0058; B = 16'h0049; #100;
A = 16'h0058; B = 16'h004A; #100;
A = 16'h0058; B = 16'h004B; #100;
A = 16'h0058; B = 16'h004C; #100;
A = 16'h0058; B = 16'h004D; #100;
A = 16'h0058; B = 16'h004E; #100;
A = 16'h0058; B = 16'h004F; #100;
A = 16'h0058; B = 16'h0050; #100;
A = 16'h0058; B = 16'h0051; #100;
A = 16'h0058; B = 16'h0052; #100;
A = 16'h0058; B = 16'h0053; #100;
A = 16'h0058; B = 16'h0054; #100;
A = 16'h0058; B = 16'h0055; #100;
A = 16'h0058; B = 16'h0056; #100;
A = 16'h0058; B = 16'h0057; #100;
A = 16'h0058; B = 16'h0058; #100;
A = 16'h0058; B = 16'h0059; #100;
A = 16'h0058; B = 16'h005A; #100;
A = 16'h0058; B = 16'h005B; #100;
A = 16'h0058; B = 16'h005C; #100;
A = 16'h0058; B = 16'h005D; #100;
A = 16'h0058; B = 16'h005E; #100;
A = 16'h0058; B = 16'h005F; #100;
A = 16'h0058; B = 16'h0060; #100;
A = 16'h0058; B = 16'h0061; #100;
A = 16'h0058; B = 16'h0062; #100;
A = 16'h0058; B = 16'h0063; #100;
A = 16'h0058; B = 16'h0064; #100;
A = 16'h0058; B = 16'h0065; #100;
A = 16'h0058; B = 16'h0066; #100;
A = 16'h0058; B = 16'h0067; #100;
A = 16'h0058; B = 16'h0068; #100;
A = 16'h0058; B = 16'h0069; #100;
A = 16'h0058; B = 16'h006A; #100;
A = 16'h0058; B = 16'h006B; #100;
A = 16'h0058; B = 16'h006C; #100;
A = 16'h0058; B = 16'h006D; #100;
A = 16'h0058; B = 16'h006E; #100;
A = 16'h0058; B = 16'h006F; #100;
A = 16'h0058; B = 16'h0070; #100;
A = 16'h0058; B = 16'h0071; #100;
A = 16'h0058; B = 16'h0072; #100;
A = 16'h0058; B = 16'h0073; #100;
A = 16'h0058; B = 16'h0074; #100;
A = 16'h0058; B = 16'h0075; #100;
A = 16'h0058; B = 16'h0076; #100;
A = 16'h0058; B = 16'h0077; #100;
A = 16'h0058; B = 16'h0078; #100;
A = 16'h0058; B = 16'h0079; #100;
A = 16'h0058; B = 16'h007A; #100;
A = 16'h0058; B = 16'h007B; #100;
A = 16'h0058; B = 16'h007C; #100;
A = 16'h0058; B = 16'h007D; #100;
A = 16'h0058; B = 16'h007E; #100;
A = 16'h0058; B = 16'h007F; #100;
A = 16'h0058; B = 16'h0080; #100;
A = 16'h0058; B = 16'h0081; #100;
A = 16'h0058; B = 16'h0082; #100;
A = 16'h0058; B = 16'h0083; #100;
A = 16'h0058; B = 16'h0084; #100;
A = 16'h0058; B = 16'h0085; #100;
A = 16'h0058; B = 16'h0086; #100;
A = 16'h0058; B = 16'h0087; #100;
A = 16'h0058; B = 16'h0088; #100;
A = 16'h0058; B = 16'h0089; #100;
A = 16'h0058; B = 16'h008A; #100;
A = 16'h0058; B = 16'h008B; #100;
A = 16'h0058; B = 16'h008C; #100;
A = 16'h0058; B = 16'h008D; #100;
A = 16'h0058; B = 16'h008E; #100;
A = 16'h0058; B = 16'h008F; #100;
A = 16'h0058; B = 16'h0090; #100;
A = 16'h0058; B = 16'h0091; #100;
A = 16'h0058; B = 16'h0092; #100;
A = 16'h0058; B = 16'h0093; #100;
A = 16'h0058; B = 16'h0094; #100;
A = 16'h0058; B = 16'h0095; #100;
A = 16'h0058; B = 16'h0096; #100;
A = 16'h0058; B = 16'h0097; #100;
A = 16'h0058; B = 16'h0098; #100;
A = 16'h0058; B = 16'h0099; #100;
A = 16'h0058; B = 16'h009A; #100;
A = 16'h0058; B = 16'h009B; #100;
A = 16'h0058; B = 16'h009C; #100;
A = 16'h0058; B = 16'h009D; #100;
A = 16'h0058; B = 16'h009E; #100;
A = 16'h0058; B = 16'h009F; #100;
A = 16'h0058; B = 16'h00A0; #100;
A = 16'h0058; B = 16'h00A1; #100;
A = 16'h0058; B = 16'h00A2; #100;
A = 16'h0058; B = 16'h00A3; #100;
A = 16'h0058; B = 16'h00A4; #100;
A = 16'h0058; B = 16'h00A5; #100;
A = 16'h0058; B = 16'h00A6; #100;
A = 16'h0058; B = 16'h00A7; #100;
A = 16'h0058; B = 16'h00A8; #100;
A = 16'h0058; B = 16'h00A9; #100;
A = 16'h0058; B = 16'h00AA; #100;
A = 16'h0058; B = 16'h00AB; #100;
A = 16'h0058; B = 16'h00AC; #100;
A = 16'h0058; B = 16'h00AD; #100;
A = 16'h0058; B = 16'h00AE; #100;
A = 16'h0058; B = 16'h00AF; #100;
A = 16'h0058; B = 16'h00B0; #100;
A = 16'h0058; B = 16'h00B1; #100;
A = 16'h0058; B = 16'h00B2; #100;
A = 16'h0058; B = 16'h00B3; #100;
A = 16'h0058; B = 16'h00B4; #100;
A = 16'h0058; B = 16'h00B5; #100;
A = 16'h0058; B = 16'h00B6; #100;
A = 16'h0058; B = 16'h00B7; #100;
A = 16'h0058; B = 16'h00B8; #100;
A = 16'h0058; B = 16'h00B9; #100;
A = 16'h0058; B = 16'h00BA; #100;
A = 16'h0058; B = 16'h00BB; #100;
A = 16'h0058; B = 16'h00BC; #100;
A = 16'h0058; B = 16'h00BD; #100;
A = 16'h0058; B = 16'h00BE; #100;
A = 16'h0058; B = 16'h00BF; #100;
A = 16'h0058; B = 16'h00C0; #100;
A = 16'h0058; B = 16'h00C1; #100;
A = 16'h0058; B = 16'h00C2; #100;
A = 16'h0058; B = 16'h00C3; #100;
A = 16'h0058; B = 16'h00C4; #100;
A = 16'h0058; B = 16'h00C5; #100;
A = 16'h0058; B = 16'h00C6; #100;
A = 16'h0058; B = 16'h00C7; #100;
A = 16'h0058; B = 16'h00C8; #100;
A = 16'h0058; B = 16'h00C9; #100;
A = 16'h0058; B = 16'h00CA; #100;
A = 16'h0058; B = 16'h00CB; #100;
A = 16'h0058; B = 16'h00CC; #100;
A = 16'h0058; B = 16'h00CD; #100;
A = 16'h0058; B = 16'h00CE; #100;
A = 16'h0058; B = 16'h00CF; #100;
A = 16'h0058; B = 16'h00D0; #100;
A = 16'h0058; B = 16'h00D1; #100;
A = 16'h0058; B = 16'h00D2; #100;
A = 16'h0058; B = 16'h00D3; #100;
A = 16'h0058; B = 16'h00D4; #100;
A = 16'h0058; B = 16'h00D5; #100;
A = 16'h0058; B = 16'h00D6; #100;
A = 16'h0058; B = 16'h00D7; #100;
A = 16'h0058; B = 16'h00D8; #100;
A = 16'h0058; B = 16'h00D9; #100;
A = 16'h0058; B = 16'h00DA; #100;
A = 16'h0058; B = 16'h00DB; #100;
A = 16'h0058; B = 16'h00DC; #100;
A = 16'h0058; B = 16'h00DD; #100;
A = 16'h0058; B = 16'h00DE; #100;
A = 16'h0058; B = 16'h00DF; #100;
A = 16'h0058; B = 16'h00E0; #100;
A = 16'h0058; B = 16'h00E1; #100;
A = 16'h0058; B = 16'h00E2; #100;
A = 16'h0058; B = 16'h00E3; #100;
A = 16'h0058; B = 16'h00E4; #100;
A = 16'h0058; B = 16'h00E5; #100;
A = 16'h0058; B = 16'h00E6; #100;
A = 16'h0058; B = 16'h00E7; #100;
A = 16'h0058; B = 16'h00E8; #100;
A = 16'h0058; B = 16'h00E9; #100;
A = 16'h0058; B = 16'h00EA; #100;
A = 16'h0058; B = 16'h00EB; #100;
A = 16'h0058; B = 16'h00EC; #100;
A = 16'h0058; B = 16'h00ED; #100;
A = 16'h0058; B = 16'h00EE; #100;
A = 16'h0058; B = 16'h00EF; #100;
A = 16'h0058; B = 16'h00F0; #100;
A = 16'h0058; B = 16'h00F1; #100;
A = 16'h0058; B = 16'h00F2; #100;
A = 16'h0058; B = 16'h00F3; #100;
A = 16'h0058; B = 16'h00F4; #100;
A = 16'h0058; B = 16'h00F5; #100;
A = 16'h0058; B = 16'h00F6; #100;
A = 16'h0058; B = 16'h00F7; #100;
A = 16'h0058; B = 16'h00F8; #100;
A = 16'h0058; B = 16'h00F9; #100;
A = 16'h0058; B = 16'h00FA; #100;
A = 16'h0058; B = 16'h00FB; #100;
A = 16'h0058; B = 16'h00FC; #100;
A = 16'h0058; B = 16'h00FD; #100;
A = 16'h0058; B = 16'h00FE; #100;
A = 16'h0058; B = 16'h00FF; #100;
A = 16'h0059; B = 16'h000; #100;
A = 16'h0059; B = 16'h001; #100;
A = 16'h0059; B = 16'h002; #100;
A = 16'h0059; B = 16'h003; #100;
A = 16'h0059; B = 16'h004; #100;
A = 16'h0059; B = 16'h005; #100;
A = 16'h0059; B = 16'h006; #100;
A = 16'h0059; B = 16'h007; #100;
A = 16'h0059; B = 16'h008; #100;
A = 16'h0059; B = 16'h009; #100;
A = 16'h0059; B = 16'h00A; #100;
A = 16'h0059; B = 16'h00B; #100;
A = 16'h0059; B = 16'h00C; #100;
A = 16'h0059; B = 16'h00D; #100;
A = 16'h0059; B = 16'h00E; #100;
A = 16'h0059; B = 16'h00F; #100;
A = 16'h0059; B = 16'h0010; #100;
A = 16'h0059; B = 16'h0011; #100;
A = 16'h0059; B = 16'h0012; #100;
A = 16'h0059; B = 16'h0013; #100;
A = 16'h0059; B = 16'h0014; #100;
A = 16'h0059; B = 16'h0015; #100;
A = 16'h0059; B = 16'h0016; #100;
A = 16'h0059; B = 16'h0017; #100;
A = 16'h0059; B = 16'h0018; #100;
A = 16'h0059; B = 16'h0019; #100;
A = 16'h0059; B = 16'h001A; #100;
A = 16'h0059; B = 16'h001B; #100;
A = 16'h0059; B = 16'h001C; #100;
A = 16'h0059; B = 16'h001D; #100;
A = 16'h0059; B = 16'h001E; #100;
A = 16'h0059; B = 16'h001F; #100;
A = 16'h0059; B = 16'h0020; #100;
A = 16'h0059; B = 16'h0021; #100;
A = 16'h0059; B = 16'h0022; #100;
A = 16'h0059; B = 16'h0023; #100;
A = 16'h0059; B = 16'h0024; #100;
A = 16'h0059; B = 16'h0025; #100;
A = 16'h0059; B = 16'h0026; #100;
A = 16'h0059; B = 16'h0027; #100;
A = 16'h0059; B = 16'h0028; #100;
A = 16'h0059; B = 16'h0029; #100;
A = 16'h0059; B = 16'h002A; #100;
A = 16'h0059; B = 16'h002B; #100;
A = 16'h0059; B = 16'h002C; #100;
A = 16'h0059; B = 16'h002D; #100;
A = 16'h0059; B = 16'h002E; #100;
A = 16'h0059; B = 16'h002F; #100;
A = 16'h0059; B = 16'h0030; #100;
A = 16'h0059; B = 16'h0031; #100;
A = 16'h0059; B = 16'h0032; #100;
A = 16'h0059; B = 16'h0033; #100;
A = 16'h0059; B = 16'h0034; #100;
A = 16'h0059; B = 16'h0035; #100;
A = 16'h0059; B = 16'h0036; #100;
A = 16'h0059; B = 16'h0037; #100;
A = 16'h0059; B = 16'h0038; #100;
A = 16'h0059; B = 16'h0039; #100;
A = 16'h0059; B = 16'h003A; #100;
A = 16'h0059; B = 16'h003B; #100;
A = 16'h0059; B = 16'h003C; #100;
A = 16'h0059; B = 16'h003D; #100;
A = 16'h0059; B = 16'h003E; #100;
A = 16'h0059; B = 16'h003F; #100;
A = 16'h0059; B = 16'h0040; #100;
A = 16'h0059; B = 16'h0041; #100;
A = 16'h0059; B = 16'h0042; #100;
A = 16'h0059; B = 16'h0043; #100;
A = 16'h0059; B = 16'h0044; #100;
A = 16'h0059; B = 16'h0045; #100;
A = 16'h0059; B = 16'h0046; #100;
A = 16'h0059; B = 16'h0047; #100;
A = 16'h0059; B = 16'h0048; #100;
A = 16'h0059; B = 16'h0049; #100;
A = 16'h0059; B = 16'h004A; #100;
A = 16'h0059; B = 16'h004B; #100;
A = 16'h0059; B = 16'h004C; #100;
A = 16'h0059; B = 16'h004D; #100;
A = 16'h0059; B = 16'h004E; #100;
A = 16'h0059; B = 16'h004F; #100;
A = 16'h0059; B = 16'h0050; #100;
A = 16'h0059; B = 16'h0051; #100;
A = 16'h0059; B = 16'h0052; #100;
A = 16'h0059; B = 16'h0053; #100;
A = 16'h0059; B = 16'h0054; #100;
A = 16'h0059; B = 16'h0055; #100;
A = 16'h0059; B = 16'h0056; #100;
A = 16'h0059; B = 16'h0057; #100;
A = 16'h0059; B = 16'h0058; #100;
A = 16'h0059; B = 16'h0059; #100;
A = 16'h0059; B = 16'h005A; #100;
A = 16'h0059; B = 16'h005B; #100;
A = 16'h0059; B = 16'h005C; #100;
A = 16'h0059; B = 16'h005D; #100;
A = 16'h0059; B = 16'h005E; #100;
A = 16'h0059; B = 16'h005F; #100;
A = 16'h0059; B = 16'h0060; #100;
A = 16'h0059; B = 16'h0061; #100;
A = 16'h0059; B = 16'h0062; #100;
A = 16'h0059; B = 16'h0063; #100;
A = 16'h0059; B = 16'h0064; #100;
A = 16'h0059; B = 16'h0065; #100;
A = 16'h0059; B = 16'h0066; #100;
A = 16'h0059; B = 16'h0067; #100;
A = 16'h0059; B = 16'h0068; #100;
A = 16'h0059; B = 16'h0069; #100;
A = 16'h0059; B = 16'h006A; #100;
A = 16'h0059; B = 16'h006B; #100;
A = 16'h0059; B = 16'h006C; #100;
A = 16'h0059; B = 16'h006D; #100;
A = 16'h0059; B = 16'h006E; #100;
A = 16'h0059; B = 16'h006F; #100;
A = 16'h0059; B = 16'h0070; #100;
A = 16'h0059; B = 16'h0071; #100;
A = 16'h0059; B = 16'h0072; #100;
A = 16'h0059; B = 16'h0073; #100;
A = 16'h0059; B = 16'h0074; #100;
A = 16'h0059; B = 16'h0075; #100;
A = 16'h0059; B = 16'h0076; #100;
A = 16'h0059; B = 16'h0077; #100;
A = 16'h0059; B = 16'h0078; #100;
A = 16'h0059; B = 16'h0079; #100;
A = 16'h0059; B = 16'h007A; #100;
A = 16'h0059; B = 16'h007B; #100;
A = 16'h0059; B = 16'h007C; #100;
A = 16'h0059; B = 16'h007D; #100;
A = 16'h0059; B = 16'h007E; #100;
A = 16'h0059; B = 16'h007F; #100;
A = 16'h0059; B = 16'h0080; #100;
A = 16'h0059; B = 16'h0081; #100;
A = 16'h0059; B = 16'h0082; #100;
A = 16'h0059; B = 16'h0083; #100;
A = 16'h0059; B = 16'h0084; #100;
A = 16'h0059; B = 16'h0085; #100;
A = 16'h0059; B = 16'h0086; #100;
A = 16'h0059; B = 16'h0087; #100;
A = 16'h0059; B = 16'h0088; #100;
A = 16'h0059; B = 16'h0089; #100;
A = 16'h0059; B = 16'h008A; #100;
A = 16'h0059; B = 16'h008B; #100;
A = 16'h0059; B = 16'h008C; #100;
A = 16'h0059; B = 16'h008D; #100;
A = 16'h0059; B = 16'h008E; #100;
A = 16'h0059; B = 16'h008F; #100;
A = 16'h0059; B = 16'h0090; #100;
A = 16'h0059; B = 16'h0091; #100;
A = 16'h0059; B = 16'h0092; #100;
A = 16'h0059; B = 16'h0093; #100;
A = 16'h0059; B = 16'h0094; #100;
A = 16'h0059; B = 16'h0095; #100;
A = 16'h0059; B = 16'h0096; #100;
A = 16'h0059; B = 16'h0097; #100;
A = 16'h0059; B = 16'h0098; #100;
A = 16'h0059; B = 16'h0099; #100;
A = 16'h0059; B = 16'h009A; #100;
A = 16'h0059; B = 16'h009B; #100;
A = 16'h0059; B = 16'h009C; #100;
A = 16'h0059; B = 16'h009D; #100;
A = 16'h0059; B = 16'h009E; #100;
A = 16'h0059; B = 16'h009F; #100;
A = 16'h0059; B = 16'h00A0; #100;
A = 16'h0059; B = 16'h00A1; #100;
A = 16'h0059; B = 16'h00A2; #100;
A = 16'h0059; B = 16'h00A3; #100;
A = 16'h0059; B = 16'h00A4; #100;
A = 16'h0059; B = 16'h00A5; #100;
A = 16'h0059; B = 16'h00A6; #100;
A = 16'h0059; B = 16'h00A7; #100;
A = 16'h0059; B = 16'h00A8; #100;
A = 16'h0059; B = 16'h00A9; #100;
A = 16'h0059; B = 16'h00AA; #100;
A = 16'h0059; B = 16'h00AB; #100;
A = 16'h0059; B = 16'h00AC; #100;
A = 16'h0059; B = 16'h00AD; #100;
A = 16'h0059; B = 16'h00AE; #100;
A = 16'h0059; B = 16'h00AF; #100;
A = 16'h0059; B = 16'h00B0; #100;
A = 16'h0059; B = 16'h00B1; #100;
A = 16'h0059; B = 16'h00B2; #100;
A = 16'h0059; B = 16'h00B3; #100;
A = 16'h0059; B = 16'h00B4; #100;
A = 16'h0059; B = 16'h00B5; #100;
A = 16'h0059; B = 16'h00B6; #100;
A = 16'h0059; B = 16'h00B7; #100;
A = 16'h0059; B = 16'h00B8; #100;
A = 16'h0059; B = 16'h00B9; #100;
A = 16'h0059; B = 16'h00BA; #100;
A = 16'h0059; B = 16'h00BB; #100;
A = 16'h0059; B = 16'h00BC; #100;
A = 16'h0059; B = 16'h00BD; #100;
A = 16'h0059; B = 16'h00BE; #100;
A = 16'h0059; B = 16'h00BF; #100;
A = 16'h0059; B = 16'h00C0; #100;
A = 16'h0059; B = 16'h00C1; #100;
A = 16'h0059; B = 16'h00C2; #100;
A = 16'h0059; B = 16'h00C3; #100;
A = 16'h0059; B = 16'h00C4; #100;
A = 16'h0059; B = 16'h00C5; #100;
A = 16'h0059; B = 16'h00C6; #100;
A = 16'h0059; B = 16'h00C7; #100;
A = 16'h0059; B = 16'h00C8; #100;
A = 16'h0059; B = 16'h00C9; #100;
A = 16'h0059; B = 16'h00CA; #100;
A = 16'h0059; B = 16'h00CB; #100;
A = 16'h0059; B = 16'h00CC; #100;
A = 16'h0059; B = 16'h00CD; #100;
A = 16'h0059; B = 16'h00CE; #100;
A = 16'h0059; B = 16'h00CF; #100;
A = 16'h0059; B = 16'h00D0; #100;
A = 16'h0059; B = 16'h00D1; #100;
A = 16'h0059; B = 16'h00D2; #100;
A = 16'h0059; B = 16'h00D3; #100;
A = 16'h0059; B = 16'h00D4; #100;
A = 16'h0059; B = 16'h00D5; #100;
A = 16'h0059; B = 16'h00D6; #100;
A = 16'h0059; B = 16'h00D7; #100;
A = 16'h0059; B = 16'h00D8; #100;
A = 16'h0059; B = 16'h00D9; #100;
A = 16'h0059; B = 16'h00DA; #100;
A = 16'h0059; B = 16'h00DB; #100;
A = 16'h0059; B = 16'h00DC; #100;
A = 16'h0059; B = 16'h00DD; #100;
A = 16'h0059; B = 16'h00DE; #100;
A = 16'h0059; B = 16'h00DF; #100;
A = 16'h0059; B = 16'h00E0; #100;
A = 16'h0059; B = 16'h00E1; #100;
A = 16'h0059; B = 16'h00E2; #100;
A = 16'h0059; B = 16'h00E3; #100;
A = 16'h0059; B = 16'h00E4; #100;
A = 16'h0059; B = 16'h00E5; #100;
A = 16'h0059; B = 16'h00E6; #100;
A = 16'h0059; B = 16'h00E7; #100;
A = 16'h0059; B = 16'h00E8; #100;
A = 16'h0059; B = 16'h00E9; #100;
A = 16'h0059; B = 16'h00EA; #100;
A = 16'h0059; B = 16'h00EB; #100;
A = 16'h0059; B = 16'h00EC; #100;
A = 16'h0059; B = 16'h00ED; #100;
A = 16'h0059; B = 16'h00EE; #100;
A = 16'h0059; B = 16'h00EF; #100;
A = 16'h0059; B = 16'h00F0; #100;
A = 16'h0059; B = 16'h00F1; #100;
A = 16'h0059; B = 16'h00F2; #100;
A = 16'h0059; B = 16'h00F3; #100;
A = 16'h0059; B = 16'h00F4; #100;
A = 16'h0059; B = 16'h00F5; #100;
A = 16'h0059; B = 16'h00F6; #100;
A = 16'h0059; B = 16'h00F7; #100;
A = 16'h0059; B = 16'h00F8; #100;
A = 16'h0059; B = 16'h00F9; #100;
A = 16'h0059; B = 16'h00FA; #100;
A = 16'h0059; B = 16'h00FB; #100;
A = 16'h0059; B = 16'h00FC; #100;
A = 16'h0059; B = 16'h00FD; #100;
A = 16'h0059; B = 16'h00FE; #100;
A = 16'h0059; B = 16'h00FF; #100;
A = 16'h005A; B = 16'h000; #100;
A = 16'h005A; B = 16'h001; #100;
A = 16'h005A; B = 16'h002; #100;
A = 16'h005A; B = 16'h003; #100;
A = 16'h005A; B = 16'h004; #100;
A = 16'h005A; B = 16'h005; #100;
A = 16'h005A; B = 16'h006; #100;
A = 16'h005A; B = 16'h007; #100;
A = 16'h005A; B = 16'h008; #100;
A = 16'h005A; B = 16'h009; #100;
A = 16'h005A; B = 16'h00A; #100;
A = 16'h005A; B = 16'h00B; #100;
A = 16'h005A; B = 16'h00C; #100;
A = 16'h005A; B = 16'h00D; #100;
A = 16'h005A; B = 16'h00E; #100;
A = 16'h005A; B = 16'h00F; #100;
A = 16'h005A; B = 16'h0010; #100;
A = 16'h005A; B = 16'h0011; #100;
A = 16'h005A; B = 16'h0012; #100;
A = 16'h005A; B = 16'h0013; #100;
A = 16'h005A; B = 16'h0014; #100;
A = 16'h005A; B = 16'h0015; #100;
A = 16'h005A; B = 16'h0016; #100;
A = 16'h005A; B = 16'h0017; #100;
A = 16'h005A; B = 16'h0018; #100;
A = 16'h005A; B = 16'h0019; #100;
A = 16'h005A; B = 16'h001A; #100;
A = 16'h005A; B = 16'h001B; #100;
A = 16'h005A; B = 16'h001C; #100;
A = 16'h005A; B = 16'h001D; #100;
A = 16'h005A; B = 16'h001E; #100;
A = 16'h005A; B = 16'h001F; #100;
A = 16'h005A; B = 16'h0020; #100;
A = 16'h005A; B = 16'h0021; #100;
A = 16'h005A; B = 16'h0022; #100;
A = 16'h005A; B = 16'h0023; #100;
A = 16'h005A; B = 16'h0024; #100;
A = 16'h005A; B = 16'h0025; #100;
A = 16'h005A; B = 16'h0026; #100;
A = 16'h005A; B = 16'h0027; #100;
A = 16'h005A; B = 16'h0028; #100;
A = 16'h005A; B = 16'h0029; #100;
A = 16'h005A; B = 16'h002A; #100;
A = 16'h005A; B = 16'h002B; #100;
A = 16'h005A; B = 16'h002C; #100;
A = 16'h005A; B = 16'h002D; #100;
A = 16'h005A; B = 16'h002E; #100;
A = 16'h005A; B = 16'h002F; #100;
A = 16'h005A; B = 16'h0030; #100;
A = 16'h005A; B = 16'h0031; #100;
A = 16'h005A; B = 16'h0032; #100;
A = 16'h005A; B = 16'h0033; #100;
A = 16'h005A; B = 16'h0034; #100;
A = 16'h005A; B = 16'h0035; #100;
A = 16'h005A; B = 16'h0036; #100;
A = 16'h005A; B = 16'h0037; #100;
A = 16'h005A; B = 16'h0038; #100;
A = 16'h005A; B = 16'h0039; #100;
A = 16'h005A; B = 16'h003A; #100;
A = 16'h005A; B = 16'h003B; #100;
A = 16'h005A; B = 16'h003C; #100;
A = 16'h005A; B = 16'h003D; #100;
A = 16'h005A; B = 16'h003E; #100;
A = 16'h005A; B = 16'h003F; #100;
A = 16'h005A; B = 16'h0040; #100;
A = 16'h005A; B = 16'h0041; #100;
A = 16'h005A; B = 16'h0042; #100;
A = 16'h005A; B = 16'h0043; #100;
A = 16'h005A; B = 16'h0044; #100;
A = 16'h005A; B = 16'h0045; #100;
A = 16'h005A; B = 16'h0046; #100;
A = 16'h005A; B = 16'h0047; #100;
A = 16'h005A; B = 16'h0048; #100;
A = 16'h005A; B = 16'h0049; #100;
A = 16'h005A; B = 16'h004A; #100;
A = 16'h005A; B = 16'h004B; #100;
A = 16'h005A; B = 16'h004C; #100;
A = 16'h005A; B = 16'h004D; #100;
A = 16'h005A; B = 16'h004E; #100;
A = 16'h005A; B = 16'h004F; #100;
A = 16'h005A; B = 16'h0050; #100;
A = 16'h005A; B = 16'h0051; #100;
A = 16'h005A; B = 16'h0052; #100;
A = 16'h005A; B = 16'h0053; #100;
A = 16'h005A; B = 16'h0054; #100;
A = 16'h005A; B = 16'h0055; #100;
A = 16'h005A; B = 16'h0056; #100;
A = 16'h005A; B = 16'h0057; #100;
A = 16'h005A; B = 16'h0058; #100;
A = 16'h005A; B = 16'h0059; #100;
A = 16'h005A; B = 16'h005A; #100;
A = 16'h005A; B = 16'h005B; #100;
A = 16'h005A; B = 16'h005C; #100;
A = 16'h005A; B = 16'h005D; #100;
A = 16'h005A; B = 16'h005E; #100;
A = 16'h005A; B = 16'h005F; #100;
A = 16'h005A; B = 16'h0060; #100;
A = 16'h005A; B = 16'h0061; #100;
A = 16'h005A; B = 16'h0062; #100;
A = 16'h005A; B = 16'h0063; #100;
A = 16'h005A; B = 16'h0064; #100;
A = 16'h005A; B = 16'h0065; #100;
A = 16'h005A; B = 16'h0066; #100;
A = 16'h005A; B = 16'h0067; #100;
A = 16'h005A; B = 16'h0068; #100;
A = 16'h005A; B = 16'h0069; #100;
A = 16'h005A; B = 16'h006A; #100;
A = 16'h005A; B = 16'h006B; #100;
A = 16'h005A; B = 16'h006C; #100;
A = 16'h005A; B = 16'h006D; #100;
A = 16'h005A; B = 16'h006E; #100;
A = 16'h005A; B = 16'h006F; #100;
A = 16'h005A; B = 16'h0070; #100;
A = 16'h005A; B = 16'h0071; #100;
A = 16'h005A; B = 16'h0072; #100;
A = 16'h005A; B = 16'h0073; #100;
A = 16'h005A; B = 16'h0074; #100;
A = 16'h005A; B = 16'h0075; #100;
A = 16'h005A; B = 16'h0076; #100;
A = 16'h005A; B = 16'h0077; #100;
A = 16'h005A; B = 16'h0078; #100;
A = 16'h005A; B = 16'h0079; #100;
A = 16'h005A; B = 16'h007A; #100;
A = 16'h005A; B = 16'h007B; #100;
A = 16'h005A; B = 16'h007C; #100;
A = 16'h005A; B = 16'h007D; #100;
A = 16'h005A; B = 16'h007E; #100;
A = 16'h005A; B = 16'h007F; #100;
A = 16'h005A; B = 16'h0080; #100;
A = 16'h005A; B = 16'h0081; #100;
A = 16'h005A; B = 16'h0082; #100;
A = 16'h005A; B = 16'h0083; #100;
A = 16'h005A; B = 16'h0084; #100;
A = 16'h005A; B = 16'h0085; #100;
A = 16'h005A; B = 16'h0086; #100;
A = 16'h005A; B = 16'h0087; #100;
A = 16'h005A; B = 16'h0088; #100;
A = 16'h005A; B = 16'h0089; #100;
A = 16'h005A; B = 16'h008A; #100;
A = 16'h005A; B = 16'h008B; #100;
A = 16'h005A; B = 16'h008C; #100;
A = 16'h005A; B = 16'h008D; #100;
A = 16'h005A; B = 16'h008E; #100;
A = 16'h005A; B = 16'h008F; #100;
A = 16'h005A; B = 16'h0090; #100;
A = 16'h005A; B = 16'h0091; #100;
A = 16'h005A; B = 16'h0092; #100;
A = 16'h005A; B = 16'h0093; #100;
A = 16'h005A; B = 16'h0094; #100;
A = 16'h005A; B = 16'h0095; #100;
A = 16'h005A; B = 16'h0096; #100;
A = 16'h005A; B = 16'h0097; #100;
A = 16'h005A; B = 16'h0098; #100;
A = 16'h005A; B = 16'h0099; #100;
A = 16'h005A; B = 16'h009A; #100;
A = 16'h005A; B = 16'h009B; #100;
A = 16'h005A; B = 16'h009C; #100;
A = 16'h005A; B = 16'h009D; #100;
A = 16'h005A; B = 16'h009E; #100;
A = 16'h005A; B = 16'h009F; #100;
A = 16'h005A; B = 16'h00A0; #100;
A = 16'h005A; B = 16'h00A1; #100;
A = 16'h005A; B = 16'h00A2; #100;
A = 16'h005A; B = 16'h00A3; #100;
A = 16'h005A; B = 16'h00A4; #100;
A = 16'h005A; B = 16'h00A5; #100;
A = 16'h005A; B = 16'h00A6; #100;
A = 16'h005A; B = 16'h00A7; #100;
A = 16'h005A; B = 16'h00A8; #100;
A = 16'h005A; B = 16'h00A9; #100;
A = 16'h005A; B = 16'h00AA; #100;
A = 16'h005A; B = 16'h00AB; #100;
A = 16'h005A; B = 16'h00AC; #100;
A = 16'h005A; B = 16'h00AD; #100;
A = 16'h005A; B = 16'h00AE; #100;
A = 16'h005A; B = 16'h00AF; #100;
A = 16'h005A; B = 16'h00B0; #100;
A = 16'h005A; B = 16'h00B1; #100;
A = 16'h005A; B = 16'h00B2; #100;
A = 16'h005A; B = 16'h00B3; #100;
A = 16'h005A; B = 16'h00B4; #100;
A = 16'h005A; B = 16'h00B5; #100;
A = 16'h005A; B = 16'h00B6; #100;
A = 16'h005A; B = 16'h00B7; #100;
A = 16'h005A; B = 16'h00B8; #100;
A = 16'h005A; B = 16'h00B9; #100;
A = 16'h005A; B = 16'h00BA; #100;
A = 16'h005A; B = 16'h00BB; #100;
A = 16'h005A; B = 16'h00BC; #100;
A = 16'h005A; B = 16'h00BD; #100;
A = 16'h005A; B = 16'h00BE; #100;
A = 16'h005A; B = 16'h00BF; #100;
A = 16'h005A; B = 16'h00C0; #100;
A = 16'h005A; B = 16'h00C1; #100;
A = 16'h005A; B = 16'h00C2; #100;
A = 16'h005A; B = 16'h00C3; #100;
A = 16'h005A; B = 16'h00C4; #100;
A = 16'h005A; B = 16'h00C5; #100;
A = 16'h005A; B = 16'h00C6; #100;
A = 16'h005A; B = 16'h00C7; #100;
A = 16'h005A; B = 16'h00C8; #100;
A = 16'h005A; B = 16'h00C9; #100;
A = 16'h005A; B = 16'h00CA; #100;
A = 16'h005A; B = 16'h00CB; #100;
A = 16'h005A; B = 16'h00CC; #100;
A = 16'h005A; B = 16'h00CD; #100;
A = 16'h005A; B = 16'h00CE; #100;
A = 16'h005A; B = 16'h00CF; #100;
A = 16'h005A; B = 16'h00D0; #100;
A = 16'h005A; B = 16'h00D1; #100;
A = 16'h005A; B = 16'h00D2; #100;
A = 16'h005A; B = 16'h00D3; #100;
A = 16'h005A; B = 16'h00D4; #100;
A = 16'h005A; B = 16'h00D5; #100;
A = 16'h005A; B = 16'h00D6; #100;
A = 16'h005A; B = 16'h00D7; #100;
A = 16'h005A; B = 16'h00D8; #100;
A = 16'h005A; B = 16'h00D9; #100;
A = 16'h005A; B = 16'h00DA; #100;
A = 16'h005A; B = 16'h00DB; #100;
A = 16'h005A; B = 16'h00DC; #100;
A = 16'h005A; B = 16'h00DD; #100;
A = 16'h005A; B = 16'h00DE; #100;
A = 16'h005A; B = 16'h00DF; #100;
A = 16'h005A; B = 16'h00E0; #100;
A = 16'h005A; B = 16'h00E1; #100;
A = 16'h005A; B = 16'h00E2; #100;
A = 16'h005A; B = 16'h00E3; #100;
A = 16'h005A; B = 16'h00E4; #100;
A = 16'h005A; B = 16'h00E5; #100;
A = 16'h005A; B = 16'h00E6; #100;
A = 16'h005A; B = 16'h00E7; #100;
A = 16'h005A; B = 16'h00E8; #100;
A = 16'h005A; B = 16'h00E9; #100;
A = 16'h005A; B = 16'h00EA; #100;
A = 16'h005A; B = 16'h00EB; #100;
A = 16'h005A; B = 16'h00EC; #100;
A = 16'h005A; B = 16'h00ED; #100;
A = 16'h005A; B = 16'h00EE; #100;
A = 16'h005A; B = 16'h00EF; #100;
A = 16'h005A; B = 16'h00F0; #100;
A = 16'h005A; B = 16'h00F1; #100;
A = 16'h005A; B = 16'h00F2; #100;
A = 16'h005A; B = 16'h00F3; #100;
A = 16'h005A; B = 16'h00F4; #100;
A = 16'h005A; B = 16'h00F5; #100;
A = 16'h005A; B = 16'h00F6; #100;
A = 16'h005A; B = 16'h00F7; #100;
A = 16'h005A; B = 16'h00F8; #100;
A = 16'h005A; B = 16'h00F9; #100;
A = 16'h005A; B = 16'h00FA; #100;
A = 16'h005A; B = 16'h00FB; #100;
A = 16'h005A; B = 16'h00FC; #100;
A = 16'h005A; B = 16'h00FD; #100;
A = 16'h005A; B = 16'h00FE; #100;
A = 16'h005A; B = 16'h00FF; #100;
A = 16'h005B; B = 16'h000; #100;
A = 16'h005B; B = 16'h001; #100;
A = 16'h005B; B = 16'h002; #100;
A = 16'h005B; B = 16'h003; #100;
A = 16'h005B; B = 16'h004; #100;
A = 16'h005B; B = 16'h005; #100;
A = 16'h005B; B = 16'h006; #100;
A = 16'h005B; B = 16'h007; #100;
A = 16'h005B; B = 16'h008; #100;
A = 16'h005B; B = 16'h009; #100;
A = 16'h005B; B = 16'h00A; #100;
A = 16'h005B; B = 16'h00B; #100;
A = 16'h005B; B = 16'h00C; #100;
A = 16'h005B; B = 16'h00D; #100;
A = 16'h005B; B = 16'h00E; #100;
A = 16'h005B; B = 16'h00F; #100;
A = 16'h005B; B = 16'h0010; #100;
A = 16'h005B; B = 16'h0011; #100;
A = 16'h005B; B = 16'h0012; #100;
A = 16'h005B; B = 16'h0013; #100;
A = 16'h005B; B = 16'h0014; #100;
A = 16'h005B; B = 16'h0015; #100;
A = 16'h005B; B = 16'h0016; #100;
A = 16'h005B; B = 16'h0017; #100;
A = 16'h005B; B = 16'h0018; #100;
A = 16'h005B; B = 16'h0019; #100;
A = 16'h005B; B = 16'h001A; #100;
A = 16'h005B; B = 16'h001B; #100;
A = 16'h005B; B = 16'h001C; #100;
A = 16'h005B; B = 16'h001D; #100;
A = 16'h005B; B = 16'h001E; #100;
A = 16'h005B; B = 16'h001F; #100;
A = 16'h005B; B = 16'h0020; #100;
A = 16'h005B; B = 16'h0021; #100;
A = 16'h005B; B = 16'h0022; #100;
A = 16'h005B; B = 16'h0023; #100;
A = 16'h005B; B = 16'h0024; #100;
A = 16'h005B; B = 16'h0025; #100;
A = 16'h005B; B = 16'h0026; #100;
A = 16'h005B; B = 16'h0027; #100;
A = 16'h005B; B = 16'h0028; #100;
A = 16'h005B; B = 16'h0029; #100;
A = 16'h005B; B = 16'h002A; #100;
A = 16'h005B; B = 16'h002B; #100;
A = 16'h005B; B = 16'h002C; #100;
A = 16'h005B; B = 16'h002D; #100;
A = 16'h005B; B = 16'h002E; #100;
A = 16'h005B; B = 16'h002F; #100;
A = 16'h005B; B = 16'h0030; #100;
A = 16'h005B; B = 16'h0031; #100;
A = 16'h005B; B = 16'h0032; #100;
A = 16'h005B; B = 16'h0033; #100;
A = 16'h005B; B = 16'h0034; #100;
A = 16'h005B; B = 16'h0035; #100;
A = 16'h005B; B = 16'h0036; #100;
A = 16'h005B; B = 16'h0037; #100;
A = 16'h005B; B = 16'h0038; #100;
A = 16'h005B; B = 16'h0039; #100;
A = 16'h005B; B = 16'h003A; #100;
A = 16'h005B; B = 16'h003B; #100;
A = 16'h005B; B = 16'h003C; #100;
A = 16'h005B; B = 16'h003D; #100;
A = 16'h005B; B = 16'h003E; #100;
A = 16'h005B; B = 16'h003F; #100;
A = 16'h005B; B = 16'h0040; #100;
A = 16'h005B; B = 16'h0041; #100;
A = 16'h005B; B = 16'h0042; #100;
A = 16'h005B; B = 16'h0043; #100;
A = 16'h005B; B = 16'h0044; #100;
A = 16'h005B; B = 16'h0045; #100;
A = 16'h005B; B = 16'h0046; #100;
A = 16'h005B; B = 16'h0047; #100;
A = 16'h005B; B = 16'h0048; #100;
A = 16'h005B; B = 16'h0049; #100;
A = 16'h005B; B = 16'h004A; #100;
A = 16'h005B; B = 16'h004B; #100;
A = 16'h005B; B = 16'h004C; #100;
A = 16'h005B; B = 16'h004D; #100;
A = 16'h005B; B = 16'h004E; #100;
A = 16'h005B; B = 16'h004F; #100;
A = 16'h005B; B = 16'h0050; #100;
A = 16'h005B; B = 16'h0051; #100;
A = 16'h005B; B = 16'h0052; #100;
A = 16'h005B; B = 16'h0053; #100;
A = 16'h005B; B = 16'h0054; #100;
A = 16'h005B; B = 16'h0055; #100;
A = 16'h005B; B = 16'h0056; #100;
A = 16'h005B; B = 16'h0057; #100;
A = 16'h005B; B = 16'h0058; #100;
A = 16'h005B; B = 16'h0059; #100;
A = 16'h005B; B = 16'h005A; #100;
A = 16'h005B; B = 16'h005B; #100;
A = 16'h005B; B = 16'h005C; #100;
A = 16'h005B; B = 16'h005D; #100;
A = 16'h005B; B = 16'h005E; #100;
A = 16'h005B; B = 16'h005F; #100;
A = 16'h005B; B = 16'h0060; #100;
A = 16'h005B; B = 16'h0061; #100;
A = 16'h005B; B = 16'h0062; #100;
A = 16'h005B; B = 16'h0063; #100;
A = 16'h005B; B = 16'h0064; #100;
A = 16'h005B; B = 16'h0065; #100;
A = 16'h005B; B = 16'h0066; #100;
A = 16'h005B; B = 16'h0067; #100;
A = 16'h005B; B = 16'h0068; #100;
A = 16'h005B; B = 16'h0069; #100;
A = 16'h005B; B = 16'h006A; #100;
A = 16'h005B; B = 16'h006B; #100;
A = 16'h005B; B = 16'h006C; #100;
A = 16'h005B; B = 16'h006D; #100;
A = 16'h005B; B = 16'h006E; #100;
A = 16'h005B; B = 16'h006F; #100;
A = 16'h005B; B = 16'h0070; #100;
A = 16'h005B; B = 16'h0071; #100;
A = 16'h005B; B = 16'h0072; #100;
A = 16'h005B; B = 16'h0073; #100;
A = 16'h005B; B = 16'h0074; #100;
A = 16'h005B; B = 16'h0075; #100;
A = 16'h005B; B = 16'h0076; #100;
A = 16'h005B; B = 16'h0077; #100;
A = 16'h005B; B = 16'h0078; #100;
A = 16'h005B; B = 16'h0079; #100;
A = 16'h005B; B = 16'h007A; #100;
A = 16'h005B; B = 16'h007B; #100;
A = 16'h005B; B = 16'h007C; #100;
A = 16'h005B; B = 16'h007D; #100;
A = 16'h005B; B = 16'h007E; #100;
A = 16'h005B; B = 16'h007F; #100;
A = 16'h005B; B = 16'h0080; #100;
A = 16'h005B; B = 16'h0081; #100;
A = 16'h005B; B = 16'h0082; #100;
A = 16'h005B; B = 16'h0083; #100;
A = 16'h005B; B = 16'h0084; #100;
A = 16'h005B; B = 16'h0085; #100;
A = 16'h005B; B = 16'h0086; #100;
A = 16'h005B; B = 16'h0087; #100;
A = 16'h005B; B = 16'h0088; #100;
A = 16'h005B; B = 16'h0089; #100;
A = 16'h005B; B = 16'h008A; #100;
A = 16'h005B; B = 16'h008B; #100;
A = 16'h005B; B = 16'h008C; #100;
A = 16'h005B; B = 16'h008D; #100;
A = 16'h005B; B = 16'h008E; #100;
A = 16'h005B; B = 16'h008F; #100;
A = 16'h005B; B = 16'h0090; #100;
A = 16'h005B; B = 16'h0091; #100;
A = 16'h005B; B = 16'h0092; #100;
A = 16'h005B; B = 16'h0093; #100;
A = 16'h005B; B = 16'h0094; #100;
A = 16'h005B; B = 16'h0095; #100;
A = 16'h005B; B = 16'h0096; #100;
A = 16'h005B; B = 16'h0097; #100;
A = 16'h005B; B = 16'h0098; #100;
A = 16'h005B; B = 16'h0099; #100;
A = 16'h005B; B = 16'h009A; #100;
A = 16'h005B; B = 16'h009B; #100;
A = 16'h005B; B = 16'h009C; #100;
A = 16'h005B; B = 16'h009D; #100;
A = 16'h005B; B = 16'h009E; #100;
A = 16'h005B; B = 16'h009F; #100;
A = 16'h005B; B = 16'h00A0; #100;
A = 16'h005B; B = 16'h00A1; #100;
A = 16'h005B; B = 16'h00A2; #100;
A = 16'h005B; B = 16'h00A3; #100;
A = 16'h005B; B = 16'h00A4; #100;
A = 16'h005B; B = 16'h00A5; #100;
A = 16'h005B; B = 16'h00A6; #100;
A = 16'h005B; B = 16'h00A7; #100;
A = 16'h005B; B = 16'h00A8; #100;
A = 16'h005B; B = 16'h00A9; #100;
A = 16'h005B; B = 16'h00AA; #100;
A = 16'h005B; B = 16'h00AB; #100;
A = 16'h005B; B = 16'h00AC; #100;
A = 16'h005B; B = 16'h00AD; #100;
A = 16'h005B; B = 16'h00AE; #100;
A = 16'h005B; B = 16'h00AF; #100;
A = 16'h005B; B = 16'h00B0; #100;
A = 16'h005B; B = 16'h00B1; #100;
A = 16'h005B; B = 16'h00B2; #100;
A = 16'h005B; B = 16'h00B3; #100;
A = 16'h005B; B = 16'h00B4; #100;
A = 16'h005B; B = 16'h00B5; #100;
A = 16'h005B; B = 16'h00B6; #100;
A = 16'h005B; B = 16'h00B7; #100;
A = 16'h005B; B = 16'h00B8; #100;
A = 16'h005B; B = 16'h00B9; #100;
A = 16'h005B; B = 16'h00BA; #100;
A = 16'h005B; B = 16'h00BB; #100;
A = 16'h005B; B = 16'h00BC; #100;
A = 16'h005B; B = 16'h00BD; #100;
A = 16'h005B; B = 16'h00BE; #100;
A = 16'h005B; B = 16'h00BF; #100;
A = 16'h005B; B = 16'h00C0; #100;
A = 16'h005B; B = 16'h00C1; #100;
A = 16'h005B; B = 16'h00C2; #100;
A = 16'h005B; B = 16'h00C3; #100;
A = 16'h005B; B = 16'h00C4; #100;
A = 16'h005B; B = 16'h00C5; #100;
A = 16'h005B; B = 16'h00C6; #100;
A = 16'h005B; B = 16'h00C7; #100;
A = 16'h005B; B = 16'h00C8; #100;
A = 16'h005B; B = 16'h00C9; #100;
A = 16'h005B; B = 16'h00CA; #100;
A = 16'h005B; B = 16'h00CB; #100;
A = 16'h005B; B = 16'h00CC; #100;
A = 16'h005B; B = 16'h00CD; #100;
A = 16'h005B; B = 16'h00CE; #100;
A = 16'h005B; B = 16'h00CF; #100;
A = 16'h005B; B = 16'h00D0; #100;
A = 16'h005B; B = 16'h00D1; #100;
A = 16'h005B; B = 16'h00D2; #100;
A = 16'h005B; B = 16'h00D3; #100;
A = 16'h005B; B = 16'h00D4; #100;
A = 16'h005B; B = 16'h00D5; #100;
A = 16'h005B; B = 16'h00D6; #100;
A = 16'h005B; B = 16'h00D7; #100;
A = 16'h005B; B = 16'h00D8; #100;
A = 16'h005B; B = 16'h00D9; #100;
A = 16'h005B; B = 16'h00DA; #100;
A = 16'h005B; B = 16'h00DB; #100;
A = 16'h005B; B = 16'h00DC; #100;
A = 16'h005B; B = 16'h00DD; #100;
A = 16'h005B; B = 16'h00DE; #100;
A = 16'h005B; B = 16'h00DF; #100;
A = 16'h005B; B = 16'h00E0; #100;
A = 16'h005B; B = 16'h00E1; #100;
A = 16'h005B; B = 16'h00E2; #100;
A = 16'h005B; B = 16'h00E3; #100;
A = 16'h005B; B = 16'h00E4; #100;
A = 16'h005B; B = 16'h00E5; #100;
A = 16'h005B; B = 16'h00E6; #100;
A = 16'h005B; B = 16'h00E7; #100;
A = 16'h005B; B = 16'h00E8; #100;
A = 16'h005B; B = 16'h00E9; #100;
A = 16'h005B; B = 16'h00EA; #100;
A = 16'h005B; B = 16'h00EB; #100;
A = 16'h005B; B = 16'h00EC; #100;
A = 16'h005B; B = 16'h00ED; #100;
A = 16'h005B; B = 16'h00EE; #100;
A = 16'h005B; B = 16'h00EF; #100;
A = 16'h005B; B = 16'h00F0; #100;
A = 16'h005B; B = 16'h00F1; #100;
A = 16'h005B; B = 16'h00F2; #100;
A = 16'h005B; B = 16'h00F3; #100;
A = 16'h005B; B = 16'h00F4; #100;
A = 16'h005B; B = 16'h00F5; #100;
A = 16'h005B; B = 16'h00F6; #100;
A = 16'h005B; B = 16'h00F7; #100;
A = 16'h005B; B = 16'h00F8; #100;
A = 16'h005B; B = 16'h00F9; #100;
A = 16'h005B; B = 16'h00FA; #100;
A = 16'h005B; B = 16'h00FB; #100;
A = 16'h005B; B = 16'h00FC; #100;
A = 16'h005B; B = 16'h00FD; #100;
A = 16'h005B; B = 16'h00FE; #100;
A = 16'h005B; B = 16'h00FF; #100;
A = 16'h005C; B = 16'h000; #100;
A = 16'h005C; B = 16'h001; #100;
A = 16'h005C; B = 16'h002; #100;
A = 16'h005C; B = 16'h003; #100;
A = 16'h005C; B = 16'h004; #100;
A = 16'h005C; B = 16'h005; #100;
A = 16'h005C; B = 16'h006; #100;
A = 16'h005C; B = 16'h007; #100;
A = 16'h005C; B = 16'h008; #100;
A = 16'h005C; B = 16'h009; #100;
A = 16'h005C; B = 16'h00A; #100;
A = 16'h005C; B = 16'h00B; #100;
A = 16'h005C; B = 16'h00C; #100;
A = 16'h005C; B = 16'h00D; #100;
A = 16'h005C; B = 16'h00E; #100;
A = 16'h005C; B = 16'h00F; #100;
A = 16'h005C; B = 16'h0010; #100;
A = 16'h005C; B = 16'h0011; #100;
A = 16'h005C; B = 16'h0012; #100;
A = 16'h005C; B = 16'h0013; #100;
A = 16'h005C; B = 16'h0014; #100;
A = 16'h005C; B = 16'h0015; #100;
A = 16'h005C; B = 16'h0016; #100;
A = 16'h005C; B = 16'h0017; #100;
A = 16'h005C; B = 16'h0018; #100;
A = 16'h005C; B = 16'h0019; #100;
A = 16'h005C; B = 16'h001A; #100;
A = 16'h005C; B = 16'h001B; #100;
A = 16'h005C; B = 16'h001C; #100;
A = 16'h005C; B = 16'h001D; #100;
A = 16'h005C; B = 16'h001E; #100;
A = 16'h005C; B = 16'h001F; #100;
A = 16'h005C; B = 16'h0020; #100;
A = 16'h005C; B = 16'h0021; #100;
A = 16'h005C; B = 16'h0022; #100;
A = 16'h005C; B = 16'h0023; #100;
A = 16'h005C; B = 16'h0024; #100;
A = 16'h005C; B = 16'h0025; #100;
A = 16'h005C; B = 16'h0026; #100;
A = 16'h005C; B = 16'h0027; #100;
A = 16'h005C; B = 16'h0028; #100;
A = 16'h005C; B = 16'h0029; #100;
A = 16'h005C; B = 16'h002A; #100;
A = 16'h005C; B = 16'h002B; #100;
A = 16'h005C; B = 16'h002C; #100;
A = 16'h005C; B = 16'h002D; #100;
A = 16'h005C; B = 16'h002E; #100;
A = 16'h005C; B = 16'h002F; #100;
A = 16'h005C; B = 16'h0030; #100;
A = 16'h005C; B = 16'h0031; #100;
A = 16'h005C; B = 16'h0032; #100;
A = 16'h005C; B = 16'h0033; #100;
A = 16'h005C; B = 16'h0034; #100;
A = 16'h005C; B = 16'h0035; #100;
A = 16'h005C; B = 16'h0036; #100;
A = 16'h005C; B = 16'h0037; #100;
A = 16'h005C; B = 16'h0038; #100;
A = 16'h005C; B = 16'h0039; #100;
A = 16'h005C; B = 16'h003A; #100;
A = 16'h005C; B = 16'h003B; #100;
A = 16'h005C; B = 16'h003C; #100;
A = 16'h005C; B = 16'h003D; #100;
A = 16'h005C; B = 16'h003E; #100;
A = 16'h005C; B = 16'h003F; #100;
A = 16'h005C; B = 16'h0040; #100;
A = 16'h005C; B = 16'h0041; #100;
A = 16'h005C; B = 16'h0042; #100;
A = 16'h005C; B = 16'h0043; #100;
A = 16'h005C; B = 16'h0044; #100;
A = 16'h005C; B = 16'h0045; #100;
A = 16'h005C; B = 16'h0046; #100;
A = 16'h005C; B = 16'h0047; #100;
A = 16'h005C; B = 16'h0048; #100;
A = 16'h005C; B = 16'h0049; #100;
A = 16'h005C; B = 16'h004A; #100;
A = 16'h005C; B = 16'h004B; #100;
A = 16'h005C; B = 16'h004C; #100;
A = 16'h005C; B = 16'h004D; #100;
A = 16'h005C; B = 16'h004E; #100;
A = 16'h005C; B = 16'h004F; #100;
A = 16'h005C; B = 16'h0050; #100;
A = 16'h005C; B = 16'h0051; #100;
A = 16'h005C; B = 16'h0052; #100;
A = 16'h005C; B = 16'h0053; #100;
A = 16'h005C; B = 16'h0054; #100;
A = 16'h005C; B = 16'h0055; #100;
A = 16'h005C; B = 16'h0056; #100;
A = 16'h005C; B = 16'h0057; #100;
A = 16'h005C; B = 16'h0058; #100;
A = 16'h005C; B = 16'h0059; #100;
A = 16'h005C; B = 16'h005A; #100;
A = 16'h005C; B = 16'h005B; #100;
A = 16'h005C; B = 16'h005C; #100;
A = 16'h005C; B = 16'h005D; #100;
A = 16'h005C; B = 16'h005E; #100;
A = 16'h005C; B = 16'h005F; #100;
A = 16'h005C; B = 16'h0060; #100;
A = 16'h005C; B = 16'h0061; #100;
A = 16'h005C; B = 16'h0062; #100;
A = 16'h005C; B = 16'h0063; #100;
A = 16'h005C; B = 16'h0064; #100;
A = 16'h005C; B = 16'h0065; #100;
A = 16'h005C; B = 16'h0066; #100;
A = 16'h005C; B = 16'h0067; #100;
A = 16'h005C; B = 16'h0068; #100;
A = 16'h005C; B = 16'h0069; #100;
A = 16'h005C; B = 16'h006A; #100;
A = 16'h005C; B = 16'h006B; #100;
A = 16'h005C; B = 16'h006C; #100;
A = 16'h005C; B = 16'h006D; #100;
A = 16'h005C; B = 16'h006E; #100;
A = 16'h005C; B = 16'h006F; #100;
A = 16'h005C; B = 16'h0070; #100;
A = 16'h005C; B = 16'h0071; #100;
A = 16'h005C; B = 16'h0072; #100;
A = 16'h005C; B = 16'h0073; #100;
A = 16'h005C; B = 16'h0074; #100;
A = 16'h005C; B = 16'h0075; #100;
A = 16'h005C; B = 16'h0076; #100;
A = 16'h005C; B = 16'h0077; #100;
A = 16'h005C; B = 16'h0078; #100;
A = 16'h005C; B = 16'h0079; #100;
A = 16'h005C; B = 16'h007A; #100;
A = 16'h005C; B = 16'h007B; #100;
A = 16'h005C; B = 16'h007C; #100;
A = 16'h005C; B = 16'h007D; #100;
A = 16'h005C; B = 16'h007E; #100;
A = 16'h005C; B = 16'h007F; #100;
A = 16'h005C; B = 16'h0080; #100;
A = 16'h005C; B = 16'h0081; #100;
A = 16'h005C; B = 16'h0082; #100;
A = 16'h005C; B = 16'h0083; #100;
A = 16'h005C; B = 16'h0084; #100;
A = 16'h005C; B = 16'h0085; #100;
A = 16'h005C; B = 16'h0086; #100;
A = 16'h005C; B = 16'h0087; #100;
A = 16'h005C; B = 16'h0088; #100;
A = 16'h005C; B = 16'h0089; #100;
A = 16'h005C; B = 16'h008A; #100;
A = 16'h005C; B = 16'h008B; #100;
A = 16'h005C; B = 16'h008C; #100;
A = 16'h005C; B = 16'h008D; #100;
A = 16'h005C; B = 16'h008E; #100;
A = 16'h005C; B = 16'h008F; #100;
A = 16'h005C; B = 16'h0090; #100;
A = 16'h005C; B = 16'h0091; #100;
A = 16'h005C; B = 16'h0092; #100;
A = 16'h005C; B = 16'h0093; #100;
A = 16'h005C; B = 16'h0094; #100;
A = 16'h005C; B = 16'h0095; #100;
A = 16'h005C; B = 16'h0096; #100;
A = 16'h005C; B = 16'h0097; #100;
A = 16'h005C; B = 16'h0098; #100;
A = 16'h005C; B = 16'h0099; #100;
A = 16'h005C; B = 16'h009A; #100;
A = 16'h005C; B = 16'h009B; #100;
A = 16'h005C; B = 16'h009C; #100;
A = 16'h005C; B = 16'h009D; #100;
A = 16'h005C; B = 16'h009E; #100;
A = 16'h005C; B = 16'h009F; #100;
A = 16'h005C; B = 16'h00A0; #100;
A = 16'h005C; B = 16'h00A1; #100;
A = 16'h005C; B = 16'h00A2; #100;
A = 16'h005C; B = 16'h00A3; #100;
A = 16'h005C; B = 16'h00A4; #100;
A = 16'h005C; B = 16'h00A5; #100;
A = 16'h005C; B = 16'h00A6; #100;
A = 16'h005C; B = 16'h00A7; #100;
A = 16'h005C; B = 16'h00A8; #100;
A = 16'h005C; B = 16'h00A9; #100;
A = 16'h005C; B = 16'h00AA; #100;
A = 16'h005C; B = 16'h00AB; #100;
A = 16'h005C; B = 16'h00AC; #100;
A = 16'h005C; B = 16'h00AD; #100;
A = 16'h005C; B = 16'h00AE; #100;
A = 16'h005C; B = 16'h00AF; #100;
A = 16'h005C; B = 16'h00B0; #100;
A = 16'h005C; B = 16'h00B1; #100;
A = 16'h005C; B = 16'h00B2; #100;
A = 16'h005C; B = 16'h00B3; #100;
A = 16'h005C; B = 16'h00B4; #100;
A = 16'h005C; B = 16'h00B5; #100;
A = 16'h005C; B = 16'h00B6; #100;
A = 16'h005C; B = 16'h00B7; #100;
A = 16'h005C; B = 16'h00B8; #100;
A = 16'h005C; B = 16'h00B9; #100;
A = 16'h005C; B = 16'h00BA; #100;
A = 16'h005C; B = 16'h00BB; #100;
A = 16'h005C; B = 16'h00BC; #100;
A = 16'h005C; B = 16'h00BD; #100;
A = 16'h005C; B = 16'h00BE; #100;
A = 16'h005C; B = 16'h00BF; #100;
A = 16'h005C; B = 16'h00C0; #100;
A = 16'h005C; B = 16'h00C1; #100;
A = 16'h005C; B = 16'h00C2; #100;
A = 16'h005C; B = 16'h00C3; #100;
A = 16'h005C; B = 16'h00C4; #100;
A = 16'h005C; B = 16'h00C5; #100;
A = 16'h005C; B = 16'h00C6; #100;
A = 16'h005C; B = 16'h00C7; #100;
A = 16'h005C; B = 16'h00C8; #100;
A = 16'h005C; B = 16'h00C9; #100;
A = 16'h005C; B = 16'h00CA; #100;
A = 16'h005C; B = 16'h00CB; #100;
A = 16'h005C; B = 16'h00CC; #100;
A = 16'h005C; B = 16'h00CD; #100;
A = 16'h005C; B = 16'h00CE; #100;
A = 16'h005C; B = 16'h00CF; #100;
A = 16'h005C; B = 16'h00D0; #100;
A = 16'h005C; B = 16'h00D1; #100;
A = 16'h005C; B = 16'h00D2; #100;
A = 16'h005C; B = 16'h00D3; #100;
A = 16'h005C; B = 16'h00D4; #100;
A = 16'h005C; B = 16'h00D5; #100;
A = 16'h005C; B = 16'h00D6; #100;
A = 16'h005C; B = 16'h00D7; #100;
A = 16'h005C; B = 16'h00D8; #100;
A = 16'h005C; B = 16'h00D9; #100;
A = 16'h005C; B = 16'h00DA; #100;
A = 16'h005C; B = 16'h00DB; #100;
A = 16'h005C; B = 16'h00DC; #100;
A = 16'h005C; B = 16'h00DD; #100;
A = 16'h005C; B = 16'h00DE; #100;
A = 16'h005C; B = 16'h00DF; #100;
A = 16'h005C; B = 16'h00E0; #100;
A = 16'h005C; B = 16'h00E1; #100;
A = 16'h005C; B = 16'h00E2; #100;
A = 16'h005C; B = 16'h00E3; #100;
A = 16'h005C; B = 16'h00E4; #100;
A = 16'h005C; B = 16'h00E5; #100;
A = 16'h005C; B = 16'h00E6; #100;
A = 16'h005C; B = 16'h00E7; #100;
A = 16'h005C; B = 16'h00E8; #100;
A = 16'h005C; B = 16'h00E9; #100;
A = 16'h005C; B = 16'h00EA; #100;
A = 16'h005C; B = 16'h00EB; #100;
A = 16'h005C; B = 16'h00EC; #100;
A = 16'h005C; B = 16'h00ED; #100;
A = 16'h005C; B = 16'h00EE; #100;
A = 16'h005C; B = 16'h00EF; #100;
A = 16'h005C; B = 16'h00F0; #100;
A = 16'h005C; B = 16'h00F1; #100;
A = 16'h005C; B = 16'h00F2; #100;
A = 16'h005C; B = 16'h00F3; #100;
A = 16'h005C; B = 16'h00F4; #100;
A = 16'h005C; B = 16'h00F5; #100;
A = 16'h005C; B = 16'h00F6; #100;
A = 16'h005C; B = 16'h00F7; #100;
A = 16'h005C; B = 16'h00F8; #100;
A = 16'h005C; B = 16'h00F9; #100;
A = 16'h005C; B = 16'h00FA; #100;
A = 16'h005C; B = 16'h00FB; #100;
A = 16'h005C; B = 16'h00FC; #100;
A = 16'h005C; B = 16'h00FD; #100;
A = 16'h005C; B = 16'h00FE; #100;
A = 16'h005C; B = 16'h00FF; #100;
A = 16'h005D; B = 16'h000; #100;
A = 16'h005D; B = 16'h001; #100;
A = 16'h005D; B = 16'h002; #100;
A = 16'h005D; B = 16'h003; #100;
A = 16'h005D; B = 16'h004; #100;
A = 16'h005D; B = 16'h005; #100;
A = 16'h005D; B = 16'h006; #100;
A = 16'h005D; B = 16'h007; #100;
A = 16'h005D; B = 16'h008; #100;
A = 16'h005D; B = 16'h009; #100;
A = 16'h005D; B = 16'h00A; #100;
A = 16'h005D; B = 16'h00B; #100;
A = 16'h005D; B = 16'h00C; #100;
A = 16'h005D; B = 16'h00D; #100;
A = 16'h005D; B = 16'h00E; #100;
A = 16'h005D; B = 16'h00F; #100;
A = 16'h005D; B = 16'h0010; #100;
A = 16'h005D; B = 16'h0011; #100;
A = 16'h005D; B = 16'h0012; #100;
A = 16'h005D; B = 16'h0013; #100;
A = 16'h005D; B = 16'h0014; #100;
A = 16'h005D; B = 16'h0015; #100;
A = 16'h005D; B = 16'h0016; #100;
A = 16'h005D; B = 16'h0017; #100;
A = 16'h005D; B = 16'h0018; #100;
A = 16'h005D; B = 16'h0019; #100;
A = 16'h005D; B = 16'h001A; #100;
A = 16'h005D; B = 16'h001B; #100;
A = 16'h005D; B = 16'h001C; #100;
A = 16'h005D; B = 16'h001D; #100;
A = 16'h005D; B = 16'h001E; #100;
A = 16'h005D; B = 16'h001F; #100;
A = 16'h005D; B = 16'h0020; #100;
A = 16'h005D; B = 16'h0021; #100;
A = 16'h005D; B = 16'h0022; #100;
A = 16'h005D; B = 16'h0023; #100;
A = 16'h005D; B = 16'h0024; #100;
A = 16'h005D; B = 16'h0025; #100;
A = 16'h005D; B = 16'h0026; #100;
A = 16'h005D; B = 16'h0027; #100;
A = 16'h005D; B = 16'h0028; #100;
A = 16'h005D; B = 16'h0029; #100;
A = 16'h005D; B = 16'h002A; #100;
A = 16'h005D; B = 16'h002B; #100;
A = 16'h005D; B = 16'h002C; #100;
A = 16'h005D; B = 16'h002D; #100;
A = 16'h005D; B = 16'h002E; #100;
A = 16'h005D; B = 16'h002F; #100;
A = 16'h005D; B = 16'h0030; #100;
A = 16'h005D; B = 16'h0031; #100;
A = 16'h005D; B = 16'h0032; #100;
A = 16'h005D; B = 16'h0033; #100;
A = 16'h005D; B = 16'h0034; #100;
A = 16'h005D; B = 16'h0035; #100;
A = 16'h005D; B = 16'h0036; #100;
A = 16'h005D; B = 16'h0037; #100;
A = 16'h005D; B = 16'h0038; #100;
A = 16'h005D; B = 16'h0039; #100;
A = 16'h005D; B = 16'h003A; #100;
A = 16'h005D; B = 16'h003B; #100;
A = 16'h005D; B = 16'h003C; #100;
A = 16'h005D; B = 16'h003D; #100;
A = 16'h005D; B = 16'h003E; #100;
A = 16'h005D; B = 16'h003F; #100;
A = 16'h005D; B = 16'h0040; #100;
A = 16'h005D; B = 16'h0041; #100;
A = 16'h005D; B = 16'h0042; #100;
A = 16'h005D; B = 16'h0043; #100;
A = 16'h005D; B = 16'h0044; #100;
A = 16'h005D; B = 16'h0045; #100;
A = 16'h005D; B = 16'h0046; #100;
A = 16'h005D; B = 16'h0047; #100;
A = 16'h005D; B = 16'h0048; #100;
A = 16'h005D; B = 16'h0049; #100;
A = 16'h005D; B = 16'h004A; #100;
A = 16'h005D; B = 16'h004B; #100;
A = 16'h005D; B = 16'h004C; #100;
A = 16'h005D; B = 16'h004D; #100;
A = 16'h005D; B = 16'h004E; #100;
A = 16'h005D; B = 16'h004F; #100;
A = 16'h005D; B = 16'h0050; #100;
A = 16'h005D; B = 16'h0051; #100;
A = 16'h005D; B = 16'h0052; #100;
A = 16'h005D; B = 16'h0053; #100;
A = 16'h005D; B = 16'h0054; #100;
A = 16'h005D; B = 16'h0055; #100;
A = 16'h005D; B = 16'h0056; #100;
A = 16'h005D; B = 16'h0057; #100;
A = 16'h005D; B = 16'h0058; #100;
A = 16'h005D; B = 16'h0059; #100;
A = 16'h005D; B = 16'h005A; #100;
A = 16'h005D; B = 16'h005B; #100;
A = 16'h005D; B = 16'h005C; #100;
A = 16'h005D; B = 16'h005D; #100;
A = 16'h005D; B = 16'h005E; #100;
A = 16'h005D; B = 16'h005F; #100;
A = 16'h005D; B = 16'h0060; #100;
A = 16'h005D; B = 16'h0061; #100;
A = 16'h005D; B = 16'h0062; #100;
A = 16'h005D; B = 16'h0063; #100;
A = 16'h005D; B = 16'h0064; #100;
A = 16'h005D; B = 16'h0065; #100;
A = 16'h005D; B = 16'h0066; #100;
A = 16'h005D; B = 16'h0067; #100;
A = 16'h005D; B = 16'h0068; #100;
A = 16'h005D; B = 16'h0069; #100;
A = 16'h005D; B = 16'h006A; #100;
A = 16'h005D; B = 16'h006B; #100;
A = 16'h005D; B = 16'h006C; #100;
A = 16'h005D; B = 16'h006D; #100;
A = 16'h005D; B = 16'h006E; #100;
A = 16'h005D; B = 16'h006F; #100;
A = 16'h005D; B = 16'h0070; #100;
A = 16'h005D; B = 16'h0071; #100;
A = 16'h005D; B = 16'h0072; #100;
A = 16'h005D; B = 16'h0073; #100;
A = 16'h005D; B = 16'h0074; #100;
A = 16'h005D; B = 16'h0075; #100;
A = 16'h005D; B = 16'h0076; #100;
A = 16'h005D; B = 16'h0077; #100;
A = 16'h005D; B = 16'h0078; #100;
A = 16'h005D; B = 16'h0079; #100;
A = 16'h005D; B = 16'h007A; #100;
A = 16'h005D; B = 16'h007B; #100;
A = 16'h005D; B = 16'h007C; #100;
A = 16'h005D; B = 16'h007D; #100;
A = 16'h005D; B = 16'h007E; #100;
A = 16'h005D; B = 16'h007F; #100;
A = 16'h005D; B = 16'h0080; #100;
A = 16'h005D; B = 16'h0081; #100;
A = 16'h005D; B = 16'h0082; #100;
A = 16'h005D; B = 16'h0083; #100;
A = 16'h005D; B = 16'h0084; #100;
A = 16'h005D; B = 16'h0085; #100;
A = 16'h005D; B = 16'h0086; #100;
A = 16'h005D; B = 16'h0087; #100;
A = 16'h005D; B = 16'h0088; #100;
A = 16'h005D; B = 16'h0089; #100;
A = 16'h005D; B = 16'h008A; #100;
A = 16'h005D; B = 16'h008B; #100;
A = 16'h005D; B = 16'h008C; #100;
A = 16'h005D; B = 16'h008D; #100;
A = 16'h005D; B = 16'h008E; #100;
A = 16'h005D; B = 16'h008F; #100;
A = 16'h005D; B = 16'h0090; #100;
A = 16'h005D; B = 16'h0091; #100;
A = 16'h005D; B = 16'h0092; #100;
A = 16'h005D; B = 16'h0093; #100;
A = 16'h005D; B = 16'h0094; #100;
A = 16'h005D; B = 16'h0095; #100;
A = 16'h005D; B = 16'h0096; #100;
A = 16'h005D; B = 16'h0097; #100;
A = 16'h005D; B = 16'h0098; #100;
A = 16'h005D; B = 16'h0099; #100;
A = 16'h005D; B = 16'h009A; #100;
A = 16'h005D; B = 16'h009B; #100;
A = 16'h005D; B = 16'h009C; #100;
A = 16'h005D; B = 16'h009D; #100;
A = 16'h005D; B = 16'h009E; #100;
A = 16'h005D; B = 16'h009F; #100;
A = 16'h005D; B = 16'h00A0; #100;
A = 16'h005D; B = 16'h00A1; #100;
A = 16'h005D; B = 16'h00A2; #100;
A = 16'h005D; B = 16'h00A3; #100;
A = 16'h005D; B = 16'h00A4; #100;
A = 16'h005D; B = 16'h00A5; #100;
A = 16'h005D; B = 16'h00A6; #100;
A = 16'h005D; B = 16'h00A7; #100;
A = 16'h005D; B = 16'h00A8; #100;
A = 16'h005D; B = 16'h00A9; #100;
A = 16'h005D; B = 16'h00AA; #100;
A = 16'h005D; B = 16'h00AB; #100;
A = 16'h005D; B = 16'h00AC; #100;
A = 16'h005D; B = 16'h00AD; #100;
A = 16'h005D; B = 16'h00AE; #100;
A = 16'h005D; B = 16'h00AF; #100;
A = 16'h005D; B = 16'h00B0; #100;
A = 16'h005D; B = 16'h00B1; #100;
A = 16'h005D; B = 16'h00B2; #100;
A = 16'h005D; B = 16'h00B3; #100;
A = 16'h005D; B = 16'h00B4; #100;
A = 16'h005D; B = 16'h00B5; #100;
A = 16'h005D; B = 16'h00B6; #100;
A = 16'h005D; B = 16'h00B7; #100;
A = 16'h005D; B = 16'h00B8; #100;
A = 16'h005D; B = 16'h00B9; #100;
A = 16'h005D; B = 16'h00BA; #100;
A = 16'h005D; B = 16'h00BB; #100;
A = 16'h005D; B = 16'h00BC; #100;
A = 16'h005D; B = 16'h00BD; #100;
A = 16'h005D; B = 16'h00BE; #100;
A = 16'h005D; B = 16'h00BF; #100;
A = 16'h005D; B = 16'h00C0; #100;
A = 16'h005D; B = 16'h00C1; #100;
A = 16'h005D; B = 16'h00C2; #100;
A = 16'h005D; B = 16'h00C3; #100;
A = 16'h005D; B = 16'h00C4; #100;
A = 16'h005D; B = 16'h00C5; #100;
A = 16'h005D; B = 16'h00C6; #100;
A = 16'h005D; B = 16'h00C7; #100;
A = 16'h005D; B = 16'h00C8; #100;
A = 16'h005D; B = 16'h00C9; #100;
A = 16'h005D; B = 16'h00CA; #100;
A = 16'h005D; B = 16'h00CB; #100;
A = 16'h005D; B = 16'h00CC; #100;
A = 16'h005D; B = 16'h00CD; #100;
A = 16'h005D; B = 16'h00CE; #100;
A = 16'h005D; B = 16'h00CF; #100;
A = 16'h005D; B = 16'h00D0; #100;
A = 16'h005D; B = 16'h00D1; #100;
A = 16'h005D; B = 16'h00D2; #100;
A = 16'h005D; B = 16'h00D3; #100;
A = 16'h005D; B = 16'h00D4; #100;
A = 16'h005D; B = 16'h00D5; #100;
A = 16'h005D; B = 16'h00D6; #100;
A = 16'h005D; B = 16'h00D7; #100;
A = 16'h005D; B = 16'h00D8; #100;
A = 16'h005D; B = 16'h00D9; #100;
A = 16'h005D; B = 16'h00DA; #100;
A = 16'h005D; B = 16'h00DB; #100;
A = 16'h005D; B = 16'h00DC; #100;
A = 16'h005D; B = 16'h00DD; #100;
A = 16'h005D; B = 16'h00DE; #100;
A = 16'h005D; B = 16'h00DF; #100;
A = 16'h005D; B = 16'h00E0; #100;
A = 16'h005D; B = 16'h00E1; #100;
A = 16'h005D; B = 16'h00E2; #100;
A = 16'h005D; B = 16'h00E3; #100;
A = 16'h005D; B = 16'h00E4; #100;
A = 16'h005D; B = 16'h00E5; #100;
A = 16'h005D; B = 16'h00E6; #100;
A = 16'h005D; B = 16'h00E7; #100;
A = 16'h005D; B = 16'h00E8; #100;
A = 16'h005D; B = 16'h00E9; #100;
A = 16'h005D; B = 16'h00EA; #100;
A = 16'h005D; B = 16'h00EB; #100;
A = 16'h005D; B = 16'h00EC; #100;
A = 16'h005D; B = 16'h00ED; #100;
A = 16'h005D; B = 16'h00EE; #100;
A = 16'h005D; B = 16'h00EF; #100;
A = 16'h005D; B = 16'h00F0; #100;
A = 16'h005D; B = 16'h00F1; #100;
A = 16'h005D; B = 16'h00F2; #100;
A = 16'h005D; B = 16'h00F3; #100;
A = 16'h005D; B = 16'h00F4; #100;
A = 16'h005D; B = 16'h00F5; #100;
A = 16'h005D; B = 16'h00F6; #100;
A = 16'h005D; B = 16'h00F7; #100;
A = 16'h005D; B = 16'h00F8; #100;
A = 16'h005D; B = 16'h00F9; #100;
A = 16'h005D; B = 16'h00FA; #100;
A = 16'h005D; B = 16'h00FB; #100;
A = 16'h005D; B = 16'h00FC; #100;
A = 16'h005D; B = 16'h00FD; #100;
A = 16'h005D; B = 16'h00FE; #100;
A = 16'h005D; B = 16'h00FF; #100;
A = 16'h005E; B = 16'h000; #100;
A = 16'h005E; B = 16'h001; #100;
A = 16'h005E; B = 16'h002; #100;
A = 16'h005E; B = 16'h003; #100;
A = 16'h005E; B = 16'h004; #100;
A = 16'h005E; B = 16'h005; #100;
A = 16'h005E; B = 16'h006; #100;
A = 16'h005E; B = 16'h007; #100;
A = 16'h005E; B = 16'h008; #100;
A = 16'h005E; B = 16'h009; #100;
A = 16'h005E; B = 16'h00A; #100;
A = 16'h005E; B = 16'h00B; #100;
A = 16'h005E; B = 16'h00C; #100;
A = 16'h005E; B = 16'h00D; #100;
A = 16'h005E; B = 16'h00E; #100;
A = 16'h005E; B = 16'h00F; #100;
A = 16'h005E; B = 16'h0010; #100;
A = 16'h005E; B = 16'h0011; #100;
A = 16'h005E; B = 16'h0012; #100;
A = 16'h005E; B = 16'h0013; #100;
A = 16'h005E; B = 16'h0014; #100;
A = 16'h005E; B = 16'h0015; #100;
A = 16'h005E; B = 16'h0016; #100;
A = 16'h005E; B = 16'h0017; #100;
A = 16'h005E; B = 16'h0018; #100;
A = 16'h005E; B = 16'h0019; #100;
A = 16'h005E; B = 16'h001A; #100;
A = 16'h005E; B = 16'h001B; #100;
A = 16'h005E; B = 16'h001C; #100;
A = 16'h005E; B = 16'h001D; #100;
A = 16'h005E; B = 16'h001E; #100;
A = 16'h005E; B = 16'h001F; #100;
A = 16'h005E; B = 16'h0020; #100;
A = 16'h005E; B = 16'h0021; #100;
A = 16'h005E; B = 16'h0022; #100;
A = 16'h005E; B = 16'h0023; #100;
A = 16'h005E; B = 16'h0024; #100;
A = 16'h005E; B = 16'h0025; #100;
A = 16'h005E; B = 16'h0026; #100;
A = 16'h005E; B = 16'h0027; #100;
A = 16'h005E; B = 16'h0028; #100;
A = 16'h005E; B = 16'h0029; #100;
A = 16'h005E; B = 16'h002A; #100;
A = 16'h005E; B = 16'h002B; #100;
A = 16'h005E; B = 16'h002C; #100;
A = 16'h005E; B = 16'h002D; #100;
A = 16'h005E; B = 16'h002E; #100;
A = 16'h005E; B = 16'h002F; #100;
A = 16'h005E; B = 16'h0030; #100;
A = 16'h005E; B = 16'h0031; #100;
A = 16'h005E; B = 16'h0032; #100;
A = 16'h005E; B = 16'h0033; #100;
A = 16'h005E; B = 16'h0034; #100;
A = 16'h005E; B = 16'h0035; #100;
A = 16'h005E; B = 16'h0036; #100;
A = 16'h005E; B = 16'h0037; #100;
A = 16'h005E; B = 16'h0038; #100;
A = 16'h005E; B = 16'h0039; #100;
A = 16'h005E; B = 16'h003A; #100;
A = 16'h005E; B = 16'h003B; #100;
A = 16'h005E; B = 16'h003C; #100;
A = 16'h005E; B = 16'h003D; #100;
A = 16'h005E; B = 16'h003E; #100;
A = 16'h005E; B = 16'h003F; #100;
A = 16'h005E; B = 16'h0040; #100;
A = 16'h005E; B = 16'h0041; #100;
A = 16'h005E; B = 16'h0042; #100;
A = 16'h005E; B = 16'h0043; #100;
A = 16'h005E; B = 16'h0044; #100;
A = 16'h005E; B = 16'h0045; #100;
A = 16'h005E; B = 16'h0046; #100;
A = 16'h005E; B = 16'h0047; #100;
A = 16'h005E; B = 16'h0048; #100;
A = 16'h005E; B = 16'h0049; #100;
A = 16'h005E; B = 16'h004A; #100;
A = 16'h005E; B = 16'h004B; #100;
A = 16'h005E; B = 16'h004C; #100;
A = 16'h005E; B = 16'h004D; #100;
A = 16'h005E; B = 16'h004E; #100;
A = 16'h005E; B = 16'h004F; #100;
A = 16'h005E; B = 16'h0050; #100;
A = 16'h005E; B = 16'h0051; #100;
A = 16'h005E; B = 16'h0052; #100;
A = 16'h005E; B = 16'h0053; #100;
A = 16'h005E; B = 16'h0054; #100;
A = 16'h005E; B = 16'h0055; #100;
A = 16'h005E; B = 16'h0056; #100;
A = 16'h005E; B = 16'h0057; #100;
A = 16'h005E; B = 16'h0058; #100;
A = 16'h005E; B = 16'h0059; #100;
A = 16'h005E; B = 16'h005A; #100;
A = 16'h005E; B = 16'h005B; #100;
A = 16'h005E; B = 16'h005C; #100;
A = 16'h005E; B = 16'h005D; #100;
A = 16'h005E; B = 16'h005E; #100;
A = 16'h005E; B = 16'h005F; #100;
A = 16'h005E; B = 16'h0060; #100;
A = 16'h005E; B = 16'h0061; #100;
A = 16'h005E; B = 16'h0062; #100;
A = 16'h005E; B = 16'h0063; #100;
A = 16'h005E; B = 16'h0064; #100;
A = 16'h005E; B = 16'h0065; #100;
A = 16'h005E; B = 16'h0066; #100;
A = 16'h005E; B = 16'h0067; #100;
A = 16'h005E; B = 16'h0068; #100;
A = 16'h005E; B = 16'h0069; #100;
A = 16'h005E; B = 16'h006A; #100;
A = 16'h005E; B = 16'h006B; #100;
A = 16'h005E; B = 16'h006C; #100;
A = 16'h005E; B = 16'h006D; #100;
A = 16'h005E; B = 16'h006E; #100;
A = 16'h005E; B = 16'h006F; #100;
A = 16'h005E; B = 16'h0070; #100;
A = 16'h005E; B = 16'h0071; #100;
A = 16'h005E; B = 16'h0072; #100;
A = 16'h005E; B = 16'h0073; #100;
A = 16'h005E; B = 16'h0074; #100;
A = 16'h005E; B = 16'h0075; #100;
A = 16'h005E; B = 16'h0076; #100;
A = 16'h005E; B = 16'h0077; #100;
A = 16'h005E; B = 16'h0078; #100;
A = 16'h005E; B = 16'h0079; #100;
A = 16'h005E; B = 16'h007A; #100;
A = 16'h005E; B = 16'h007B; #100;
A = 16'h005E; B = 16'h007C; #100;
A = 16'h005E; B = 16'h007D; #100;
A = 16'h005E; B = 16'h007E; #100;
A = 16'h005E; B = 16'h007F; #100;
A = 16'h005E; B = 16'h0080; #100;
A = 16'h005E; B = 16'h0081; #100;
A = 16'h005E; B = 16'h0082; #100;
A = 16'h005E; B = 16'h0083; #100;
A = 16'h005E; B = 16'h0084; #100;
A = 16'h005E; B = 16'h0085; #100;
A = 16'h005E; B = 16'h0086; #100;
A = 16'h005E; B = 16'h0087; #100;
A = 16'h005E; B = 16'h0088; #100;
A = 16'h005E; B = 16'h0089; #100;
A = 16'h005E; B = 16'h008A; #100;
A = 16'h005E; B = 16'h008B; #100;
A = 16'h005E; B = 16'h008C; #100;
A = 16'h005E; B = 16'h008D; #100;
A = 16'h005E; B = 16'h008E; #100;
A = 16'h005E; B = 16'h008F; #100;
A = 16'h005E; B = 16'h0090; #100;
A = 16'h005E; B = 16'h0091; #100;
A = 16'h005E; B = 16'h0092; #100;
A = 16'h005E; B = 16'h0093; #100;
A = 16'h005E; B = 16'h0094; #100;
A = 16'h005E; B = 16'h0095; #100;
A = 16'h005E; B = 16'h0096; #100;
A = 16'h005E; B = 16'h0097; #100;
A = 16'h005E; B = 16'h0098; #100;
A = 16'h005E; B = 16'h0099; #100;
A = 16'h005E; B = 16'h009A; #100;
A = 16'h005E; B = 16'h009B; #100;
A = 16'h005E; B = 16'h009C; #100;
A = 16'h005E; B = 16'h009D; #100;
A = 16'h005E; B = 16'h009E; #100;
A = 16'h005E; B = 16'h009F; #100;
A = 16'h005E; B = 16'h00A0; #100;
A = 16'h005E; B = 16'h00A1; #100;
A = 16'h005E; B = 16'h00A2; #100;
A = 16'h005E; B = 16'h00A3; #100;
A = 16'h005E; B = 16'h00A4; #100;
A = 16'h005E; B = 16'h00A5; #100;
A = 16'h005E; B = 16'h00A6; #100;
A = 16'h005E; B = 16'h00A7; #100;
A = 16'h005E; B = 16'h00A8; #100;
A = 16'h005E; B = 16'h00A9; #100;
A = 16'h005E; B = 16'h00AA; #100;
A = 16'h005E; B = 16'h00AB; #100;
A = 16'h005E; B = 16'h00AC; #100;
A = 16'h005E; B = 16'h00AD; #100;
A = 16'h005E; B = 16'h00AE; #100;
A = 16'h005E; B = 16'h00AF; #100;
A = 16'h005E; B = 16'h00B0; #100;
A = 16'h005E; B = 16'h00B1; #100;
A = 16'h005E; B = 16'h00B2; #100;
A = 16'h005E; B = 16'h00B3; #100;
A = 16'h005E; B = 16'h00B4; #100;
A = 16'h005E; B = 16'h00B5; #100;
A = 16'h005E; B = 16'h00B6; #100;
A = 16'h005E; B = 16'h00B7; #100;
A = 16'h005E; B = 16'h00B8; #100;
A = 16'h005E; B = 16'h00B9; #100;
A = 16'h005E; B = 16'h00BA; #100;
A = 16'h005E; B = 16'h00BB; #100;
A = 16'h005E; B = 16'h00BC; #100;
A = 16'h005E; B = 16'h00BD; #100;
A = 16'h005E; B = 16'h00BE; #100;
A = 16'h005E; B = 16'h00BF; #100;
A = 16'h005E; B = 16'h00C0; #100;
A = 16'h005E; B = 16'h00C1; #100;
A = 16'h005E; B = 16'h00C2; #100;
A = 16'h005E; B = 16'h00C3; #100;
A = 16'h005E; B = 16'h00C4; #100;
A = 16'h005E; B = 16'h00C5; #100;
A = 16'h005E; B = 16'h00C6; #100;
A = 16'h005E; B = 16'h00C7; #100;
A = 16'h005E; B = 16'h00C8; #100;
A = 16'h005E; B = 16'h00C9; #100;
A = 16'h005E; B = 16'h00CA; #100;
A = 16'h005E; B = 16'h00CB; #100;
A = 16'h005E; B = 16'h00CC; #100;
A = 16'h005E; B = 16'h00CD; #100;
A = 16'h005E; B = 16'h00CE; #100;
A = 16'h005E; B = 16'h00CF; #100;
A = 16'h005E; B = 16'h00D0; #100;
A = 16'h005E; B = 16'h00D1; #100;
A = 16'h005E; B = 16'h00D2; #100;
A = 16'h005E; B = 16'h00D3; #100;
A = 16'h005E; B = 16'h00D4; #100;
A = 16'h005E; B = 16'h00D5; #100;
A = 16'h005E; B = 16'h00D6; #100;
A = 16'h005E; B = 16'h00D7; #100;
A = 16'h005E; B = 16'h00D8; #100;
A = 16'h005E; B = 16'h00D9; #100;
A = 16'h005E; B = 16'h00DA; #100;
A = 16'h005E; B = 16'h00DB; #100;
A = 16'h005E; B = 16'h00DC; #100;
A = 16'h005E; B = 16'h00DD; #100;
A = 16'h005E; B = 16'h00DE; #100;
A = 16'h005E; B = 16'h00DF; #100;
A = 16'h005E; B = 16'h00E0; #100;
A = 16'h005E; B = 16'h00E1; #100;
A = 16'h005E; B = 16'h00E2; #100;
A = 16'h005E; B = 16'h00E3; #100;
A = 16'h005E; B = 16'h00E4; #100;
A = 16'h005E; B = 16'h00E5; #100;
A = 16'h005E; B = 16'h00E6; #100;
A = 16'h005E; B = 16'h00E7; #100;
A = 16'h005E; B = 16'h00E8; #100;
A = 16'h005E; B = 16'h00E9; #100;
A = 16'h005E; B = 16'h00EA; #100;
A = 16'h005E; B = 16'h00EB; #100;
A = 16'h005E; B = 16'h00EC; #100;
A = 16'h005E; B = 16'h00ED; #100;
A = 16'h005E; B = 16'h00EE; #100;
A = 16'h005E; B = 16'h00EF; #100;
A = 16'h005E; B = 16'h00F0; #100;
A = 16'h005E; B = 16'h00F1; #100;
A = 16'h005E; B = 16'h00F2; #100;
A = 16'h005E; B = 16'h00F3; #100;
A = 16'h005E; B = 16'h00F4; #100;
A = 16'h005E; B = 16'h00F5; #100;
A = 16'h005E; B = 16'h00F6; #100;
A = 16'h005E; B = 16'h00F7; #100;
A = 16'h005E; B = 16'h00F8; #100;
A = 16'h005E; B = 16'h00F9; #100;
A = 16'h005E; B = 16'h00FA; #100;
A = 16'h005E; B = 16'h00FB; #100;
A = 16'h005E; B = 16'h00FC; #100;
A = 16'h005E; B = 16'h00FD; #100;
A = 16'h005E; B = 16'h00FE; #100;
A = 16'h005E; B = 16'h00FF; #100;
A = 16'h005F; B = 16'h000; #100;
A = 16'h005F; B = 16'h001; #100;
A = 16'h005F; B = 16'h002; #100;
A = 16'h005F; B = 16'h003; #100;
A = 16'h005F; B = 16'h004; #100;
A = 16'h005F; B = 16'h005; #100;
A = 16'h005F; B = 16'h006; #100;
A = 16'h005F; B = 16'h007; #100;
A = 16'h005F; B = 16'h008; #100;
A = 16'h005F; B = 16'h009; #100;
A = 16'h005F; B = 16'h00A; #100;
A = 16'h005F; B = 16'h00B; #100;
A = 16'h005F; B = 16'h00C; #100;
A = 16'h005F; B = 16'h00D; #100;
A = 16'h005F; B = 16'h00E; #100;
A = 16'h005F; B = 16'h00F; #100;
A = 16'h005F; B = 16'h0010; #100;
A = 16'h005F; B = 16'h0011; #100;
A = 16'h005F; B = 16'h0012; #100;
A = 16'h005F; B = 16'h0013; #100;
A = 16'h005F; B = 16'h0014; #100;
A = 16'h005F; B = 16'h0015; #100;
A = 16'h005F; B = 16'h0016; #100;
A = 16'h005F; B = 16'h0017; #100;
A = 16'h005F; B = 16'h0018; #100;
A = 16'h005F; B = 16'h0019; #100;
A = 16'h005F; B = 16'h001A; #100;
A = 16'h005F; B = 16'h001B; #100;
A = 16'h005F; B = 16'h001C; #100;
A = 16'h005F; B = 16'h001D; #100;
A = 16'h005F; B = 16'h001E; #100;
A = 16'h005F; B = 16'h001F; #100;
A = 16'h005F; B = 16'h0020; #100;
A = 16'h005F; B = 16'h0021; #100;
A = 16'h005F; B = 16'h0022; #100;
A = 16'h005F; B = 16'h0023; #100;
A = 16'h005F; B = 16'h0024; #100;
A = 16'h005F; B = 16'h0025; #100;
A = 16'h005F; B = 16'h0026; #100;
A = 16'h005F; B = 16'h0027; #100;
A = 16'h005F; B = 16'h0028; #100;
A = 16'h005F; B = 16'h0029; #100;
A = 16'h005F; B = 16'h002A; #100;
A = 16'h005F; B = 16'h002B; #100;
A = 16'h005F; B = 16'h002C; #100;
A = 16'h005F; B = 16'h002D; #100;
A = 16'h005F; B = 16'h002E; #100;
A = 16'h005F; B = 16'h002F; #100;
A = 16'h005F; B = 16'h0030; #100;
A = 16'h005F; B = 16'h0031; #100;
A = 16'h005F; B = 16'h0032; #100;
A = 16'h005F; B = 16'h0033; #100;
A = 16'h005F; B = 16'h0034; #100;
A = 16'h005F; B = 16'h0035; #100;
A = 16'h005F; B = 16'h0036; #100;
A = 16'h005F; B = 16'h0037; #100;
A = 16'h005F; B = 16'h0038; #100;
A = 16'h005F; B = 16'h0039; #100;
A = 16'h005F; B = 16'h003A; #100;
A = 16'h005F; B = 16'h003B; #100;
A = 16'h005F; B = 16'h003C; #100;
A = 16'h005F; B = 16'h003D; #100;
A = 16'h005F; B = 16'h003E; #100;
A = 16'h005F; B = 16'h003F; #100;
A = 16'h005F; B = 16'h0040; #100;
A = 16'h005F; B = 16'h0041; #100;
A = 16'h005F; B = 16'h0042; #100;
A = 16'h005F; B = 16'h0043; #100;
A = 16'h005F; B = 16'h0044; #100;
A = 16'h005F; B = 16'h0045; #100;
A = 16'h005F; B = 16'h0046; #100;
A = 16'h005F; B = 16'h0047; #100;
A = 16'h005F; B = 16'h0048; #100;
A = 16'h005F; B = 16'h0049; #100;
A = 16'h005F; B = 16'h004A; #100;
A = 16'h005F; B = 16'h004B; #100;
A = 16'h005F; B = 16'h004C; #100;
A = 16'h005F; B = 16'h004D; #100;
A = 16'h005F; B = 16'h004E; #100;
A = 16'h005F; B = 16'h004F; #100;
A = 16'h005F; B = 16'h0050; #100;
A = 16'h005F; B = 16'h0051; #100;
A = 16'h005F; B = 16'h0052; #100;
A = 16'h005F; B = 16'h0053; #100;
A = 16'h005F; B = 16'h0054; #100;
A = 16'h005F; B = 16'h0055; #100;
A = 16'h005F; B = 16'h0056; #100;
A = 16'h005F; B = 16'h0057; #100;
A = 16'h005F; B = 16'h0058; #100;
A = 16'h005F; B = 16'h0059; #100;
A = 16'h005F; B = 16'h005A; #100;
A = 16'h005F; B = 16'h005B; #100;
A = 16'h005F; B = 16'h005C; #100;
A = 16'h005F; B = 16'h005D; #100;
A = 16'h005F; B = 16'h005E; #100;
A = 16'h005F; B = 16'h005F; #100;
A = 16'h005F; B = 16'h0060; #100;
A = 16'h005F; B = 16'h0061; #100;
A = 16'h005F; B = 16'h0062; #100;
A = 16'h005F; B = 16'h0063; #100;
A = 16'h005F; B = 16'h0064; #100;
A = 16'h005F; B = 16'h0065; #100;
A = 16'h005F; B = 16'h0066; #100;
A = 16'h005F; B = 16'h0067; #100;
A = 16'h005F; B = 16'h0068; #100;
A = 16'h005F; B = 16'h0069; #100;
A = 16'h005F; B = 16'h006A; #100;
A = 16'h005F; B = 16'h006B; #100;
A = 16'h005F; B = 16'h006C; #100;
A = 16'h005F; B = 16'h006D; #100;
A = 16'h005F; B = 16'h006E; #100;
A = 16'h005F; B = 16'h006F; #100;
A = 16'h005F; B = 16'h0070; #100;
A = 16'h005F; B = 16'h0071; #100;
A = 16'h005F; B = 16'h0072; #100;
A = 16'h005F; B = 16'h0073; #100;
A = 16'h005F; B = 16'h0074; #100;
A = 16'h005F; B = 16'h0075; #100;
A = 16'h005F; B = 16'h0076; #100;
A = 16'h005F; B = 16'h0077; #100;
A = 16'h005F; B = 16'h0078; #100;
A = 16'h005F; B = 16'h0079; #100;
A = 16'h005F; B = 16'h007A; #100;
A = 16'h005F; B = 16'h007B; #100;
A = 16'h005F; B = 16'h007C; #100;
A = 16'h005F; B = 16'h007D; #100;
A = 16'h005F; B = 16'h007E; #100;
A = 16'h005F; B = 16'h007F; #100;
A = 16'h005F; B = 16'h0080; #100;
A = 16'h005F; B = 16'h0081; #100;
A = 16'h005F; B = 16'h0082; #100;
A = 16'h005F; B = 16'h0083; #100;
A = 16'h005F; B = 16'h0084; #100;
A = 16'h005F; B = 16'h0085; #100;
A = 16'h005F; B = 16'h0086; #100;
A = 16'h005F; B = 16'h0087; #100;
A = 16'h005F; B = 16'h0088; #100;
A = 16'h005F; B = 16'h0089; #100;
A = 16'h005F; B = 16'h008A; #100;
A = 16'h005F; B = 16'h008B; #100;
A = 16'h005F; B = 16'h008C; #100;
A = 16'h005F; B = 16'h008D; #100;
A = 16'h005F; B = 16'h008E; #100;
A = 16'h005F; B = 16'h008F; #100;
A = 16'h005F; B = 16'h0090; #100;
A = 16'h005F; B = 16'h0091; #100;
A = 16'h005F; B = 16'h0092; #100;
A = 16'h005F; B = 16'h0093; #100;
A = 16'h005F; B = 16'h0094; #100;
A = 16'h005F; B = 16'h0095; #100;
A = 16'h005F; B = 16'h0096; #100;
A = 16'h005F; B = 16'h0097; #100;
A = 16'h005F; B = 16'h0098; #100;
A = 16'h005F; B = 16'h0099; #100;
A = 16'h005F; B = 16'h009A; #100;
A = 16'h005F; B = 16'h009B; #100;
A = 16'h005F; B = 16'h009C; #100;
A = 16'h005F; B = 16'h009D; #100;
A = 16'h005F; B = 16'h009E; #100;
A = 16'h005F; B = 16'h009F; #100;
A = 16'h005F; B = 16'h00A0; #100;
A = 16'h005F; B = 16'h00A1; #100;
A = 16'h005F; B = 16'h00A2; #100;
A = 16'h005F; B = 16'h00A3; #100;
A = 16'h005F; B = 16'h00A4; #100;
A = 16'h005F; B = 16'h00A5; #100;
A = 16'h005F; B = 16'h00A6; #100;
A = 16'h005F; B = 16'h00A7; #100;
A = 16'h005F; B = 16'h00A8; #100;
A = 16'h005F; B = 16'h00A9; #100;
A = 16'h005F; B = 16'h00AA; #100;
A = 16'h005F; B = 16'h00AB; #100;
A = 16'h005F; B = 16'h00AC; #100;
A = 16'h005F; B = 16'h00AD; #100;
A = 16'h005F; B = 16'h00AE; #100;
A = 16'h005F; B = 16'h00AF; #100;
A = 16'h005F; B = 16'h00B0; #100;
A = 16'h005F; B = 16'h00B1; #100;
A = 16'h005F; B = 16'h00B2; #100;
A = 16'h005F; B = 16'h00B3; #100;
A = 16'h005F; B = 16'h00B4; #100;
A = 16'h005F; B = 16'h00B5; #100;
A = 16'h005F; B = 16'h00B6; #100;
A = 16'h005F; B = 16'h00B7; #100;
A = 16'h005F; B = 16'h00B8; #100;
A = 16'h005F; B = 16'h00B9; #100;
A = 16'h005F; B = 16'h00BA; #100;
A = 16'h005F; B = 16'h00BB; #100;
A = 16'h005F; B = 16'h00BC; #100;
A = 16'h005F; B = 16'h00BD; #100;
A = 16'h005F; B = 16'h00BE; #100;
A = 16'h005F; B = 16'h00BF; #100;
A = 16'h005F; B = 16'h00C0; #100;
A = 16'h005F; B = 16'h00C1; #100;
A = 16'h005F; B = 16'h00C2; #100;
A = 16'h005F; B = 16'h00C3; #100;
A = 16'h005F; B = 16'h00C4; #100;
A = 16'h005F; B = 16'h00C5; #100;
A = 16'h005F; B = 16'h00C6; #100;
A = 16'h005F; B = 16'h00C7; #100;
A = 16'h005F; B = 16'h00C8; #100;
A = 16'h005F; B = 16'h00C9; #100;
A = 16'h005F; B = 16'h00CA; #100;
A = 16'h005F; B = 16'h00CB; #100;
A = 16'h005F; B = 16'h00CC; #100;
A = 16'h005F; B = 16'h00CD; #100;
A = 16'h005F; B = 16'h00CE; #100;
A = 16'h005F; B = 16'h00CF; #100;
A = 16'h005F; B = 16'h00D0; #100;
A = 16'h005F; B = 16'h00D1; #100;
A = 16'h005F; B = 16'h00D2; #100;
A = 16'h005F; B = 16'h00D3; #100;
A = 16'h005F; B = 16'h00D4; #100;
A = 16'h005F; B = 16'h00D5; #100;
A = 16'h005F; B = 16'h00D6; #100;
A = 16'h005F; B = 16'h00D7; #100;
A = 16'h005F; B = 16'h00D8; #100;
A = 16'h005F; B = 16'h00D9; #100;
A = 16'h005F; B = 16'h00DA; #100;
A = 16'h005F; B = 16'h00DB; #100;
A = 16'h005F; B = 16'h00DC; #100;
A = 16'h005F; B = 16'h00DD; #100;
A = 16'h005F; B = 16'h00DE; #100;
A = 16'h005F; B = 16'h00DF; #100;
A = 16'h005F; B = 16'h00E0; #100;
A = 16'h005F; B = 16'h00E1; #100;
A = 16'h005F; B = 16'h00E2; #100;
A = 16'h005F; B = 16'h00E3; #100;
A = 16'h005F; B = 16'h00E4; #100;
A = 16'h005F; B = 16'h00E5; #100;
A = 16'h005F; B = 16'h00E6; #100;
A = 16'h005F; B = 16'h00E7; #100;
A = 16'h005F; B = 16'h00E8; #100;
A = 16'h005F; B = 16'h00E9; #100;
A = 16'h005F; B = 16'h00EA; #100;
A = 16'h005F; B = 16'h00EB; #100;
A = 16'h005F; B = 16'h00EC; #100;
A = 16'h005F; B = 16'h00ED; #100;
A = 16'h005F; B = 16'h00EE; #100;
A = 16'h005F; B = 16'h00EF; #100;
A = 16'h005F; B = 16'h00F0; #100;
A = 16'h005F; B = 16'h00F1; #100;
A = 16'h005F; B = 16'h00F2; #100;
A = 16'h005F; B = 16'h00F3; #100;
A = 16'h005F; B = 16'h00F4; #100;
A = 16'h005F; B = 16'h00F5; #100;
A = 16'h005F; B = 16'h00F6; #100;
A = 16'h005F; B = 16'h00F7; #100;
A = 16'h005F; B = 16'h00F8; #100;
A = 16'h005F; B = 16'h00F9; #100;
A = 16'h005F; B = 16'h00FA; #100;
A = 16'h005F; B = 16'h00FB; #100;
A = 16'h005F; B = 16'h00FC; #100;
A = 16'h005F; B = 16'h00FD; #100;
A = 16'h005F; B = 16'h00FE; #100;
A = 16'h005F; B = 16'h00FF; #100;
A = 16'h0060; B = 16'h000; #100;
A = 16'h0060; B = 16'h001; #100;
A = 16'h0060; B = 16'h002; #100;
A = 16'h0060; B = 16'h003; #100;
A = 16'h0060; B = 16'h004; #100;
A = 16'h0060; B = 16'h005; #100;
A = 16'h0060; B = 16'h006; #100;
A = 16'h0060; B = 16'h007; #100;
A = 16'h0060; B = 16'h008; #100;
A = 16'h0060; B = 16'h009; #100;
A = 16'h0060; B = 16'h00A; #100;
A = 16'h0060; B = 16'h00B; #100;
A = 16'h0060; B = 16'h00C; #100;
A = 16'h0060; B = 16'h00D; #100;
A = 16'h0060; B = 16'h00E; #100;
A = 16'h0060; B = 16'h00F; #100;
A = 16'h0060; B = 16'h0010; #100;
A = 16'h0060; B = 16'h0011; #100;
A = 16'h0060; B = 16'h0012; #100;
A = 16'h0060; B = 16'h0013; #100;
A = 16'h0060; B = 16'h0014; #100;
A = 16'h0060; B = 16'h0015; #100;
A = 16'h0060; B = 16'h0016; #100;
A = 16'h0060; B = 16'h0017; #100;
A = 16'h0060; B = 16'h0018; #100;
A = 16'h0060; B = 16'h0019; #100;
A = 16'h0060; B = 16'h001A; #100;
A = 16'h0060; B = 16'h001B; #100;
A = 16'h0060; B = 16'h001C; #100;
A = 16'h0060; B = 16'h001D; #100;
A = 16'h0060; B = 16'h001E; #100;
A = 16'h0060; B = 16'h001F; #100;
A = 16'h0060; B = 16'h0020; #100;
A = 16'h0060; B = 16'h0021; #100;
A = 16'h0060; B = 16'h0022; #100;
A = 16'h0060; B = 16'h0023; #100;
A = 16'h0060; B = 16'h0024; #100;
A = 16'h0060; B = 16'h0025; #100;
A = 16'h0060; B = 16'h0026; #100;
A = 16'h0060; B = 16'h0027; #100;
A = 16'h0060; B = 16'h0028; #100;
A = 16'h0060; B = 16'h0029; #100;
A = 16'h0060; B = 16'h002A; #100;
A = 16'h0060; B = 16'h002B; #100;
A = 16'h0060; B = 16'h002C; #100;
A = 16'h0060; B = 16'h002D; #100;
A = 16'h0060; B = 16'h002E; #100;
A = 16'h0060; B = 16'h002F; #100;
A = 16'h0060; B = 16'h0030; #100;
A = 16'h0060; B = 16'h0031; #100;
A = 16'h0060; B = 16'h0032; #100;
A = 16'h0060; B = 16'h0033; #100;
A = 16'h0060; B = 16'h0034; #100;
A = 16'h0060; B = 16'h0035; #100;
A = 16'h0060; B = 16'h0036; #100;
A = 16'h0060; B = 16'h0037; #100;
A = 16'h0060; B = 16'h0038; #100;
A = 16'h0060; B = 16'h0039; #100;
A = 16'h0060; B = 16'h003A; #100;
A = 16'h0060; B = 16'h003B; #100;
A = 16'h0060; B = 16'h003C; #100;
A = 16'h0060; B = 16'h003D; #100;
A = 16'h0060; B = 16'h003E; #100;
A = 16'h0060; B = 16'h003F; #100;
A = 16'h0060; B = 16'h0040; #100;
A = 16'h0060; B = 16'h0041; #100;
A = 16'h0060; B = 16'h0042; #100;
A = 16'h0060; B = 16'h0043; #100;
A = 16'h0060; B = 16'h0044; #100;
A = 16'h0060; B = 16'h0045; #100;
A = 16'h0060; B = 16'h0046; #100;
A = 16'h0060; B = 16'h0047; #100;
A = 16'h0060; B = 16'h0048; #100;
A = 16'h0060; B = 16'h0049; #100;
A = 16'h0060; B = 16'h004A; #100;
A = 16'h0060; B = 16'h004B; #100;
A = 16'h0060; B = 16'h004C; #100;
A = 16'h0060; B = 16'h004D; #100;
A = 16'h0060; B = 16'h004E; #100;
A = 16'h0060; B = 16'h004F; #100;
A = 16'h0060; B = 16'h0050; #100;
A = 16'h0060; B = 16'h0051; #100;
A = 16'h0060; B = 16'h0052; #100;
A = 16'h0060; B = 16'h0053; #100;
A = 16'h0060; B = 16'h0054; #100;
A = 16'h0060; B = 16'h0055; #100;
A = 16'h0060; B = 16'h0056; #100;
A = 16'h0060; B = 16'h0057; #100;
A = 16'h0060; B = 16'h0058; #100;
A = 16'h0060; B = 16'h0059; #100;
A = 16'h0060; B = 16'h005A; #100;
A = 16'h0060; B = 16'h005B; #100;
A = 16'h0060; B = 16'h005C; #100;
A = 16'h0060; B = 16'h005D; #100;
A = 16'h0060; B = 16'h005E; #100;
A = 16'h0060; B = 16'h005F; #100;
A = 16'h0060; B = 16'h0060; #100;
A = 16'h0060; B = 16'h0061; #100;
A = 16'h0060; B = 16'h0062; #100;
A = 16'h0060; B = 16'h0063; #100;
A = 16'h0060; B = 16'h0064; #100;
A = 16'h0060; B = 16'h0065; #100;
A = 16'h0060; B = 16'h0066; #100;
A = 16'h0060; B = 16'h0067; #100;
A = 16'h0060; B = 16'h0068; #100;
A = 16'h0060; B = 16'h0069; #100;
A = 16'h0060; B = 16'h006A; #100;
A = 16'h0060; B = 16'h006B; #100;
A = 16'h0060; B = 16'h006C; #100;
A = 16'h0060; B = 16'h006D; #100;
A = 16'h0060; B = 16'h006E; #100;
A = 16'h0060; B = 16'h006F; #100;
A = 16'h0060; B = 16'h0070; #100;
A = 16'h0060; B = 16'h0071; #100;
A = 16'h0060; B = 16'h0072; #100;
A = 16'h0060; B = 16'h0073; #100;
A = 16'h0060; B = 16'h0074; #100;
A = 16'h0060; B = 16'h0075; #100;
A = 16'h0060; B = 16'h0076; #100;
A = 16'h0060; B = 16'h0077; #100;
A = 16'h0060; B = 16'h0078; #100;
A = 16'h0060; B = 16'h0079; #100;
A = 16'h0060; B = 16'h007A; #100;
A = 16'h0060; B = 16'h007B; #100;
A = 16'h0060; B = 16'h007C; #100;
A = 16'h0060; B = 16'h007D; #100;
A = 16'h0060; B = 16'h007E; #100;
A = 16'h0060; B = 16'h007F; #100;
A = 16'h0060; B = 16'h0080; #100;
A = 16'h0060; B = 16'h0081; #100;
A = 16'h0060; B = 16'h0082; #100;
A = 16'h0060; B = 16'h0083; #100;
A = 16'h0060; B = 16'h0084; #100;
A = 16'h0060; B = 16'h0085; #100;
A = 16'h0060; B = 16'h0086; #100;
A = 16'h0060; B = 16'h0087; #100;
A = 16'h0060; B = 16'h0088; #100;
A = 16'h0060; B = 16'h0089; #100;
A = 16'h0060; B = 16'h008A; #100;
A = 16'h0060; B = 16'h008B; #100;
A = 16'h0060; B = 16'h008C; #100;
A = 16'h0060; B = 16'h008D; #100;
A = 16'h0060; B = 16'h008E; #100;
A = 16'h0060; B = 16'h008F; #100;
A = 16'h0060; B = 16'h0090; #100;
A = 16'h0060; B = 16'h0091; #100;
A = 16'h0060; B = 16'h0092; #100;
A = 16'h0060; B = 16'h0093; #100;
A = 16'h0060; B = 16'h0094; #100;
A = 16'h0060; B = 16'h0095; #100;
A = 16'h0060; B = 16'h0096; #100;
A = 16'h0060; B = 16'h0097; #100;
A = 16'h0060; B = 16'h0098; #100;
A = 16'h0060; B = 16'h0099; #100;
A = 16'h0060; B = 16'h009A; #100;
A = 16'h0060; B = 16'h009B; #100;
A = 16'h0060; B = 16'h009C; #100;
A = 16'h0060; B = 16'h009D; #100;
A = 16'h0060; B = 16'h009E; #100;
A = 16'h0060; B = 16'h009F; #100;
A = 16'h0060; B = 16'h00A0; #100;
A = 16'h0060; B = 16'h00A1; #100;
A = 16'h0060; B = 16'h00A2; #100;
A = 16'h0060; B = 16'h00A3; #100;
A = 16'h0060; B = 16'h00A4; #100;
A = 16'h0060; B = 16'h00A5; #100;
A = 16'h0060; B = 16'h00A6; #100;
A = 16'h0060; B = 16'h00A7; #100;
A = 16'h0060; B = 16'h00A8; #100;
A = 16'h0060; B = 16'h00A9; #100;
A = 16'h0060; B = 16'h00AA; #100;
A = 16'h0060; B = 16'h00AB; #100;
A = 16'h0060; B = 16'h00AC; #100;
A = 16'h0060; B = 16'h00AD; #100;
A = 16'h0060; B = 16'h00AE; #100;
A = 16'h0060; B = 16'h00AF; #100;
A = 16'h0060; B = 16'h00B0; #100;
A = 16'h0060; B = 16'h00B1; #100;
A = 16'h0060; B = 16'h00B2; #100;
A = 16'h0060; B = 16'h00B3; #100;
A = 16'h0060; B = 16'h00B4; #100;
A = 16'h0060; B = 16'h00B5; #100;
A = 16'h0060; B = 16'h00B6; #100;
A = 16'h0060; B = 16'h00B7; #100;
A = 16'h0060; B = 16'h00B8; #100;
A = 16'h0060; B = 16'h00B9; #100;
A = 16'h0060; B = 16'h00BA; #100;
A = 16'h0060; B = 16'h00BB; #100;
A = 16'h0060; B = 16'h00BC; #100;
A = 16'h0060; B = 16'h00BD; #100;
A = 16'h0060; B = 16'h00BE; #100;
A = 16'h0060; B = 16'h00BF; #100;
A = 16'h0060; B = 16'h00C0; #100;
A = 16'h0060; B = 16'h00C1; #100;
A = 16'h0060; B = 16'h00C2; #100;
A = 16'h0060; B = 16'h00C3; #100;
A = 16'h0060; B = 16'h00C4; #100;
A = 16'h0060; B = 16'h00C5; #100;
A = 16'h0060; B = 16'h00C6; #100;
A = 16'h0060; B = 16'h00C7; #100;
A = 16'h0060; B = 16'h00C8; #100;
A = 16'h0060; B = 16'h00C9; #100;
A = 16'h0060; B = 16'h00CA; #100;
A = 16'h0060; B = 16'h00CB; #100;
A = 16'h0060; B = 16'h00CC; #100;
A = 16'h0060; B = 16'h00CD; #100;
A = 16'h0060; B = 16'h00CE; #100;
A = 16'h0060; B = 16'h00CF; #100;
A = 16'h0060; B = 16'h00D0; #100;
A = 16'h0060; B = 16'h00D1; #100;
A = 16'h0060; B = 16'h00D2; #100;
A = 16'h0060; B = 16'h00D3; #100;
A = 16'h0060; B = 16'h00D4; #100;
A = 16'h0060; B = 16'h00D5; #100;
A = 16'h0060; B = 16'h00D6; #100;
A = 16'h0060; B = 16'h00D7; #100;
A = 16'h0060; B = 16'h00D8; #100;
A = 16'h0060; B = 16'h00D9; #100;
A = 16'h0060; B = 16'h00DA; #100;
A = 16'h0060; B = 16'h00DB; #100;
A = 16'h0060; B = 16'h00DC; #100;
A = 16'h0060; B = 16'h00DD; #100;
A = 16'h0060; B = 16'h00DE; #100;
A = 16'h0060; B = 16'h00DF; #100;
A = 16'h0060; B = 16'h00E0; #100;
A = 16'h0060; B = 16'h00E1; #100;
A = 16'h0060; B = 16'h00E2; #100;
A = 16'h0060; B = 16'h00E3; #100;
A = 16'h0060; B = 16'h00E4; #100;
A = 16'h0060; B = 16'h00E5; #100;
A = 16'h0060; B = 16'h00E6; #100;
A = 16'h0060; B = 16'h00E7; #100;
A = 16'h0060; B = 16'h00E8; #100;
A = 16'h0060; B = 16'h00E9; #100;
A = 16'h0060; B = 16'h00EA; #100;
A = 16'h0060; B = 16'h00EB; #100;
A = 16'h0060; B = 16'h00EC; #100;
A = 16'h0060; B = 16'h00ED; #100;
A = 16'h0060; B = 16'h00EE; #100;
A = 16'h0060; B = 16'h00EF; #100;
A = 16'h0060; B = 16'h00F0; #100;
A = 16'h0060; B = 16'h00F1; #100;
A = 16'h0060; B = 16'h00F2; #100;
A = 16'h0060; B = 16'h00F3; #100;
A = 16'h0060; B = 16'h00F4; #100;
A = 16'h0060; B = 16'h00F5; #100;
A = 16'h0060; B = 16'h00F6; #100;
A = 16'h0060; B = 16'h00F7; #100;
A = 16'h0060; B = 16'h00F8; #100;
A = 16'h0060; B = 16'h00F9; #100;
A = 16'h0060; B = 16'h00FA; #100;
A = 16'h0060; B = 16'h00FB; #100;
A = 16'h0060; B = 16'h00FC; #100;
A = 16'h0060; B = 16'h00FD; #100;
A = 16'h0060; B = 16'h00FE; #100;
A = 16'h0060; B = 16'h00FF; #100;
A = 16'h0061; B = 16'h000; #100;
A = 16'h0061; B = 16'h001; #100;
A = 16'h0061; B = 16'h002; #100;
A = 16'h0061; B = 16'h003; #100;
A = 16'h0061; B = 16'h004; #100;
A = 16'h0061; B = 16'h005; #100;
A = 16'h0061; B = 16'h006; #100;
A = 16'h0061; B = 16'h007; #100;
A = 16'h0061; B = 16'h008; #100;
A = 16'h0061; B = 16'h009; #100;
A = 16'h0061; B = 16'h00A; #100;
A = 16'h0061; B = 16'h00B; #100;
A = 16'h0061; B = 16'h00C; #100;
A = 16'h0061; B = 16'h00D; #100;
A = 16'h0061; B = 16'h00E; #100;
A = 16'h0061; B = 16'h00F; #100;
A = 16'h0061; B = 16'h0010; #100;
A = 16'h0061; B = 16'h0011; #100;
A = 16'h0061; B = 16'h0012; #100;
A = 16'h0061; B = 16'h0013; #100;
A = 16'h0061; B = 16'h0014; #100;
A = 16'h0061; B = 16'h0015; #100;
A = 16'h0061; B = 16'h0016; #100;
A = 16'h0061; B = 16'h0017; #100;
A = 16'h0061; B = 16'h0018; #100;
A = 16'h0061; B = 16'h0019; #100;
A = 16'h0061; B = 16'h001A; #100;
A = 16'h0061; B = 16'h001B; #100;
A = 16'h0061; B = 16'h001C; #100;
A = 16'h0061; B = 16'h001D; #100;
A = 16'h0061; B = 16'h001E; #100;
A = 16'h0061; B = 16'h001F; #100;
A = 16'h0061; B = 16'h0020; #100;
A = 16'h0061; B = 16'h0021; #100;
A = 16'h0061; B = 16'h0022; #100;
A = 16'h0061; B = 16'h0023; #100;
A = 16'h0061; B = 16'h0024; #100;
A = 16'h0061; B = 16'h0025; #100;
A = 16'h0061; B = 16'h0026; #100;
A = 16'h0061; B = 16'h0027; #100;
A = 16'h0061; B = 16'h0028; #100;
A = 16'h0061; B = 16'h0029; #100;
A = 16'h0061; B = 16'h002A; #100;
A = 16'h0061; B = 16'h002B; #100;
A = 16'h0061; B = 16'h002C; #100;
A = 16'h0061; B = 16'h002D; #100;
A = 16'h0061; B = 16'h002E; #100;
A = 16'h0061; B = 16'h002F; #100;
A = 16'h0061; B = 16'h0030; #100;
A = 16'h0061; B = 16'h0031; #100;
A = 16'h0061; B = 16'h0032; #100;
A = 16'h0061; B = 16'h0033; #100;
A = 16'h0061; B = 16'h0034; #100;
A = 16'h0061; B = 16'h0035; #100;
A = 16'h0061; B = 16'h0036; #100;
A = 16'h0061; B = 16'h0037; #100;
A = 16'h0061; B = 16'h0038; #100;
A = 16'h0061; B = 16'h0039; #100;
A = 16'h0061; B = 16'h003A; #100;
A = 16'h0061; B = 16'h003B; #100;
A = 16'h0061; B = 16'h003C; #100;
A = 16'h0061; B = 16'h003D; #100;
A = 16'h0061; B = 16'h003E; #100;
A = 16'h0061; B = 16'h003F; #100;
A = 16'h0061; B = 16'h0040; #100;
A = 16'h0061; B = 16'h0041; #100;
A = 16'h0061; B = 16'h0042; #100;
A = 16'h0061; B = 16'h0043; #100;
A = 16'h0061; B = 16'h0044; #100;
A = 16'h0061; B = 16'h0045; #100;
A = 16'h0061; B = 16'h0046; #100;
A = 16'h0061; B = 16'h0047; #100;
A = 16'h0061; B = 16'h0048; #100;
A = 16'h0061; B = 16'h0049; #100;
A = 16'h0061; B = 16'h004A; #100;
A = 16'h0061; B = 16'h004B; #100;
A = 16'h0061; B = 16'h004C; #100;
A = 16'h0061; B = 16'h004D; #100;
A = 16'h0061; B = 16'h004E; #100;
A = 16'h0061; B = 16'h004F; #100;
A = 16'h0061; B = 16'h0050; #100;
A = 16'h0061; B = 16'h0051; #100;
A = 16'h0061; B = 16'h0052; #100;
A = 16'h0061; B = 16'h0053; #100;
A = 16'h0061; B = 16'h0054; #100;
A = 16'h0061; B = 16'h0055; #100;
A = 16'h0061; B = 16'h0056; #100;
A = 16'h0061; B = 16'h0057; #100;
A = 16'h0061; B = 16'h0058; #100;
A = 16'h0061; B = 16'h0059; #100;
A = 16'h0061; B = 16'h005A; #100;
A = 16'h0061; B = 16'h005B; #100;
A = 16'h0061; B = 16'h005C; #100;
A = 16'h0061; B = 16'h005D; #100;
A = 16'h0061; B = 16'h005E; #100;
A = 16'h0061; B = 16'h005F; #100;
A = 16'h0061; B = 16'h0060; #100;
A = 16'h0061; B = 16'h0061; #100;
A = 16'h0061; B = 16'h0062; #100;
A = 16'h0061; B = 16'h0063; #100;
A = 16'h0061; B = 16'h0064; #100;
A = 16'h0061; B = 16'h0065; #100;
A = 16'h0061; B = 16'h0066; #100;
A = 16'h0061; B = 16'h0067; #100;
A = 16'h0061; B = 16'h0068; #100;
A = 16'h0061; B = 16'h0069; #100;
A = 16'h0061; B = 16'h006A; #100;
A = 16'h0061; B = 16'h006B; #100;
A = 16'h0061; B = 16'h006C; #100;
A = 16'h0061; B = 16'h006D; #100;
A = 16'h0061; B = 16'h006E; #100;
A = 16'h0061; B = 16'h006F; #100;
A = 16'h0061; B = 16'h0070; #100;
A = 16'h0061; B = 16'h0071; #100;
A = 16'h0061; B = 16'h0072; #100;
A = 16'h0061; B = 16'h0073; #100;
A = 16'h0061; B = 16'h0074; #100;
A = 16'h0061; B = 16'h0075; #100;
A = 16'h0061; B = 16'h0076; #100;
A = 16'h0061; B = 16'h0077; #100;
A = 16'h0061; B = 16'h0078; #100;
A = 16'h0061; B = 16'h0079; #100;
A = 16'h0061; B = 16'h007A; #100;
A = 16'h0061; B = 16'h007B; #100;
A = 16'h0061; B = 16'h007C; #100;
A = 16'h0061; B = 16'h007D; #100;
A = 16'h0061; B = 16'h007E; #100;
A = 16'h0061; B = 16'h007F; #100;
A = 16'h0061; B = 16'h0080; #100;
A = 16'h0061; B = 16'h0081; #100;
A = 16'h0061; B = 16'h0082; #100;
A = 16'h0061; B = 16'h0083; #100;
A = 16'h0061; B = 16'h0084; #100;
A = 16'h0061; B = 16'h0085; #100;
A = 16'h0061; B = 16'h0086; #100;
A = 16'h0061; B = 16'h0087; #100;
A = 16'h0061; B = 16'h0088; #100;
A = 16'h0061; B = 16'h0089; #100;
A = 16'h0061; B = 16'h008A; #100;
A = 16'h0061; B = 16'h008B; #100;
A = 16'h0061; B = 16'h008C; #100;
A = 16'h0061; B = 16'h008D; #100;
A = 16'h0061; B = 16'h008E; #100;
A = 16'h0061; B = 16'h008F; #100;
A = 16'h0061; B = 16'h0090; #100;
A = 16'h0061; B = 16'h0091; #100;
A = 16'h0061; B = 16'h0092; #100;
A = 16'h0061; B = 16'h0093; #100;
A = 16'h0061; B = 16'h0094; #100;
A = 16'h0061; B = 16'h0095; #100;
A = 16'h0061; B = 16'h0096; #100;
A = 16'h0061; B = 16'h0097; #100;
A = 16'h0061; B = 16'h0098; #100;
A = 16'h0061; B = 16'h0099; #100;
A = 16'h0061; B = 16'h009A; #100;
A = 16'h0061; B = 16'h009B; #100;
A = 16'h0061; B = 16'h009C; #100;
A = 16'h0061; B = 16'h009D; #100;
A = 16'h0061; B = 16'h009E; #100;
A = 16'h0061; B = 16'h009F; #100;
A = 16'h0061; B = 16'h00A0; #100;
A = 16'h0061; B = 16'h00A1; #100;
A = 16'h0061; B = 16'h00A2; #100;
A = 16'h0061; B = 16'h00A3; #100;
A = 16'h0061; B = 16'h00A4; #100;
A = 16'h0061; B = 16'h00A5; #100;
A = 16'h0061; B = 16'h00A6; #100;
A = 16'h0061; B = 16'h00A7; #100;
A = 16'h0061; B = 16'h00A8; #100;
A = 16'h0061; B = 16'h00A9; #100;
A = 16'h0061; B = 16'h00AA; #100;
A = 16'h0061; B = 16'h00AB; #100;
A = 16'h0061; B = 16'h00AC; #100;
A = 16'h0061; B = 16'h00AD; #100;
A = 16'h0061; B = 16'h00AE; #100;
A = 16'h0061; B = 16'h00AF; #100;
A = 16'h0061; B = 16'h00B0; #100;
A = 16'h0061; B = 16'h00B1; #100;
A = 16'h0061; B = 16'h00B2; #100;
A = 16'h0061; B = 16'h00B3; #100;
A = 16'h0061; B = 16'h00B4; #100;
A = 16'h0061; B = 16'h00B5; #100;
A = 16'h0061; B = 16'h00B6; #100;
A = 16'h0061; B = 16'h00B7; #100;
A = 16'h0061; B = 16'h00B8; #100;
A = 16'h0061; B = 16'h00B9; #100;
A = 16'h0061; B = 16'h00BA; #100;
A = 16'h0061; B = 16'h00BB; #100;
A = 16'h0061; B = 16'h00BC; #100;
A = 16'h0061; B = 16'h00BD; #100;
A = 16'h0061; B = 16'h00BE; #100;
A = 16'h0061; B = 16'h00BF; #100;
A = 16'h0061; B = 16'h00C0; #100;
A = 16'h0061; B = 16'h00C1; #100;
A = 16'h0061; B = 16'h00C2; #100;
A = 16'h0061; B = 16'h00C3; #100;
A = 16'h0061; B = 16'h00C4; #100;
A = 16'h0061; B = 16'h00C5; #100;
A = 16'h0061; B = 16'h00C6; #100;
A = 16'h0061; B = 16'h00C7; #100;
A = 16'h0061; B = 16'h00C8; #100;
A = 16'h0061; B = 16'h00C9; #100;
A = 16'h0061; B = 16'h00CA; #100;
A = 16'h0061; B = 16'h00CB; #100;
A = 16'h0061; B = 16'h00CC; #100;
A = 16'h0061; B = 16'h00CD; #100;
A = 16'h0061; B = 16'h00CE; #100;
A = 16'h0061; B = 16'h00CF; #100;
A = 16'h0061; B = 16'h00D0; #100;
A = 16'h0061; B = 16'h00D1; #100;
A = 16'h0061; B = 16'h00D2; #100;
A = 16'h0061; B = 16'h00D3; #100;
A = 16'h0061; B = 16'h00D4; #100;
A = 16'h0061; B = 16'h00D5; #100;
A = 16'h0061; B = 16'h00D6; #100;
A = 16'h0061; B = 16'h00D7; #100;
A = 16'h0061; B = 16'h00D8; #100;
A = 16'h0061; B = 16'h00D9; #100;
A = 16'h0061; B = 16'h00DA; #100;
A = 16'h0061; B = 16'h00DB; #100;
A = 16'h0061; B = 16'h00DC; #100;
A = 16'h0061; B = 16'h00DD; #100;
A = 16'h0061; B = 16'h00DE; #100;
A = 16'h0061; B = 16'h00DF; #100;
A = 16'h0061; B = 16'h00E0; #100;
A = 16'h0061; B = 16'h00E1; #100;
A = 16'h0061; B = 16'h00E2; #100;
A = 16'h0061; B = 16'h00E3; #100;
A = 16'h0061; B = 16'h00E4; #100;
A = 16'h0061; B = 16'h00E5; #100;
A = 16'h0061; B = 16'h00E6; #100;
A = 16'h0061; B = 16'h00E7; #100;
A = 16'h0061; B = 16'h00E8; #100;
A = 16'h0061; B = 16'h00E9; #100;
A = 16'h0061; B = 16'h00EA; #100;
A = 16'h0061; B = 16'h00EB; #100;
A = 16'h0061; B = 16'h00EC; #100;
A = 16'h0061; B = 16'h00ED; #100;
A = 16'h0061; B = 16'h00EE; #100;
A = 16'h0061; B = 16'h00EF; #100;
A = 16'h0061; B = 16'h00F0; #100;
A = 16'h0061; B = 16'h00F1; #100;
A = 16'h0061; B = 16'h00F2; #100;
A = 16'h0061; B = 16'h00F3; #100;
A = 16'h0061; B = 16'h00F4; #100;
A = 16'h0061; B = 16'h00F5; #100;
A = 16'h0061; B = 16'h00F6; #100;
A = 16'h0061; B = 16'h00F7; #100;
A = 16'h0061; B = 16'h00F8; #100;
A = 16'h0061; B = 16'h00F9; #100;
A = 16'h0061; B = 16'h00FA; #100;
A = 16'h0061; B = 16'h00FB; #100;
A = 16'h0061; B = 16'h00FC; #100;
A = 16'h0061; B = 16'h00FD; #100;
A = 16'h0061; B = 16'h00FE; #100;
A = 16'h0061; B = 16'h00FF; #100;
A = 16'h0062; B = 16'h000; #100;
A = 16'h0062; B = 16'h001; #100;
A = 16'h0062; B = 16'h002; #100;
A = 16'h0062; B = 16'h003; #100;
A = 16'h0062; B = 16'h004; #100;
A = 16'h0062; B = 16'h005; #100;
A = 16'h0062; B = 16'h006; #100;
A = 16'h0062; B = 16'h007; #100;
A = 16'h0062; B = 16'h008; #100;
A = 16'h0062; B = 16'h009; #100;
A = 16'h0062; B = 16'h00A; #100;
A = 16'h0062; B = 16'h00B; #100;
A = 16'h0062; B = 16'h00C; #100;
A = 16'h0062; B = 16'h00D; #100;
A = 16'h0062; B = 16'h00E; #100;
A = 16'h0062; B = 16'h00F; #100;
A = 16'h0062; B = 16'h0010; #100;
A = 16'h0062; B = 16'h0011; #100;
A = 16'h0062; B = 16'h0012; #100;
A = 16'h0062; B = 16'h0013; #100;
A = 16'h0062; B = 16'h0014; #100;
A = 16'h0062; B = 16'h0015; #100;
A = 16'h0062; B = 16'h0016; #100;
A = 16'h0062; B = 16'h0017; #100;
A = 16'h0062; B = 16'h0018; #100;
A = 16'h0062; B = 16'h0019; #100;
A = 16'h0062; B = 16'h001A; #100;
A = 16'h0062; B = 16'h001B; #100;
A = 16'h0062; B = 16'h001C; #100;
A = 16'h0062; B = 16'h001D; #100;
A = 16'h0062; B = 16'h001E; #100;
A = 16'h0062; B = 16'h001F; #100;
A = 16'h0062; B = 16'h0020; #100;
A = 16'h0062; B = 16'h0021; #100;
A = 16'h0062; B = 16'h0022; #100;
A = 16'h0062; B = 16'h0023; #100;
A = 16'h0062; B = 16'h0024; #100;
A = 16'h0062; B = 16'h0025; #100;
A = 16'h0062; B = 16'h0026; #100;
A = 16'h0062; B = 16'h0027; #100;
A = 16'h0062; B = 16'h0028; #100;
A = 16'h0062; B = 16'h0029; #100;
A = 16'h0062; B = 16'h002A; #100;
A = 16'h0062; B = 16'h002B; #100;
A = 16'h0062; B = 16'h002C; #100;
A = 16'h0062; B = 16'h002D; #100;
A = 16'h0062; B = 16'h002E; #100;
A = 16'h0062; B = 16'h002F; #100;
A = 16'h0062; B = 16'h0030; #100;
A = 16'h0062; B = 16'h0031; #100;
A = 16'h0062; B = 16'h0032; #100;
A = 16'h0062; B = 16'h0033; #100;
A = 16'h0062; B = 16'h0034; #100;
A = 16'h0062; B = 16'h0035; #100;
A = 16'h0062; B = 16'h0036; #100;
A = 16'h0062; B = 16'h0037; #100;
A = 16'h0062; B = 16'h0038; #100;
A = 16'h0062; B = 16'h0039; #100;
A = 16'h0062; B = 16'h003A; #100;
A = 16'h0062; B = 16'h003B; #100;
A = 16'h0062; B = 16'h003C; #100;
A = 16'h0062; B = 16'h003D; #100;
A = 16'h0062; B = 16'h003E; #100;
A = 16'h0062; B = 16'h003F; #100;
A = 16'h0062; B = 16'h0040; #100;
A = 16'h0062; B = 16'h0041; #100;
A = 16'h0062; B = 16'h0042; #100;
A = 16'h0062; B = 16'h0043; #100;
A = 16'h0062; B = 16'h0044; #100;
A = 16'h0062; B = 16'h0045; #100;
A = 16'h0062; B = 16'h0046; #100;
A = 16'h0062; B = 16'h0047; #100;
A = 16'h0062; B = 16'h0048; #100;
A = 16'h0062; B = 16'h0049; #100;
A = 16'h0062; B = 16'h004A; #100;
A = 16'h0062; B = 16'h004B; #100;
A = 16'h0062; B = 16'h004C; #100;
A = 16'h0062; B = 16'h004D; #100;
A = 16'h0062; B = 16'h004E; #100;
A = 16'h0062; B = 16'h004F; #100;
A = 16'h0062; B = 16'h0050; #100;
A = 16'h0062; B = 16'h0051; #100;
A = 16'h0062; B = 16'h0052; #100;
A = 16'h0062; B = 16'h0053; #100;
A = 16'h0062; B = 16'h0054; #100;
A = 16'h0062; B = 16'h0055; #100;
A = 16'h0062; B = 16'h0056; #100;
A = 16'h0062; B = 16'h0057; #100;
A = 16'h0062; B = 16'h0058; #100;
A = 16'h0062; B = 16'h0059; #100;
A = 16'h0062; B = 16'h005A; #100;
A = 16'h0062; B = 16'h005B; #100;
A = 16'h0062; B = 16'h005C; #100;
A = 16'h0062; B = 16'h005D; #100;
A = 16'h0062; B = 16'h005E; #100;
A = 16'h0062; B = 16'h005F; #100;
A = 16'h0062; B = 16'h0060; #100;
A = 16'h0062; B = 16'h0061; #100;
A = 16'h0062; B = 16'h0062; #100;
A = 16'h0062; B = 16'h0063; #100;
A = 16'h0062; B = 16'h0064; #100;
A = 16'h0062; B = 16'h0065; #100;
A = 16'h0062; B = 16'h0066; #100;
A = 16'h0062; B = 16'h0067; #100;
A = 16'h0062; B = 16'h0068; #100;
A = 16'h0062; B = 16'h0069; #100;
A = 16'h0062; B = 16'h006A; #100;
A = 16'h0062; B = 16'h006B; #100;
A = 16'h0062; B = 16'h006C; #100;
A = 16'h0062; B = 16'h006D; #100;
A = 16'h0062; B = 16'h006E; #100;
A = 16'h0062; B = 16'h006F; #100;
A = 16'h0062; B = 16'h0070; #100;
A = 16'h0062; B = 16'h0071; #100;
A = 16'h0062; B = 16'h0072; #100;
A = 16'h0062; B = 16'h0073; #100;
A = 16'h0062; B = 16'h0074; #100;
A = 16'h0062; B = 16'h0075; #100;
A = 16'h0062; B = 16'h0076; #100;
A = 16'h0062; B = 16'h0077; #100;
A = 16'h0062; B = 16'h0078; #100;
A = 16'h0062; B = 16'h0079; #100;
A = 16'h0062; B = 16'h007A; #100;
A = 16'h0062; B = 16'h007B; #100;
A = 16'h0062; B = 16'h007C; #100;
A = 16'h0062; B = 16'h007D; #100;
A = 16'h0062; B = 16'h007E; #100;
A = 16'h0062; B = 16'h007F; #100;
A = 16'h0062; B = 16'h0080; #100;
A = 16'h0062; B = 16'h0081; #100;
A = 16'h0062; B = 16'h0082; #100;
A = 16'h0062; B = 16'h0083; #100;
A = 16'h0062; B = 16'h0084; #100;
A = 16'h0062; B = 16'h0085; #100;
A = 16'h0062; B = 16'h0086; #100;
A = 16'h0062; B = 16'h0087; #100;
A = 16'h0062; B = 16'h0088; #100;
A = 16'h0062; B = 16'h0089; #100;
A = 16'h0062; B = 16'h008A; #100;
A = 16'h0062; B = 16'h008B; #100;
A = 16'h0062; B = 16'h008C; #100;
A = 16'h0062; B = 16'h008D; #100;
A = 16'h0062; B = 16'h008E; #100;
A = 16'h0062; B = 16'h008F; #100;
A = 16'h0062; B = 16'h0090; #100;
A = 16'h0062; B = 16'h0091; #100;
A = 16'h0062; B = 16'h0092; #100;
A = 16'h0062; B = 16'h0093; #100;
A = 16'h0062; B = 16'h0094; #100;
A = 16'h0062; B = 16'h0095; #100;
A = 16'h0062; B = 16'h0096; #100;
A = 16'h0062; B = 16'h0097; #100;
A = 16'h0062; B = 16'h0098; #100;
A = 16'h0062; B = 16'h0099; #100;
A = 16'h0062; B = 16'h009A; #100;
A = 16'h0062; B = 16'h009B; #100;
A = 16'h0062; B = 16'h009C; #100;
A = 16'h0062; B = 16'h009D; #100;
A = 16'h0062; B = 16'h009E; #100;
A = 16'h0062; B = 16'h009F; #100;
A = 16'h0062; B = 16'h00A0; #100;
A = 16'h0062; B = 16'h00A1; #100;
A = 16'h0062; B = 16'h00A2; #100;
A = 16'h0062; B = 16'h00A3; #100;
A = 16'h0062; B = 16'h00A4; #100;
A = 16'h0062; B = 16'h00A5; #100;
A = 16'h0062; B = 16'h00A6; #100;
A = 16'h0062; B = 16'h00A7; #100;
A = 16'h0062; B = 16'h00A8; #100;
A = 16'h0062; B = 16'h00A9; #100;
A = 16'h0062; B = 16'h00AA; #100;
A = 16'h0062; B = 16'h00AB; #100;
A = 16'h0062; B = 16'h00AC; #100;
A = 16'h0062; B = 16'h00AD; #100;
A = 16'h0062; B = 16'h00AE; #100;
A = 16'h0062; B = 16'h00AF; #100;
A = 16'h0062; B = 16'h00B0; #100;
A = 16'h0062; B = 16'h00B1; #100;
A = 16'h0062; B = 16'h00B2; #100;
A = 16'h0062; B = 16'h00B3; #100;
A = 16'h0062; B = 16'h00B4; #100;
A = 16'h0062; B = 16'h00B5; #100;
A = 16'h0062; B = 16'h00B6; #100;
A = 16'h0062; B = 16'h00B7; #100;
A = 16'h0062; B = 16'h00B8; #100;
A = 16'h0062; B = 16'h00B9; #100;
A = 16'h0062; B = 16'h00BA; #100;
A = 16'h0062; B = 16'h00BB; #100;
A = 16'h0062; B = 16'h00BC; #100;
A = 16'h0062; B = 16'h00BD; #100;
A = 16'h0062; B = 16'h00BE; #100;
A = 16'h0062; B = 16'h00BF; #100;
A = 16'h0062; B = 16'h00C0; #100;
A = 16'h0062; B = 16'h00C1; #100;
A = 16'h0062; B = 16'h00C2; #100;
A = 16'h0062; B = 16'h00C3; #100;
A = 16'h0062; B = 16'h00C4; #100;
A = 16'h0062; B = 16'h00C5; #100;
A = 16'h0062; B = 16'h00C6; #100;
A = 16'h0062; B = 16'h00C7; #100;
A = 16'h0062; B = 16'h00C8; #100;
A = 16'h0062; B = 16'h00C9; #100;
A = 16'h0062; B = 16'h00CA; #100;
A = 16'h0062; B = 16'h00CB; #100;
A = 16'h0062; B = 16'h00CC; #100;
A = 16'h0062; B = 16'h00CD; #100;
A = 16'h0062; B = 16'h00CE; #100;
A = 16'h0062; B = 16'h00CF; #100;
A = 16'h0062; B = 16'h00D0; #100;
A = 16'h0062; B = 16'h00D1; #100;
A = 16'h0062; B = 16'h00D2; #100;
A = 16'h0062; B = 16'h00D3; #100;
A = 16'h0062; B = 16'h00D4; #100;
A = 16'h0062; B = 16'h00D5; #100;
A = 16'h0062; B = 16'h00D6; #100;
A = 16'h0062; B = 16'h00D7; #100;
A = 16'h0062; B = 16'h00D8; #100;
A = 16'h0062; B = 16'h00D9; #100;
A = 16'h0062; B = 16'h00DA; #100;
A = 16'h0062; B = 16'h00DB; #100;
A = 16'h0062; B = 16'h00DC; #100;
A = 16'h0062; B = 16'h00DD; #100;
A = 16'h0062; B = 16'h00DE; #100;
A = 16'h0062; B = 16'h00DF; #100;
A = 16'h0062; B = 16'h00E0; #100;
A = 16'h0062; B = 16'h00E1; #100;
A = 16'h0062; B = 16'h00E2; #100;
A = 16'h0062; B = 16'h00E3; #100;
A = 16'h0062; B = 16'h00E4; #100;
A = 16'h0062; B = 16'h00E5; #100;
A = 16'h0062; B = 16'h00E6; #100;
A = 16'h0062; B = 16'h00E7; #100;
A = 16'h0062; B = 16'h00E8; #100;
A = 16'h0062; B = 16'h00E9; #100;
A = 16'h0062; B = 16'h00EA; #100;
A = 16'h0062; B = 16'h00EB; #100;
A = 16'h0062; B = 16'h00EC; #100;
A = 16'h0062; B = 16'h00ED; #100;
A = 16'h0062; B = 16'h00EE; #100;
A = 16'h0062; B = 16'h00EF; #100;
A = 16'h0062; B = 16'h00F0; #100;
A = 16'h0062; B = 16'h00F1; #100;
A = 16'h0062; B = 16'h00F2; #100;
A = 16'h0062; B = 16'h00F3; #100;
A = 16'h0062; B = 16'h00F4; #100;
A = 16'h0062; B = 16'h00F5; #100;
A = 16'h0062; B = 16'h00F6; #100;
A = 16'h0062; B = 16'h00F7; #100;
A = 16'h0062; B = 16'h00F8; #100;
A = 16'h0062; B = 16'h00F9; #100;
A = 16'h0062; B = 16'h00FA; #100;
A = 16'h0062; B = 16'h00FB; #100;
A = 16'h0062; B = 16'h00FC; #100;
A = 16'h0062; B = 16'h00FD; #100;
A = 16'h0062; B = 16'h00FE; #100;
A = 16'h0062; B = 16'h00FF; #100;
A = 16'h0063; B = 16'h000; #100;
A = 16'h0063; B = 16'h001; #100;
A = 16'h0063; B = 16'h002; #100;
A = 16'h0063; B = 16'h003; #100;
A = 16'h0063; B = 16'h004; #100;
A = 16'h0063; B = 16'h005; #100;
A = 16'h0063; B = 16'h006; #100;
A = 16'h0063; B = 16'h007; #100;
A = 16'h0063; B = 16'h008; #100;
A = 16'h0063; B = 16'h009; #100;
A = 16'h0063; B = 16'h00A; #100;
A = 16'h0063; B = 16'h00B; #100;
A = 16'h0063; B = 16'h00C; #100;
A = 16'h0063; B = 16'h00D; #100;
A = 16'h0063; B = 16'h00E; #100;
A = 16'h0063; B = 16'h00F; #100;
A = 16'h0063; B = 16'h0010; #100;
A = 16'h0063; B = 16'h0011; #100;
A = 16'h0063; B = 16'h0012; #100;
A = 16'h0063; B = 16'h0013; #100;
A = 16'h0063; B = 16'h0014; #100;
A = 16'h0063; B = 16'h0015; #100;
A = 16'h0063; B = 16'h0016; #100;
A = 16'h0063; B = 16'h0017; #100;
A = 16'h0063; B = 16'h0018; #100;
A = 16'h0063; B = 16'h0019; #100;
A = 16'h0063; B = 16'h001A; #100;
A = 16'h0063; B = 16'h001B; #100;
A = 16'h0063; B = 16'h001C; #100;
A = 16'h0063; B = 16'h001D; #100;
A = 16'h0063; B = 16'h001E; #100;
A = 16'h0063; B = 16'h001F; #100;
A = 16'h0063; B = 16'h0020; #100;
A = 16'h0063; B = 16'h0021; #100;
A = 16'h0063; B = 16'h0022; #100;
A = 16'h0063; B = 16'h0023; #100;
A = 16'h0063; B = 16'h0024; #100;
A = 16'h0063; B = 16'h0025; #100;
A = 16'h0063; B = 16'h0026; #100;
A = 16'h0063; B = 16'h0027; #100;
A = 16'h0063; B = 16'h0028; #100;
A = 16'h0063; B = 16'h0029; #100;
A = 16'h0063; B = 16'h002A; #100;
A = 16'h0063; B = 16'h002B; #100;
A = 16'h0063; B = 16'h002C; #100;
A = 16'h0063; B = 16'h002D; #100;
A = 16'h0063; B = 16'h002E; #100;
A = 16'h0063; B = 16'h002F; #100;
A = 16'h0063; B = 16'h0030; #100;
A = 16'h0063; B = 16'h0031; #100;
A = 16'h0063; B = 16'h0032; #100;
A = 16'h0063; B = 16'h0033; #100;
A = 16'h0063; B = 16'h0034; #100;
A = 16'h0063; B = 16'h0035; #100;
A = 16'h0063; B = 16'h0036; #100;
A = 16'h0063; B = 16'h0037; #100;
A = 16'h0063; B = 16'h0038; #100;
A = 16'h0063; B = 16'h0039; #100;
A = 16'h0063; B = 16'h003A; #100;
A = 16'h0063; B = 16'h003B; #100;
A = 16'h0063; B = 16'h003C; #100;
A = 16'h0063; B = 16'h003D; #100;
A = 16'h0063; B = 16'h003E; #100;
A = 16'h0063; B = 16'h003F; #100;
A = 16'h0063; B = 16'h0040; #100;
A = 16'h0063; B = 16'h0041; #100;
A = 16'h0063; B = 16'h0042; #100;
A = 16'h0063; B = 16'h0043; #100;
A = 16'h0063; B = 16'h0044; #100;
A = 16'h0063; B = 16'h0045; #100;
A = 16'h0063; B = 16'h0046; #100;
A = 16'h0063; B = 16'h0047; #100;
A = 16'h0063; B = 16'h0048; #100;
A = 16'h0063; B = 16'h0049; #100;
A = 16'h0063; B = 16'h004A; #100;
A = 16'h0063; B = 16'h004B; #100;
A = 16'h0063; B = 16'h004C; #100;
A = 16'h0063; B = 16'h004D; #100;
A = 16'h0063; B = 16'h004E; #100;
A = 16'h0063; B = 16'h004F; #100;
A = 16'h0063; B = 16'h0050; #100;
A = 16'h0063; B = 16'h0051; #100;
A = 16'h0063; B = 16'h0052; #100;
A = 16'h0063; B = 16'h0053; #100;
A = 16'h0063; B = 16'h0054; #100;
A = 16'h0063; B = 16'h0055; #100;
A = 16'h0063; B = 16'h0056; #100;
A = 16'h0063; B = 16'h0057; #100;
A = 16'h0063; B = 16'h0058; #100;
A = 16'h0063; B = 16'h0059; #100;
A = 16'h0063; B = 16'h005A; #100;
A = 16'h0063; B = 16'h005B; #100;
A = 16'h0063; B = 16'h005C; #100;
A = 16'h0063; B = 16'h005D; #100;
A = 16'h0063; B = 16'h005E; #100;
A = 16'h0063; B = 16'h005F; #100;
A = 16'h0063; B = 16'h0060; #100;
A = 16'h0063; B = 16'h0061; #100;
A = 16'h0063; B = 16'h0062; #100;
A = 16'h0063; B = 16'h0063; #100;
A = 16'h0063; B = 16'h0064; #100;
A = 16'h0063; B = 16'h0065; #100;
A = 16'h0063; B = 16'h0066; #100;
A = 16'h0063; B = 16'h0067; #100;
A = 16'h0063; B = 16'h0068; #100;
A = 16'h0063; B = 16'h0069; #100;
A = 16'h0063; B = 16'h006A; #100;
A = 16'h0063; B = 16'h006B; #100;
A = 16'h0063; B = 16'h006C; #100;
A = 16'h0063; B = 16'h006D; #100;
A = 16'h0063; B = 16'h006E; #100;
A = 16'h0063; B = 16'h006F; #100;
A = 16'h0063; B = 16'h0070; #100;
A = 16'h0063; B = 16'h0071; #100;
A = 16'h0063; B = 16'h0072; #100;
A = 16'h0063; B = 16'h0073; #100;
A = 16'h0063; B = 16'h0074; #100;
A = 16'h0063; B = 16'h0075; #100;
A = 16'h0063; B = 16'h0076; #100;
A = 16'h0063; B = 16'h0077; #100;
A = 16'h0063; B = 16'h0078; #100;
A = 16'h0063; B = 16'h0079; #100;
A = 16'h0063; B = 16'h007A; #100;
A = 16'h0063; B = 16'h007B; #100;
A = 16'h0063; B = 16'h007C; #100;
A = 16'h0063; B = 16'h007D; #100;
A = 16'h0063; B = 16'h007E; #100;
A = 16'h0063; B = 16'h007F; #100;
A = 16'h0063; B = 16'h0080; #100;
A = 16'h0063; B = 16'h0081; #100;
A = 16'h0063; B = 16'h0082; #100;
A = 16'h0063; B = 16'h0083; #100;
A = 16'h0063; B = 16'h0084; #100;
A = 16'h0063; B = 16'h0085; #100;
A = 16'h0063; B = 16'h0086; #100;
A = 16'h0063; B = 16'h0087; #100;
A = 16'h0063; B = 16'h0088; #100;
A = 16'h0063; B = 16'h0089; #100;
A = 16'h0063; B = 16'h008A; #100;
A = 16'h0063; B = 16'h008B; #100;
A = 16'h0063; B = 16'h008C; #100;
A = 16'h0063; B = 16'h008D; #100;
A = 16'h0063; B = 16'h008E; #100;
A = 16'h0063; B = 16'h008F; #100;
A = 16'h0063; B = 16'h0090; #100;
A = 16'h0063; B = 16'h0091; #100;
A = 16'h0063; B = 16'h0092; #100;
A = 16'h0063; B = 16'h0093; #100;
A = 16'h0063; B = 16'h0094; #100;
A = 16'h0063; B = 16'h0095; #100;
A = 16'h0063; B = 16'h0096; #100;
A = 16'h0063; B = 16'h0097; #100;
A = 16'h0063; B = 16'h0098; #100;
A = 16'h0063; B = 16'h0099; #100;
A = 16'h0063; B = 16'h009A; #100;
A = 16'h0063; B = 16'h009B; #100;
A = 16'h0063; B = 16'h009C; #100;
A = 16'h0063; B = 16'h009D; #100;
A = 16'h0063; B = 16'h009E; #100;
A = 16'h0063; B = 16'h009F; #100;
A = 16'h0063; B = 16'h00A0; #100;
A = 16'h0063; B = 16'h00A1; #100;
A = 16'h0063; B = 16'h00A2; #100;
A = 16'h0063; B = 16'h00A3; #100;
A = 16'h0063; B = 16'h00A4; #100;
A = 16'h0063; B = 16'h00A5; #100;
A = 16'h0063; B = 16'h00A6; #100;
A = 16'h0063; B = 16'h00A7; #100;
A = 16'h0063; B = 16'h00A8; #100;
A = 16'h0063; B = 16'h00A9; #100;
A = 16'h0063; B = 16'h00AA; #100;
A = 16'h0063; B = 16'h00AB; #100;
A = 16'h0063; B = 16'h00AC; #100;
A = 16'h0063; B = 16'h00AD; #100;
A = 16'h0063; B = 16'h00AE; #100;
A = 16'h0063; B = 16'h00AF; #100;
A = 16'h0063; B = 16'h00B0; #100;
A = 16'h0063; B = 16'h00B1; #100;
A = 16'h0063; B = 16'h00B2; #100;
A = 16'h0063; B = 16'h00B3; #100;
A = 16'h0063; B = 16'h00B4; #100;
A = 16'h0063; B = 16'h00B5; #100;
A = 16'h0063; B = 16'h00B6; #100;
A = 16'h0063; B = 16'h00B7; #100;
A = 16'h0063; B = 16'h00B8; #100;
A = 16'h0063; B = 16'h00B9; #100;
A = 16'h0063; B = 16'h00BA; #100;
A = 16'h0063; B = 16'h00BB; #100;
A = 16'h0063; B = 16'h00BC; #100;
A = 16'h0063; B = 16'h00BD; #100;
A = 16'h0063; B = 16'h00BE; #100;
A = 16'h0063; B = 16'h00BF; #100;
A = 16'h0063; B = 16'h00C0; #100;
A = 16'h0063; B = 16'h00C1; #100;
A = 16'h0063; B = 16'h00C2; #100;
A = 16'h0063; B = 16'h00C3; #100;
A = 16'h0063; B = 16'h00C4; #100;
A = 16'h0063; B = 16'h00C5; #100;
A = 16'h0063; B = 16'h00C6; #100;
A = 16'h0063; B = 16'h00C7; #100;
A = 16'h0063; B = 16'h00C8; #100;
A = 16'h0063; B = 16'h00C9; #100;
A = 16'h0063; B = 16'h00CA; #100;
A = 16'h0063; B = 16'h00CB; #100;
A = 16'h0063; B = 16'h00CC; #100;
A = 16'h0063; B = 16'h00CD; #100;
A = 16'h0063; B = 16'h00CE; #100;
A = 16'h0063; B = 16'h00CF; #100;
A = 16'h0063; B = 16'h00D0; #100;
A = 16'h0063; B = 16'h00D1; #100;
A = 16'h0063; B = 16'h00D2; #100;
A = 16'h0063; B = 16'h00D3; #100;
A = 16'h0063; B = 16'h00D4; #100;
A = 16'h0063; B = 16'h00D5; #100;
A = 16'h0063; B = 16'h00D6; #100;
A = 16'h0063; B = 16'h00D7; #100;
A = 16'h0063; B = 16'h00D8; #100;
A = 16'h0063; B = 16'h00D9; #100;
A = 16'h0063; B = 16'h00DA; #100;
A = 16'h0063; B = 16'h00DB; #100;
A = 16'h0063; B = 16'h00DC; #100;
A = 16'h0063; B = 16'h00DD; #100;
A = 16'h0063; B = 16'h00DE; #100;
A = 16'h0063; B = 16'h00DF; #100;
A = 16'h0063; B = 16'h00E0; #100;
A = 16'h0063; B = 16'h00E1; #100;
A = 16'h0063; B = 16'h00E2; #100;
A = 16'h0063; B = 16'h00E3; #100;
A = 16'h0063; B = 16'h00E4; #100;
A = 16'h0063; B = 16'h00E5; #100;
A = 16'h0063; B = 16'h00E6; #100;
A = 16'h0063; B = 16'h00E7; #100;
A = 16'h0063; B = 16'h00E8; #100;
A = 16'h0063; B = 16'h00E9; #100;
A = 16'h0063; B = 16'h00EA; #100;
A = 16'h0063; B = 16'h00EB; #100;
A = 16'h0063; B = 16'h00EC; #100;
A = 16'h0063; B = 16'h00ED; #100;
A = 16'h0063; B = 16'h00EE; #100;
A = 16'h0063; B = 16'h00EF; #100;
A = 16'h0063; B = 16'h00F0; #100;
A = 16'h0063; B = 16'h00F1; #100;
A = 16'h0063; B = 16'h00F2; #100;
A = 16'h0063; B = 16'h00F3; #100;
A = 16'h0063; B = 16'h00F4; #100;
A = 16'h0063; B = 16'h00F5; #100;
A = 16'h0063; B = 16'h00F6; #100;
A = 16'h0063; B = 16'h00F7; #100;
A = 16'h0063; B = 16'h00F8; #100;
A = 16'h0063; B = 16'h00F9; #100;
A = 16'h0063; B = 16'h00FA; #100;
A = 16'h0063; B = 16'h00FB; #100;
A = 16'h0063; B = 16'h00FC; #100;
A = 16'h0063; B = 16'h00FD; #100;
A = 16'h0063; B = 16'h00FE; #100;
A = 16'h0063; B = 16'h00FF; #100;
A = 16'h0064; B = 16'h000; #100;
A = 16'h0064; B = 16'h001; #100;
A = 16'h0064; B = 16'h002; #100;
A = 16'h0064; B = 16'h003; #100;
A = 16'h0064; B = 16'h004; #100;
A = 16'h0064; B = 16'h005; #100;
A = 16'h0064; B = 16'h006; #100;
A = 16'h0064; B = 16'h007; #100;
A = 16'h0064; B = 16'h008; #100;
A = 16'h0064; B = 16'h009; #100;
A = 16'h0064; B = 16'h00A; #100;
A = 16'h0064; B = 16'h00B; #100;
A = 16'h0064; B = 16'h00C; #100;
A = 16'h0064; B = 16'h00D; #100;
A = 16'h0064; B = 16'h00E; #100;
A = 16'h0064; B = 16'h00F; #100;
A = 16'h0064; B = 16'h0010; #100;
A = 16'h0064; B = 16'h0011; #100;
A = 16'h0064; B = 16'h0012; #100;
A = 16'h0064; B = 16'h0013; #100;
A = 16'h0064; B = 16'h0014; #100;
A = 16'h0064; B = 16'h0015; #100;
A = 16'h0064; B = 16'h0016; #100;
A = 16'h0064; B = 16'h0017; #100;
A = 16'h0064; B = 16'h0018; #100;
A = 16'h0064; B = 16'h0019; #100;
A = 16'h0064; B = 16'h001A; #100;
A = 16'h0064; B = 16'h001B; #100;
A = 16'h0064; B = 16'h001C; #100;
A = 16'h0064; B = 16'h001D; #100;
A = 16'h0064; B = 16'h001E; #100;
A = 16'h0064; B = 16'h001F; #100;
A = 16'h0064; B = 16'h0020; #100;
A = 16'h0064; B = 16'h0021; #100;
A = 16'h0064; B = 16'h0022; #100;
A = 16'h0064; B = 16'h0023; #100;
A = 16'h0064; B = 16'h0024; #100;
A = 16'h0064; B = 16'h0025; #100;
A = 16'h0064; B = 16'h0026; #100;
A = 16'h0064; B = 16'h0027; #100;
A = 16'h0064; B = 16'h0028; #100;
A = 16'h0064; B = 16'h0029; #100;
A = 16'h0064; B = 16'h002A; #100;
A = 16'h0064; B = 16'h002B; #100;
A = 16'h0064; B = 16'h002C; #100;
A = 16'h0064; B = 16'h002D; #100;
A = 16'h0064; B = 16'h002E; #100;
A = 16'h0064; B = 16'h002F; #100;
A = 16'h0064; B = 16'h0030; #100;
A = 16'h0064; B = 16'h0031; #100;
A = 16'h0064; B = 16'h0032; #100;
A = 16'h0064; B = 16'h0033; #100;
A = 16'h0064; B = 16'h0034; #100;
A = 16'h0064; B = 16'h0035; #100;
A = 16'h0064; B = 16'h0036; #100;
A = 16'h0064; B = 16'h0037; #100;
A = 16'h0064; B = 16'h0038; #100;
A = 16'h0064; B = 16'h0039; #100;
A = 16'h0064; B = 16'h003A; #100;
A = 16'h0064; B = 16'h003B; #100;
A = 16'h0064; B = 16'h003C; #100;
A = 16'h0064; B = 16'h003D; #100;
A = 16'h0064; B = 16'h003E; #100;
A = 16'h0064; B = 16'h003F; #100;
A = 16'h0064; B = 16'h0040; #100;
A = 16'h0064; B = 16'h0041; #100;
A = 16'h0064; B = 16'h0042; #100;
A = 16'h0064; B = 16'h0043; #100;
A = 16'h0064; B = 16'h0044; #100;
A = 16'h0064; B = 16'h0045; #100;
A = 16'h0064; B = 16'h0046; #100;
A = 16'h0064; B = 16'h0047; #100;
A = 16'h0064; B = 16'h0048; #100;
A = 16'h0064; B = 16'h0049; #100;
A = 16'h0064; B = 16'h004A; #100;
A = 16'h0064; B = 16'h004B; #100;
A = 16'h0064; B = 16'h004C; #100;
A = 16'h0064; B = 16'h004D; #100;
A = 16'h0064; B = 16'h004E; #100;
A = 16'h0064; B = 16'h004F; #100;
A = 16'h0064; B = 16'h0050; #100;
A = 16'h0064; B = 16'h0051; #100;
A = 16'h0064; B = 16'h0052; #100;
A = 16'h0064; B = 16'h0053; #100;
A = 16'h0064; B = 16'h0054; #100;
A = 16'h0064; B = 16'h0055; #100;
A = 16'h0064; B = 16'h0056; #100;
A = 16'h0064; B = 16'h0057; #100;
A = 16'h0064; B = 16'h0058; #100;
A = 16'h0064; B = 16'h0059; #100;
A = 16'h0064; B = 16'h005A; #100;
A = 16'h0064; B = 16'h005B; #100;
A = 16'h0064; B = 16'h005C; #100;
A = 16'h0064; B = 16'h005D; #100;
A = 16'h0064; B = 16'h005E; #100;
A = 16'h0064; B = 16'h005F; #100;
A = 16'h0064; B = 16'h0060; #100;
A = 16'h0064; B = 16'h0061; #100;
A = 16'h0064; B = 16'h0062; #100;
A = 16'h0064; B = 16'h0063; #100;
A = 16'h0064; B = 16'h0064; #100;
A = 16'h0064; B = 16'h0065; #100;
A = 16'h0064; B = 16'h0066; #100;
A = 16'h0064; B = 16'h0067; #100;
A = 16'h0064; B = 16'h0068; #100;
A = 16'h0064; B = 16'h0069; #100;
A = 16'h0064; B = 16'h006A; #100;
A = 16'h0064; B = 16'h006B; #100;
A = 16'h0064; B = 16'h006C; #100;
A = 16'h0064; B = 16'h006D; #100;
A = 16'h0064; B = 16'h006E; #100;
A = 16'h0064; B = 16'h006F; #100;
A = 16'h0064; B = 16'h0070; #100;
A = 16'h0064; B = 16'h0071; #100;
A = 16'h0064; B = 16'h0072; #100;
A = 16'h0064; B = 16'h0073; #100;
A = 16'h0064; B = 16'h0074; #100;
A = 16'h0064; B = 16'h0075; #100;
A = 16'h0064; B = 16'h0076; #100;
A = 16'h0064; B = 16'h0077; #100;
A = 16'h0064; B = 16'h0078; #100;
A = 16'h0064; B = 16'h0079; #100;
A = 16'h0064; B = 16'h007A; #100;
A = 16'h0064; B = 16'h007B; #100;
A = 16'h0064; B = 16'h007C; #100;
A = 16'h0064; B = 16'h007D; #100;
A = 16'h0064; B = 16'h007E; #100;
A = 16'h0064; B = 16'h007F; #100;
A = 16'h0064; B = 16'h0080; #100;
A = 16'h0064; B = 16'h0081; #100;
A = 16'h0064; B = 16'h0082; #100;
A = 16'h0064; B = 16'h0083; #100;
A = 16'h0064; B = 16'h0084; #100;
A = 16'h0064; B = 16'h0085; #100;
A = 16'h0064; B = 16'h0086; #100;
A = 16'h0064; B = 16'h0087; #100;
A = 16'h0064; B = 16'h0088; #100;
A = 16'h0064; B = 16'h0089; #100;
A = 16'h0064; B = 16'h008A; #100;
A = 16'h0064; B = 16'h008B; #100;
A = 16'h0064; B = 16'h008C; #100;
A = 16'h0064; B = 16'h008D; #100;
A = 16'h0064; B = 16'h008E; #100;
A = 16'h0064; B = 16'h008F; #100;
A = 16'h0064; B = 16'h0090; #100;
A = 16'h0064; B = 16'h0091; #100;
A = 16'h0064; B = 16'h0092; #100;
A = 16'h0064; B = 16'h0093; #100;
A = 16'h0064; B = 16'h0094; #100;
A = 16'h0064; B = 16'h0095; #100;
A = 16'h0064; B = 16'h0096; #100;
A = 16'h0064; B = 16'h0097; #100;
A = 16'h0064; B = 16'h0098; #100;
A = 16'h0064; B = 16'h0099; #100;
A = 16'h0064; B = 16'h009A; #100;
A = 16'h0064; B = 16'h009B; #100;
A = 16'h0064; B = 16'h009C; #100;
A = 16'h0064; B = 16'h009D; #100;
A = 16'h0064; B = 16'h009E; #100;
A = 16'h0064; B = 16'h009F; #100;
A = 16'h0064; B = 16'h00A0; #100;
A = 16'h0064; B = 16'h00A1; #100;
A = 16'h0064; B = 16'h00A2; #100;
A = 16'h0064; B = 16'h00A3; #100;
A = 16'h0064; B = 16'h00A4; #100;
A = 16'h0064; B = 16'h00A5; #100;
A = 16'h0064; B = 16'h00A6; #100;
A = 16'h0064; B = 16'h00A7; #100;
A = 16'h0064; B = 16'h00A8; #100;
A = 16'h0064; B = 16'h00A9; #100;
A = 16'h0064; B = 16'h00AA; #100;
A = 16'h0064; B = 16'h00AB; #100;
A = 16'h0064; B = 16'h00AC; #100;
A = 16'h0064; B = 16'h00AD; #100;
A = 16'h0064; B = 16'h00AE; #100;
A = 16'h0064; B = 16'h00AF; #100;
A = 16'h0064; B = 16'h00B0; #100;
A = 16'h0064; B = 16'h00B1; #100;
A = 16'h0064; B = 16'h00B2; #100;
A = 16'h0064; B = 16'h00B3; #100;
A = 16'h0064; B = 16'h00B4; #100;
A = 16'h0064; B = 16'h00B5; #100;
A = 16'h0064; B = 16'h00B6; #100;
A = 16'h0064; B = 16'h00B7; #100;
A = 16'h0064; B = 16'h00B8; #100;
A = 16'h0064; B = 16'h00B9; #100;
A = 16'h0064; B = 16'h00BA; #100;
A = 16'h0064; B = 16'h00BB; #100;
A = 16'h0064; B = 16'h00BC; #100;
A = 16'h0064; B = 16'h00BD; #100;
A = 16'h0064; B = 16'h00BE; #100;
A = 16'h0064; B = 16'h00BF; #100;
A = 16'h0064; B = 16'h00C0; #100;
A = 16'h0064; B = 16'h00C1; #100;
A = 16'h0064; B = 16'h00C2; #100;
A = 16'h0064; B = 16'h00C3; #100;
A = 16'h0064; B = 16'h00C4; #100;
A = 16'h0064; B = 16'h00C5; #100;
A = 16'h0064; B = 16'h00C6; #100;
A = 16'h0064; B = 16'h00C7; #100;
A = 16'h0064; B = 16'h00C8; #100;
A = 16'h0064; B = 16'h00C9; #100;
A = 16'h0064; B = 16'h00CA; #100;
A = 16'h0064; B = 16'h00CB; #100;
A = 16'h0064; B = 16'h00CC; #100;
A = 16'h0064; B = 16'h00CD; #100;
A = 16'h0064; B = 16'h00CE; #100;
A = 16'h0064; B = 16'h00CF; #100;
A = 16'h0064; B = 16'h00D0; #100;
A = 16'h0064; B = 16'h00D1; #100;
A = 16'h0064; B = 16'h00D2; #100;
A = 16'h0064; B = 16'h00D3; #100;
A = 16'h0064; B = 16'h00D4; #100;
A = 16'h0064; B = 16'h00D5; #100;
A = 16'h0064; B = 16'h00D6; #100;
A = 16'h0064; B = 16'h00D7; #100;
A = 16'h0064; B = 16'h00D8; #100;
A = 16'h0064; B = 16'h00D9; #100;
A = 16'h0064; B = 16'h00DA; #100;
A = 16'h0064; B = 16'h00DB; #100;
A = 16'h0064; B = 16'h00DC; #100;
A = 16'h0064; B = 16'h00DD; #100;
A = 16'h0064; B = 16'h00DE; #100;
A = 16'h0064; B = 16'h00DF; #100;
A = 16'h0064; B = 16'h00E0; #100;
A = 16'h0064; B = 16'h00E1; #100;
A = 16'h0064; B = 16'h00E2; #100;
A = 16'h0064; B = 16'h00E3; #100;
A = 16'h0064; B = 16'h00E4; #100;
A = 16'h0064; B = 16'h00E5; #100;
A = 16'h0064; B = 16'h00E6; #100;
A = 16'h0064; B = 16'h00E7; #100;
A = 16'h0064; B = 16'h00E8; #100;
A = 16'h0064; B = 16'h00E9; #100;
A = 16'h0064; B = 16'h00EA; #100;
A = 16'h0064; B = 16'h00EB; #100;
A = 16'h0064; B = 16'h00EC; #100;
A = 16'h0064; B = 16'h00ED; #100;
A = 16'h0064; B = 16'h00EE; #100;
A = 16'h0064; B = 16'h00EF; #100;
A = 16'h0064; B = 16'h00F0; #100;
A = 16'h0064; B = 16'h00F1; #100;
A = 16'h0064; B = 16'h00F2; #100;
A = 16'h0064; B = 16'h00F3; #100;
A = 16'h0064; B = 16'h00F4; #100;
A = 16'h0064; B = 16'h00F5; #100;
A = 16'h0064; B = 16'h00F6; #100;
A = 16'h0064; B = 16'h00F7; #100;
A = 16'h0064; B = 16'h00F8; #100;
A = 16'h0064; B = 16'h00F9; #100;
A = 16'h0064; B = 16'h00FA; #100;
A = 16'h0064; B = 16'h00FB; #100;
A = 16'h0064; B = 16'h00FC; #100;
A = 16'h0064; B = 16'h00FD; #100;
A = 16'h0064; B = 16'h00FE; #100;
A = 16'h0064; B = 16'h00FF; #100;
A = 16'h0065; B = 16'h000; #100;
A = 16'h0065; B = 16'h001; #100;
A = 16'h0065; B = 16'h002; #100;
A = 16'h0065; B = 16'h003; #100;
A = 16'h0065; B = 16'h004; #100;
A = 16'h0065; B = 16'h005; #100;
A = 16'h0065; B = 16'h006; #100;
A = 16'h0065; B = 16'h007; #100;
A = 16'h0065; B = 16'h008; #100;
A = 16'h0065; B = 16'h009; #100;
A = 16'h0065; B = 16'h00A; #100;
A = 16'h0065; B = 16'h00B; #100;
A = 16'h0065; B = 16'h00C; #100;
A = 16'h0065; B = 16'h00D; #100;
A = 16'h0065; B = 16'h00E; #100;
A = 16'h0065; B = 16'h00F; #100;
A = 16'h0065; B = 16'h0010; #100;
A = 16'h0065; B = 16'h0011; #100;
A = 16'h0065; B = 16'h0012; #100;
A = 16'h0065; B = 16'h0013; #100;
A = 16'h0065; B = 16'h0014; #100;
A = 16'h0065; B = 16'h0015; #100;
A = 16'h0065; B = 16'h0016; #100;
A = 16'h0065; B = 16'h0017; #100;
A = 16'h0065; B = 16'h0018; #100;
A = 16'h0065; B = 16'h0019; #100;
A = 16'h0065; B = 16'h001A; #100;
A = 16'h0065; B = 16'h001B; #100;
A = 16'h0065; B = 16'h001C; #100;
A = 16'h0065; B = 16'h001D; #100;
A = 16'h0065; B = 16'h001E; #100;
A = 16'h0065; B = 16'h001F; #100;
A = 16'h0065; B = 16'h0020; #100;
A = 16'h0065; B = 16'h0021; #100;
A = 16'h0065; B = 16'h0022; #100;
A = 16'h0065; B = 16'h0023; #100;
A = 16'h0065; B = 16'h0024; #100;
A = 16'h0065; B = 16'h0025; #100;
A = 16'h0065; B = 16'h0026; #100;
A = 16'h0065; B = 16'h0027; #100;
A = 16'h0065; B = 16'h0028; #100;
A = 16'h0065; B = 16'h0029; #100;
A = 16'h0065; B = 16'h002A; #100;
A = 16'h0065; B = 16'h002B; #100;
A = 16'h0065; B = 16'h002C; #100;
A = 16'h0065; B = 16'h002D; #100;
A = 16'h0065; B = 16'h002E; #100;
A = 16'h0065; B = 16'h002F; #100;
A = 16'h0065; B = 16'h0030; #100;
A = 16'h0065; B = 16'h0031; #100;
A = 16'h0065; B = 16'h0032; #100;
A = 16'h0065; B = 16'h0033; #100;
A = 16'h0065; B = 16'h0034; #100;
A = 16'h0065; B = 16'h0035; #100;
A = 16'h0065; B = 16'h0036; #100;
A = 16'h0065; B = 16'h0037; #100;
A = 16'h0065; B = 16'h0038; #100;
A = 16'h0065; B = 16'h0039; #100;
A = 16'h0065; B = 16'h003A; #100;
A = 16'h0065; B = 16'h003B; #100;
A = 16'h0065; B = 16'h003C; #100;
A = 16'h0065; B = 16'h003D; #100;
A = 16'h0065; B = 16'h003E; #100;
A = 16'h0065; B = 16'h003F; #100;
A = 16'h0065; B = 16'h0040; #100;
A = 16'h0065; B = 16'h0041; #100;
A = 16'h0065; B = 16'h0042; #100;
A = 16'h0065; B = 16'h0043; #100;
A = 16'h0065; B = 16'h0044; #100;
A = 16'h0065; B = 16'h0045; #100;
A = 16'h0065; B = 16'h0046; #100;
A = 16'h0065; B = 16'h0047; #100;
A = 16'h0065; B = 16'h0048; #100;
A = 16'h0065; B = 16'h0049; #100;
A = 16'h0065; B = 16'h004A; #100;
A = 16'h0065; B = 16'h004B; #100;
A = 16'h0065; B = 16'h004C; #100;
A = 16'h0065; B = 16'h004D; #100;
A = 16'h0065; B = 16'h004E; #100;
A = 16'h0065; B = 16'h004F; #100;
A = 16'h0065; B = 16'h0050; #100;
A = 16'h0065; B = 16'h0051; #100;
A = 16'h0065; B = 16'h0052; #100;
A = 16'h0065; B = 16'h0053; #100;
A = 16'h0065; B = 16'h0054; #100;
A = 16'h0065; B = 16'h0055; #100;
A = 16'h0065; B = 16'h0056; #100;
A = 16'h0065; B = 16'h0057; #100;
A = 16'h0065; B = 16'h0058; #100;
A = 16'h0065; B = 16'h0059; #100;
A = 16'h0065; B = 16'h005A; #100;
A = 16'h0065; B = 16'h005B; #100;
A = 16'h0065; B = 16'h005C; #100;
A = 16'h0065; B = 16'h005D; #100;
A = 16'h0065; B = 16'h005E; #100;
A = 16'h0065; B = 16'h005F; #100;
A = 16'h0065; B = 16'h0060; #100;
A = 16'h0065; B = 16'h0061; #100;
A = 16'h0065; B = 16'h0062; #100;
A = 16'h0065; B = 16'h0063; #100;
A = 16'h0065; B = 16'h0064; #100;
A = 16'h0065; B = 16'h0065; #100;
A = 16'h0065; B = 16'h0066; #100;
A = 16'h0065; B = 16'h0067; #100;
A = 16'h0065; B = 16'h0068; #100;
A = 16'h0065; B = 16'h0069; #100;
A = 16'h0065; B = 16'h006A; #100;
A = 16'h0065; B = 16'h006B; #100;
A = 16'h0065; B = 16'h006C; #100;
A = 16'h0065; B = 16'h006D; #100;
A = 16'h0065; B = 16'h006E; #100;
A = 16'h0065; B = 16'h006F; #100;
A = 16'h0065; B = 16'h0070; #100;
A = 16'h0065; B = 16'h0071; #100;
A = 16'h0065; B = 16'h0072; #100;
A = 16'h0065; B = 16'h0073; #100;
A = 16'h0065; B = 16'h0074; #100;
A = 16'h0065; B = 16'h0075; #100;
A = 16'h0065; B = 16'h0076; #100;
A = 16'h0065; B = 16'h0077; #100;
A = 16'h0065; B = 16'h0078; #100;
A = 16'h0065; B = 16'h0079; #100;
A = 16'h0065; B = 16'h007A; #100;
A = 16'h0065; B = 16'h007B; #100;
A = 16'h0065; B = 16'h007C; #100;
A = 16'h0065; B = 16'h007D; #100;
A = 16'h0065; B = 16'h007E; #100;
A = 16'h0065; B = 16'h007F; #100;
A = 16'h0065; B = 16'h0080; #100;
A = 16'h0065; B = 16'h0081; #100;
A = 16'h0065; B = 16'h0082; #100;
A = 16'h0065; B = 16'h0083; #100;
A = 16'h0065; B = 16'h0084; #100;
A = 16'h0065; B = 16'h0085; #100;
A = 16'h0065; B = 16'h0086; #100;
A = 16'h0065; B = 16'h0087; #100;
A = 16'h0065; B = 16'h0088; #100;
A = 16'h0065; B = 16'h0089; #100;
A = 16'h0065; B = 16'h008A; #100;
A = 16'h0065; B = 16'h008B; #100;
A = 16'h0065; B = 16'h008C; #100;
A = 16'h0065; B = 16'h008D; #100;
A = 16'h0065; B = 16'h008E; #100;
A = 16'h0065; B = 16'h008F; #100;
A = 16'h0065; B = 16'h0090; #100;
A = 16'h0065; B = 16'h0091; #100;
A = 16'h0065; B = 16'h0092; #100;
A = 16'h0065; B = 16'h0093; #100;
A = 16'h0065; B = 16'h0094; #100;
A = 16'h0065; B = 16'h0095; #100;
A = 16'h0065; B = 16'h0096; #100;
A = 16'h0065; B = 16'h0097; #100;
A = 16'h0065; B = 16'h0098; #100;
A = 16'h0065; B = 16'h0099; #100;
A = 16'h0065; B = 16'h009A; #100;
A = 16'h0065; B = 16'h009B; #100;
A = 16'h0065; B = 16'h009C; #100;
A = 16'h0065; B = 16'h009D; #100;
A = 16'h0065; B = 16'h009E; #100;
A = 16'h0065; B = 16'h009F; #100;
A = 16'h0065; B = 16'h00A0; #100;
A = 16'h0065; B = 16'h00A1; #100;
A = 16'h0065; B = 16'h00A2; #100;
A = 16'h0065; B = 16'h00A3; #100;
A = 16'h0065; B = 16'h00A4; #100;
A = 16'h0065; B = 16'h00A5; #100;
A = 16'h0065; B = 16'h00A6; #100;
A = 16'h0065; B = 16'h00A7; #100;
A = 16'h0065; B = 16'h00A8; #100;
A = 16'h0065; B = 16'h00A9; #100;
A = 16'h0065; B = 16'h00AA; #100;
A = 16'h0065; B = 16'h00AB; #100;
A = 16'h0065; B = 16'h00AC; #100;
A = 16'h0065; B = 16'h00AD; #100;
A = 16'h0065; B = 16'h00AE; #100;
A = 16'h0065; B = 16'h00AF; #100;
A = 16'h0065; B = 16'h00B0; #100;
A = 16'h0065; B = 16'h00B1; #100;
A = 16'h0065; B = 16'h00B2; #100;
A = 16'h0065; B = 16'h00B3; #100;
A = 16'h0065; B = 16'h00B4; #100;
A = 16'h0065; B = 16'h00B5; #100;
A = 16'h0065; B = 16'h00B6; #100;
A = 16'h0065; B = 16'h00B7; #100;
A = 16'h0065; B = 16'h00B8; #100;
A = 16'h0065; B = 16'h00B9; #100;
A = 16'h0065; B = 16'h00BA; #100;
A = 16'h0065; B = 16'h00BB; #100;
A = 16'h0065; B = 16'h00BC; #100;
A = 16'h0065; B = 16'h00BD; #100;
A = 16'h0065; B = 16'h00BE; #100;
A = 16'h0065; B = 16'h00BF; #100;
A = 16'h0065; B = 16'h00C0; #100;
A = 16'h0065; B = 16'h00C1; #100;
A = 16'h0065; B = 16'h00C2; #100;
A = 16'h0065; B = 16'h00C3; #100;
A = 16'h0065; B = 16'h00C4; #100;
A = 16'h0065; B = 16'h00C5; #100;
A = 16'h0065; B = 16'h00C6; #100;
A = 16'h0065; B = 16'h00C7; #100;
A = 16'h0065; B = 16'h00C8; #100;
A = 16'h0065; B = 16'h00C9; #100;
A = 16'h0065; B = 16'h00CA; #100;
A = 16'h0065; B = 16'h00CB; #100;
A = 16'h0065; B = 16'h00CC; #100;
A = 16'h0065; B = 16'h00CD; #100;
A = 16'h0065; B = 16'h00CE; #100;
A = 16'h0065; B = 16'h00CF; #100;
A = 16'h0065; B = 16'h00D0; #100;
A = 16'h0065; B = 16'h00D1; #100;
A = 16'h0065; B = 16'h00D2; #100;
A = 16'h0065; B = 16'h00D3; #100;
A = 16'h0065; B = 16'h00D4; #100;
A = 16'h0065; B = 16'h00D5; #100;
A = 16'h0065; B = 16'h00D6; #100;
A = 16'h0065; B = 16'h00D7; #100;
A = 16'h0065; B = 16'h00D8; #100;
A = 16'h0065; B = 16'h00D9; #100;
A = 16'h0065; B = 16'h00DA; #100;
A = 16'h0065; B = 16'h00DB; #100;
A = 16'h0065; B = 16'h00DC; #100;
A = 16'h0065; B = 16'h00DD; #100;
A = 16'h0065; B = 16'h00DE; #100;
A = 16'h0065; B = 16'h00DF; #100;
A = 16'h0065; B = 16'h00E0; #100;
A = 16'h0065; B = 16'h00E1; #100;
A = 16'h0065; B = 16'h00E2; #100;
A = 16'h0065; B = 16'h00E3; #100;
A = 16'h0065; B = 16'h00E4; #100;
A = 16'h0065; B = 16'h00E5; #100;
A = 16'h0065; B = 16'h00E6; #100;
A = 16'h0065; B = 16'h00E7; #100;
A = 16'h0065; B = 16'h00E8; #100;
A = 16'h0065; B = 16'h00E9; #100;
A = 16'h0065; B = 16'h00EA; #100;
A = 16'h0065; B = 16'h00EB; #100;
A = 16'h0065; B = 16'h00EC; #100;
A = 16'h0065; B = 16'h00ED; #100;
A = 16'h0065; B = 16'h00EE; #100;
A = 16'h0065; B = 16'h00EF; #100;
A = 16'h0065; B = 16'h00F0; #100;
A = 16'h0065; B = 16'h00F1; #100;
A = 16'h0065; B = 16'h00F2; #100;
A = 16'h0065; B = 16'h00F3; #100;
A = 16'h0065; B = 16'h00F4; #100;
A = 16'h0065; B = 16'h00F5; #100;
A = 16'h0065; B = 16'h00F6; #100;
A = 16'h0065; B = 16'h00F7; #100;
A = 16'h0065; B = 16'h00F8; #100;
A = 16'h0065; B = 16'h00F9; #100;
A = 16'h0065; B = 16'h00FA; #100;
A = 16'h0065; B = 16'h00FB; #100;
A = 16'h0065; B = 16'h00FC; #100;
A = 16'h0065; B = 16'h00FD; #100;
A = 16'h0065; B = 16'h00FE; #100;
A = 16'h0065; B = 16'h00FF; #100;
A = 16'h0066; B = 16'h000; #100;
A = 16'h0066; B = 16'h001; #100;
A = 16'h0066; B = 16'h002; #100;
A = 16'h0066; B = 16'h003; #100;
A = 16'h0066; B = 16'h004; #100;
A = 16'h0066; B = 16'h005; #100;
A = 16'h0066; B = 16'h006; #100;
A = 16'h0066; B = 16'h007; #100;
A = 16'h0066; B = 16'h008; #100;
A = 16'h0066; B = 16'h009; #100;
A = 16'h0066; B = 16'h00A; #100;
A = 16'h0066; B = 16'h00B; #100;
A = 16'h0066; B = 16'h00C; #100;
A = 16'h0066; B = 16'h00D; #100;
A = 16'h0066; B = 16'h00E; #100;
A = 16'h0066; B = 16'h00F; #100;
A = 16'h0066; B = 16'h0010; #100;
A = 16'h0066; B = 16'h0011; #100;
A = 16'h0066; B = 16'h0012; #100;
A = 16'h0066; B = 16'h0013; #100;
A = 16'h0066; B = 16'h0014; #100;
A = 16'h0066; B = 16'h0015; #100;
A = 16'h0066; B = 16'h0016; #100;
A = 16'h0066; B = 16'h0017; #100;
A = 16'h0066; B = 16'h0018; #100;
A = 16'h0066; B = 16'h0019; #100;
A = 16'h0066; B = 16'h001A; #100;
A = 16'h0066; B = 16'h001B; #100;
A = 16'h0066; B = 16'h001C; #100;
A = 16'h0066; B = 16'h001D; #100;
A = 16'h0066; B = 16'h001E; #100;
A = 16'h0066; B = 16'h001F; #100;
A = 16'h0066; B = 16'h0020; #100;
A = 16'h0066; B = 16'h0021; #100;
A = 16'h0066; B = 16'h0022; #100;
A = 16'h0066; B = 16'h0023; #100;
A = 16'h0066; B = 16'h0024; #100;
A = 16'h0066; B = 16'h0025; #100;
A = 16'h0066; B = 16'h0026; #100;
A = 16'h0066; B = 16'h0027; #100;
A = 16'h0066; B = 16'h0028; #100;
A = 16'h0066; B = 16'h0029; #100;
A = 16'h0066; B = 16'h002A; #100;
A = 16'h0066; B = 16'h002B; #100;
A = 16'h0066; B = 16'h002C; #100;
A = 16'h0066; B = 16'h002D; #100;
A = 16'h0066; B = 16'h002E; #100;
A = 16'h0066; B = 16'h002F; #100;
A = 16'h0066; B = 16'h0030; #100;
A = 16'h0066; B = 16'h0031; #100;
A = 16'h0066; B = 16'h0032; #100;
A = 16'h0066; B = 16'h0033; #100;
A = 16'h0066; B = 16'h0034; #100;
A = 16'h0066; B = 16'h0035; #100;
A = 16'h0066; B = 16'h0036; #100;
A = 16'h0066; B = 16'h0037; #100;
A = 16'h0066; B = 16'h0038; #100;
A = 16'h0066; B = 16'h0039; #100;
A = 16'h0066; B = 16'h003A; #100;
A = 16'h0066; B = 16'h003B; #100;
A = 16'h0066; B = 16'h003C; #100;
A = 16'h0066; B = 16'h003D; #100;
A = 16'h0066; B = 16'h003E; #100;
A = 16'h0066; B = 16'h003F; #100;
A = 16'h0066; B = 16'h0040; #100;
A = 16'h0066; B = 16'h0041; #100;
A = 16'h0066; B = 16'h0042; #100;
A = 16'h0066; B = 16'h0043; #100;
A = 16'h0066; B = 16'h0044; #100;
A = 16'h0066; B = 16'h0045; #100;
A = 16'h0066; B = 16'h0046; #100;
A = 16'h0066; B = 16'h0047; #100;
A = 16'h0066; B = 16'h0048; #100;
A = 16'h0066; B = 16'h0049; #100;
A = 16'h0066; B = 16'h004A; #100;
A = 16'h0066; B = 16'h004B; #100;
A = 16'h0066; B = 16'h004C; #100;
A = 16'h0066; B = 16'h004D; #100;
A = 16'h0066; B = 16'h004E; #100;
A = 16'h0066; B = 16'h004F; #100;
A = 16'h0066; B = 16'h0050; #100;
A = 16'h0066; B = 16'h0051; #100;
A = 16'h0066; B = 16'h0052; #100;
A = 16'h0066; B = 16'h0053; #100;
A = 16'h0066; B = 16'h0054; #100;
A = 16'h0066; B = 16'h0055; #100;
A = 16'h0066; B = 16'h0056; #100;
A = 16'h0066; B = 16'h0057; #100;
A = 16'h0066; B = 16'h0058; #100;
A = 16'h0066; B = 16'h0059; #100;
A = 16'h0066; B = 16'h005A; #100;
A = 16'h0066; B = 16'h005B; #100;
A = 16'h0066; B = 16'h005C; #100;
A = 16'h0066; B = 16'h005D; #100;
A = 16'h0066; B = 16'h005E; #100;
A = 16'h0066; B = 16'h005F; #100;
A = 16'h0066; B = 16'h0060; #100;
A = 16'h0066; B = 16'h0061; #100;
A = 16'h0066; B = 16'h0062; #100;
A = 16'h0066; B = 16'h0063; #100;
A = 16'h0066; B = 16'h0064; #100;
A = 16'h0066; B = 16'h0065; #100;
A = 16'h0066; B = 16'h0066; #100;
A = 16'h0066; B = 16'h0067; #100;
A = 16'h0066; B = 16'h0068; #100;
A = 16'h0066; B = 16'h0069; #100;
A = 16'h0066; B = 16'h006A; #100;
A = 16'h0066; B = 16'h006B; #100;
A = 16'h0066; B = 16'h006C; #100;
A = 16'h0066; B = 16'h006D; #100;
A = 16'h0066; B = 16'h006E; #100;
A = 16'h0066; B = 16'h006F; #100;
A = 16'h0066; B = 16'h0070; #100;
A = 16'h0066; B = 16'h0071; #100;
A = 16'h0066; B = 16'h0072; #100;
A = 16'h0066; B = 16'h0073; #100;
A = 16'h0066; B = 16'h0074; #100;
A = 16'h0066; B = 16'h0075; #100;
A = 16'h0066; B = 16'h0076; #100;
A = 16'h0066; B = 16'h0077; #100;
A = 16'h0066; B = 16'h0078; #100;
A = 16'h0066; B = 16'h0079; #100;
A = 16'h0066; B = 16'h007A; #100;
A = 16'h0066; B = 16'h007B; #100;
A = 16'h0066; B = 16'h007C; #100;
A = 16'h0066; B = 16'h007D; #100;
A = 16'h0066; B = 16'h007E; #100;
A = 16'h0066; B = 16'h007F; #100;
A = 16'h0066; B = 16'h0080; #100;
A = 16'h0066; B = 16'h0081; #100;
A = 16'h0066; B = 16'h0082; #100;
A = 16'h0066; B = 16'h0083; #100;
A = 16'h0066; B = 16'h0084; #100;
A = 16'h0066; B = 16'h0085; #100;
A = 16'h0066; B = 16'h0086; #100;
A = 16'h0066; B = 16'h0087; #100;
A = 16'h0066; B = 16'h0088; #100;
A = 16'h0066; B = 16'h0089; #100;
A = 16'h0066; B = 16'h008A; #100;
A = 16'h0066; B = 16'h008B; #100;
A = 16'h0066; B = 16'h008C; #100;
A = 16'h0066; B = 16'h008D; #100;
A = 16'h0066; B = 16'h008E; #100;
A = 16'h0066; B = 16'h008F; #100;
A = 16'h0066; B = 16'h0090; #100;
A = 16'h0066; B = 16'h0091; #100;
A = 16'h0066; B = 16'h0092; #100;
A = 16'h0066; B = 16'h0093; #100;
A = 16'h0066; B = 16'h0094; #100;
A = 16'h0066; B = 16'h0095; #100;
A = 16'h0066; B = 16'h0096; #100;
A = 16'h0066; B = 16'h0097; #100;
A = 16'h0066; B = 16'h0098; #100;
A = 16'h0066; B = 16'h0099; #100;
A = 16'h0066; B = 16'h009A; #100;
A = 16'h0066; B = 16'h009B; #100;
A = 16'h0066; B = 16'h009C; #100;
A = 16'h0066; B = 16'h009D; #100;
A = 16'h0066; B = 16'h009E; #100;
A = 16'h0066; B = 16'h009F; #100;
A = 16'h0066; B = 16'h00A0; #100;
A = 16'h0066; B = 16'h00A1; #100;
A = 16'h0066; B = 16'h00A2; #100;
A = 16'h0066; B = 16'h00A3; #100;
A = 16'h0066; B = 16'h00A4; #100;
A = 16'h0066; B = 16'h00A5; #100;
A = 16'h0066; B = 16'h00A6; #100;
A = 16'h0066; B = 16'h00A7; #100;
A = 16'h0066; B = 16'h00A8; #100;
A = 16'h0066; B = 16'h00A9; #100;
A = 16'h0066; B = 16'h00AA; #100;
A = 16'h0066; B = 16'h00AB; #100;
A = 16'h0066; B = 16'h00AC; #100;
A = 16'h0066; B = 16'h00AD; #100;
A = 16'h0066; B = 16'h00AE; #100;
A = 16'h0066; B = 16'h00AF; #100;
A = 16'h0066; B = 16'h00B0; #100;
A = 16'h0066; B = 16'h00B1; #100;
A = 16'h0066; B = 16'h00B2; #100;
A = 16'h0066; B = 16'h00B3; #100;
A = 16'h0066; B = 16'h00B4; #100;
A = 16'h0066; B = 16'h00B5; #100;
A = 16'h0066; B = 16'h00B6; #100;
A = 16'h0066; B = 16'h00B7; #100;
A = 16'h0066; B = 16'h00B8; #100;
A = 16'h0066; B = 16'h00B9; #100;
A = 16'h0066; B = 16'h00BA; #100;
A = 16'h0066; B = 16'h00BB; #100;
A = 16'h0066; B = 16'h00BC; #100;
A = 16'h0066; B = 16'h00BD; #100;
A = 16'h0066; B = 16'h00BE; #100;
A = 16'h0066; B = 16'h00BF; #100;
A = 16'h0066; B = 16'h00C0; #100;
A = 16'h0066; B = 16'h00C1; #100;
A = 16'h0066; B = 16'h00C2; #100;
A = 16'h0066; B = 16'h00C3; #100;
A = 16'h0066; B = 16'h00C4; #100;
A = 16'h0066; B = 16'h00C5; #100;
A = 16'h0066; B = 16'h00C6; #100;
A = 16'h0066; B = 16'h00C7; #100;
A = 16'h0066; B = 16'h00C8; #100;
A = 16'h0066; B = 16'h00C9; #100;
A = 16'h0066; B = 16'h00CA; #100;
A = 16'h0066; B = 16'h00CB; #100;
A = 16'h0066; B = 16'h00CC; #100;
A = 16'h0066; B = 16'h00CD; #100;
A = 16'h0066; B = 16'h00CE; #100;
A = 16'h0066; B = 16'h00CF; #100;
A = 16'h0066; B = 16'h00D0; #100;
A = 16'h0066; B = 16'h00D1; #100;
A = 16'h0066; B = 16'h00D2; #100;
A = 16'h0066; B = 16'h00D3; #100;
A = 16'h0066; B = 16'h00D4; #100;
A = 16'h0066; B = 16'h00D5; #100;
A = 16'h0066; B = 16'h00D6; #100;
A = 16'h0066; B = 16'h00D7; #100;
A = 16'h0066; B = 16'h00D8; #100;
A = 16'h0066; B = 16'h00D9; #100;
A = 16'h0066; B = 16'h00DA; #100;
A = 16'h0066; B = 16'h00DB; #100;
A = 16'h0066; B = 16'h00DC; #100;
A = 16'h0066; B = 16'h00DD; #100;
A = 16'h0066; B = 16'h00DE; #100;
A = 16'h0066; B = 16'h00DF; #100;
A = 16'h0066; B = 16'h00E0; #100;
A = 16'h0066; B = 16'h00E1; #100;
A = 16'h0066; B = 16'h00E2; #100;
A = 16'h0066; B = 16'h00E3; #100;
A = 16'h0066; B = 16'h00E4; #100;
A = 16'h0066; B = 16'h00E5; #100;
A = 16'h0066; B = 16'h00E6; #100;
A = 16'h0066; B = 16'h00E7; #100;
A = 16'h0066; B = 16'h00E8; #100;
A = 16'h0066; B = 16'h00E9; #100;
A = 16'h0066; B = 16'h00EA; #100;
A = 16'h0066; B = 16'h00EB; #100;
A = 16'h0066; B = 16'h00EC; #100;
A = 16'h0066; B = 16'h00ED; #100;
A = 16'h0066; B = 16'h00EE; #100;
A = 16'h0066; B = 16'h00EF; #100;
A = 16'h0066; B = 16'h00F0; #100;
A = 16'h0066; B = 16'h00F1; #100;
A = 16'h0066; B = 16'h00F2; #100;
A = 16'h0066; B = 16'h00F3; #100;
A = 16'h0066; B = 16'h00F4; #100;
A = 16'h0066; B = 16'h00F5; #100;
A = 16'h0066; B = 16'h00F6; #100;
A = 16'h0066; B = 16'h00F7; #100;
A = 16'h0066; B = 16'h00F8; #100;
A = 16'h0066; B = 16'h00F9; #100;
A = 16'h0066; B = 16'h00FA; #100;
A = 16'h0066; B = 16'h00FB; #100;
A = 16'h0066; B = 16'h00FC; #100;
A = 16'h0066; B = 16'h00FD; #100;
A = 16'h0066; B = 16'h00FE; #100;
A = 16'h0066; B = 16'h00FF; #100;
A = 16'h0067; B = 16'h000; #100;
A = 16'h0067; B = 16'h001; #100;
A = 16'h0067; B = 16'h002; #100;
A = 16'h0067; B = 16'h003; #100;
A = 16'h0067; B = 16'h004; #100;
A = 16'h0067; B = 16'h005; #100;
A = 16'h0067; B = 16'h006; #100;
A = 16'h0067; B = 16'h007; #100;
A = 16'h0067; B = 16'h008; #100;
A = 16'h0067; B = 16'h009; #100;
A = 16'h0067; B = 16'h00A; #100;
A = 16'h0067; B = 16'h00B; #100;
A = 16'h0067; B = 16'h00C; #100;
A = 16'h0067; B = 16'h00D; #100;
A = 16'h0067; B = 16'h00E; #100;
A = 16'h0067; B = 16'h00F; #100;
A = 16'h0067; B = 16'h0010; #100;
A = 16'h0067; B = 16'h0011; #100;
A = 16'h0067; B = 16'h0012; #100;
A = 16'h0067; B = 16'h0013; #100;
A = 16'h0067; B = 16'h0014; #100;
A = 16'h0067; B = 16'h0015; #100;
A = 16'h0067; B = 16'h0016; #100;
A = 16'h0067; B = 16'h0017; #100;
A = 16'h0067; B = 16'h0018; #100;
A = 16'h0067; B = 16'h0019; #100;
A = 16'h0067; B = 16'h001A; #100;
A = 16'h0067; B = 16'h001B; #100;
A = 16'h0067; B = 16'h001C; #100;
A = 16'h0067; B = 16'h001D; #100;
A = 16'h0067; B = 16'h001E; #100;
A = 16'h0067; B = 16'h001F; #100;
A = 16'h0067; B = 16'h0020; #100;
A = 16'h0067; B = 16'h0021; #100;
A = 16'h0067; B = 16'h0022; #100;
A = 16'h0067; B = 16'h0023; #100;
A = 16'h0067; B = 16'h0024; #100;
A = 16'h0067; B = 16'h0025; #100;
A = 16'h0067; B = 16'h0026; #100;
A = 16'h0067; B = 16'h0027; #100;
A = 16'h0067; B = 16'h0028; #100;
A = 16'h0067; B = 16'h0029; #100;
A = 16'h0067; B = 16'h002A; #100;
A = 16'h0067; B = 16'h002B; #100;
A = 16'h0067; B = 16'h002C; #100;
A = 16'h0067; B = 16'h002D; #100;
A = 16'h0067; B = 16'h002E; #100;
A = 16'h0067; B = 16'h002F; #100;
A = 16'h0067; B = 16'h0030; #100;
A = 16'h0067; B = 16'h0031; #100;
A = 16'h0067; B = 16'h0032; #100;
A = 16'h0067; B = 16'h0033; #100;
A = 16'h0067; B = 16'h0034; #100;
A = 16'h0067; B = 16'h0035; #100;
A = 16'h0067; B = 16'h0036; #100;
A = 16'h0067; B = 16'h0037; #100;
A = 16'h0067; B = 16'h0038; #100;
A = 16'h0067; B = 16'h0039; #100;
A = 16'h0067; B = 16'h003A; #100;
A = 16'h0067; B = 16'h003B; #100;
A = 16'h0067; B = 16'h003C; #100;
A = 16'h0067; B = 16'h003D; #100;
A = 16'h0067; B = 16'h003E; #100;
A = 16'h0067; B = 16'h003F; #100;
A = 16'h0067; B = 16'h0040; #100;
A = 16'h0067; B = 16'h0041; #100;
A = 16'h0067; B = 16'h0042; #100;
A = 16'h0067; B = 16'h0043; #100;
A = 16'h0067; B = 16'h0044; #100;
A = 16'h0067; B = 16'h0045; #100;
A = 16'h0067; B = 16'h0046; #100;
A = 16'h0067; B = 16'h0047; #100;
A = 16'h0067; B = 16'h0048; #100;
A = 16'h0067; B = 16'h0049; #100;
A = 16'h0067; B = 16'h004A; #100;
A = 16'h0067; B = 16'h004B; #100;
A = 16'h0067; B = 16'h004C; #100;
A = 16'h0067; B = 16'h004D; #100;
A = 16'h0067; B = 16'h004E; #100;
A = 16'h0067; B = 16'h004F; #100;
A = 16'h0067; B = 16'h0050; #100;
A = 16'h0067; B = 16'h0051; #100;
A = 16'h0067; B = 16'h0052; #100;
A = 16'h0067; B = 16'h0053; #100;
A = 16'h0067; B = 16'h0054; #100;
A = 16'h0067; B = 16'h0055; #100;
A = 16'h0067; B = 16'h0056; #100;
A = 16'h0067; B = 16'h0057; #100;
A = 16'h0067; B = 16'h0058; #100;
A = 16'h0067; B = 16'h0059; #100;
A = 16'h0067; B = 16'h005A; #100;
A = 16'h0067; B = 16'h005B; #100;
A = 16'h0067; B = 16'h005C; #100;
A = 16'h0067; B = 16'h005D; #100;
A = 16'h0067; B = 16'h005E; #100;
A = 16'h0067; B = 16'h005F; #100;
A = 16'h0067; B = 16'h0060; #100;
A = 16'h0067; B = 16'h0061; #100;
A = 16'h0067; B = 16'h0062; #100;
A = 16'h0067; B = 16'h0063; #100;
A = 16'h0067; B = 16'h0064; #100;
A = 16'h0067; B = 16'h0065; #100;
A = 16'h0067; B = 16'h0066; #100;
A = 16'h0067; B = 16'h0067; #100;
A = 16'h0067; B = 16'h0068; #100;
A = 16'h0067; B = 16'h0069; #100;
A = 16'h0067; B = 16'h006A; #100;
A = 16'h0067; B = 16'h006B; #100;
A = 16'h0067; B = 16'h006C; #100;
A = 16'h0067; B = 16'h006D; #100;
A = 16'h0067; B = 16'h006E; #100;
A = 16'h0067; B = 16'h006F; #100;
A = 16'h0067; B = 16'h0070; #100;
A = 16'h0067; B = 16'h0071; #100;
A = 16'h0067; B = 16'h0072; #100;
A = 16'h0067; B = 16'h0073; #100;
A = 16'h0067; B = 16'h0074; #100;
A = 16'h0067; B = 16'h0075; #100;
A = 16'h0067; B = 16'h0076; #100;
A = 16'h0067; B = 16'h0077; #100;
A = 16'h0067; B = 16'h0078; #100;
A = 16'h0067; B = 16'h0079; #100;
A = 16'h0067; B = 16'h007A; #100;
A = 16'h0067; B = 16'h007B; #100;
A = 16'h0067; B = 16'h007C; #100;
A = 16'h0067; B = 16'h007D; #100;
A = 16'h0067; B = 16'h007E; #100;
A = 16'h0067; B = 16'h007F; #100;
A = 16'h0067; B = 16'h0080; #100;
A = 16'h0067; B = 16'h0081; #100;
A = 16'h0067; B = 16'h0082; #100;
A = 16'h0067; B = 16'h0083; #100;
A = 16'h0067; B = 16'h0084; #100;
A = 16'h0067; B = 16'h0085; #100;
A = 16'h0067; B = 16'h0086; #100;
A = 16'h0067; B = 16'h0087; #100;
A = 16'h0067; B = 16'h0088; #100;
A = 16'h0067; B = 16'h0089; #100;
A = 16'h0067; B = 16'h008A; #100;
A = 16'h0067; B = 16'h008B; #100;
A = 16'h0067; B = 16'h008C; #100;
A = 16'h0067; B = 16'h008D; #100;
A = 16'h0067; B = 16'h008E; #100;
A = 16'h0067; B = 16'h008F; #100;
A = 16'h0067; B = 16'h0090; #100;
A = 16'h0067; B = 16'h0091; #100;
A = 16'h0067; B = 16'h0092; #100;
A = 16'h0067; B = 16'h0093; #100;
A = 16'h0067; B = 16'h0094; #100;
A = 16'h0067; B = 16'h0095; #100;
A = 16'h0067; B = 16'h0096; #100;
A = 16'h0067; B = 16'h0097; #100;
A = 16'h0067; B = 16'h0098; #100;
A = 16'h0067; B = 16'h0099; #100;
A = 16'h0067; B = 16'h009A; #100;
A = 16'h0067; B = 16'h009B; #100;
A = 16'h0067; B = 16'h009C; #100;
A = 16'h0067; B = 16'h009D; #100;
A = 16'h0067; B = 16'h009E; #100;
A = 16'h0067; B = 16'h009F; #100;
A = 16'h0067; B = 16'h00A0; #100;
A = 16'h0067; B = 16'h00A1; #100;
A = 16'h0067; B = 16'h00A2; #100;
A = 16'h0067; B = 16'h00A3; #100;
A = 16'h0067; B = 16'h00A4; #100;
A = 16'h0067; B = 16'h00A5; #100;
A = 16'h0067; B = 16'h00A6; #100;
A = 16'h0067; B = 16'h00A7; #100;
A = 16'h0067; B = 16'h00A8; #100;
A = 16'h0067; B = 16'h00A9; #100;
A = 16'h0067; B = 16'h00AA; #100;
A = 16'h0067; B = 16'h00AB; #100;
A = 16'h0067; B = 16'h00AC; #100;
A = 16'h0067; B = 16'h00AD; #100;
A = 16'h0067; B = 16'h00AE; #100;
A = 16'h0067; B = 16'h00AF; #100;
A = 16'h0067; B = 16'h00B0; #100;
A = 16'h0067; B = 16'h00B1; #100;
A = 16'h0067; B = 16'h00B2; #100;
A = 16'h0067; B = 16'h00B3; #100;
A = 16'h0067; B = 16'h00B4; #100;
A = 16'h0067; B = 16'h00B5; #100;
A = 16'h0067; B = 16'h00B6; #100;
A = 16'h0067; B = 16'h00B7; #100;
A = 16'h0067; B = 16'h00B8; #100;
A = 16'h0067; B = 16'h00B9; #100;
A = 16'h0067; B = 16'h00BA; #100;
A = 16'h0067; B = 16'h00BB; #100;
A = 16'h0067; B = 16'h00BC; #100;
A = 16'h0067; B = 16'h00BD; #100;
A = 16'h0067; B = 16'h00BE; #100;
A = 16'h0067; B = 16'h00BF; #100;
A = 16'h0067; B = 16'h00C0; #100;
A = 16'h0067; B = 16'h00C1; #100;
A = 16'h0067; B = 16'h00C2; #100;
A = 16'h0067; B = 16'h00C3; #100;
A = 16'h0067; B = 16'h00C4; #100;
A = 16'h0067; B = 16'h00C5; #100;
A = 16'h0067; B = 16'h00C6; #100;
A = 16'h0067; B = 16'h00C7; #100;
A = 16'h0067; B = 16'h00C8; #100;
A = 16'h0067; B = 16'h00C9; #100;
A = 16'h0067; B = 16'h00CA; #100;
A = 16'h0067; B = 16'h00CB; #100;
A = 16'h0067; B = 16'h00CC; #100;
A = 16'h0067; B = 16'h00CD; #100;
A = 16'h0067; B = 16'h00CE; #100;
A = 16'h0067; B = 16'h00CF; #100;
A = 16'h0067; B = 16'h00D0; #100;
A = 16'h0067; B = 16'h00D1; #100;
A = 16'h0067; B = 16'h00D2; #100;
A = 16'h0067; B = 16'h00D3; #100;
A = 16'h0067; B = 16'h00D4; #100;
A = 16'h0067; B = 16'h00D5; #100;
A = 16'h0067; B = 16'h00D6; #100;
A = 16'h0067; B = 16'h00D7; #100;
A = 16'h0067; B = 16'h00D8; #100;
A = 16'h0067; B = 16'h00D9; #100;
A = 16'h0067; B = 16'h00DA; #100;
A = 16'h0067; B = 16'h00DB; #100;
A = 16'h0067; B = 16'h00DC; #100;
A = 16'h0067; B = 16'h00DD; #100;
A = 16'h0067; B = 16'h00DE; #100;
A = 16'h0067; B = 16'h00DF; #100;
A = 16'h0067; B = 16'h00E0; #100;
A = 16'h0067; B = 16'h00E1; #100;
A = 16'h0067; B = 16'h00E2; #100;
A = 16'h0067; B = 16'h00E3; #100;
A = 16'h0067; B = 16'h00E4; #100;
A = 16'h0067; B = 16'h00E5; #100;
A = 16'h0067; B = 16'h00E6; #100;
A = 16'h0067; B = 16'h00E7; #100;
A = 16'h0067; B = 16'h00E8; #100;
A = 16'h0067; B = 16'h00E9; #100;
A = 16'h0067; B = 16'h00EA; #100;
A = 16'h0067; B = 16'h00EB; #100;
A = 16'h0067; B = 16'h00EC; #100;
A = 16'h0067; B = 16'h00ED; #100;
A = 16'h0067; B = 16'h00EE; #100;
A = 16'h0067; B = 16'h00EF; #100;
A = 16'h0067; B = 16'h00F0; #100;
A = 16'h0067; B = 16'h00F1; #100;
A = 16'h0067; B = 16'h00F2; #100;
A = 16'h0067; B = 16'h00F3; #100;
A = 16'h0067; B = 16'h00F4; #100;
A = 16'h0067; B = 16'h00F5; #100;
A = 16'h0067; B = 16'h00F6; #100;
A = 16'h0067; B = 16'h00F7; #100;
A = 16'h0067; B = 16'h00F8; #100;
A = 16'h0067; B = 16'h00F9; #100;
A = 16'h0067; B = 16'h00FA; #100;
A = 16'h0067; B = 16'h00FB; #100;
A = 16'h0067; B = 16'h00FC; #100;
A = 16'h0067; B = 16'h00FD; #100;
A = 16'h0067; B = 16'h00FE; #100;
A = 16'h0067; B = 16'h00FF; #100;
A = 16'h0068; B = 16'h000; #100;
A = 16'h0068; B = 16'h001; #100;
A = 16'h0068; B = 16'h002; #100;
A = 16'h0068; B = 16'h003; #100;
A = 16'h0068; B = 16'h004; #100;
A = 16'h0068; B = 16'h005; #100;
A = 16'h0068; B = 16'h006; #100;
A = 16'h0068; B = 16'h007; #100;
A = 16'h0068; B = 16'h008; #100;
A = 16'h0068; B = 16'h009; #100;
A = 16'h0068; B = 16'h00A; #100;
A = 16'h0068; B = 16'h00B; #100;
A = 16'h0068; B = 16'h00C; #100;
A = 16'h0068; B = 16'h00D; #100;
A = 16'h0068; B = 16'h00E; #100;
A = 16'h0068; B = 16'h00F; #100;
A = 16'h0068; B = 16'h0010; #100;
A = 16'h0068; B = 16'h0011; #100;
A = 16'h0068; B = 16'h0012; #100;
A = 16'h0068; B = 16'h0013; #100;
A = 16'h0068; B = 16'h0014; #100;
A = 16'h0068; B = 16'h0015; #100;
A = 16'h0068; B = 16'h0016; #100;
A = 16'h0068; B = 16'h0017; #100;
A = 16'h0068; B = 16'h0018; #100;
A = 16'h0068; B = 16'h0019; #100;
A = 16'h0068; B = 16'h001A; #100;
A = 16'h0068; B = 16'h001B; #100;
A = 16'h0068; B = 16'h001C; #100;
A = 16'h0068; B = 16'h001D; #100;
A = 16'h0068; B = 16'h001E; #100;
A = 16'h0068; B = 16'h001F; #100;
A = 16'h0068; B = 16'h0020; #100;
A = 16'h0068; B = 16'h0021; #100;
A = 16'h0068; B = 16'h0022; #100;
A = 16'h0068; B = 16'h0023; #100;
A = 16'h0068; B = 16'h0024; #100;
A = 16'h0068; B = 16'h0025; #100;
A = 16'h0068; B = 16'h0026; #100;
A = 16'h0068; B = 16'h0027; #100;
A = 16'h0068; B = 16'h0028; #100;
A = 16'h0068; B = 16'h0029; #100;
A = 16'h0068; B = 16'h002A; #100;
A = 16'h0068; B = 16'h002B; #100;
A = 16'h0068; B = 16'h002C; #100;
A = 16'h0068; B = 16'h002D; #100;
A = 16'h0068; B = 16'h002E; #100;
A = 16'h0068; B = 16'h002F; #100;
A = 16'h0068; B = 16'h0030; #100;
A = 16'h0068; B = 16'h0031; #100;
A = 16'h0068; B = 16'h0032; #100;
A = 16'h0068; B = 16'h0033; #100;
A = 16'h0068; B = 16'h0034; #100;
A = 16'h0068; B = 16'h0035; #100;
A = 16'h0068; B = 16'h0036; #100;
A = 16'h0068; B = 16'h0037; #100;
A = 16'h0068; B = 16'h0038; #100;
A = 16'h0068; B = 16'h0039; #100;
A = 16'h0068; B = 16'h003A; #100;
A = 16'h0068; B = 16'h003B; #100;
A = 16'h0068; B = 16'h003C; #100;
A = 16'h0068; B = 16'h003D; #100;
A = 16'h0068; B = 16'h003E; #100;
A = 16'h0068; B = 16'h003F; #100;
A = 16'h0068; B = 16'h0040; #100;
A = 16'h0068; B = 16'h0041; #100;
A = 16'h0068; B = 16'h0042; #100;
A = 16'h0068; B = 16'h0043; #100;
A = 16'h0068; B = 16'h0044; #100;
A = 16'h0068; B = 16'h0045; #100;
A = 16'h0068; B = 16'h0046; #100;
A = 16'h0068; B = 16'h0047; #100;
A = 16'h0068; B = 16'h0048; #100;
A = 16'h0068; B = 16'h0049; #100;
A = 16'h0068; B = 16'h004A; #100;
A = 16'h0068; B = 16'h004B; #100;
A = 16'h0068; B = 16'h004C; #100;
A = 16'h0068; B = 16'h004D; #100;
A = 16'h0068; B = 16'h004E; #100;
A = 16'h0068; B = 16'h004F; #100;
A = 16'h0068; B = 16'h0050; #100;
A = 16'h0068; B = 16'h0051; #100;
A = 16'h0068; B = 16'h0052; #100;
A = 16'h0068; B = 16'h0053; #100;
A = 16'h0068; B = 16'h0054; #100;
A = 16'h0068; B = 16'h0055; #100;
A = 16'h0068; B = 16'h0056; #100;
A = 16'h0068; B = 16'h0057; #100;
A = 16'h0068; B = 16'h0058; #100;
A = 16'h0068; B = 16'h0059; #100;
A = 16'h0068; B = 16'h005A; #100;
A = 16'h0068; B = 16'h005B; #100;
A = 16'h0068; B = 16'h005C; #100;
A = 16'h0068; B = 16'h005D; #100;
A = 16'h0068; B = 16'h005E; #100;
A = 16'h0068; B = 16'h005F; #100;
A = 16'h0068; B = 16'h0060; #100;
A = 16'h0068; B = 16'h0061; #100;
A = 16'h0068; B = 16'h0062; #100;
A = 16'h0068; B = 16'h0063; #100;
A = 16'h0068; B = 16'h0064; #100;
A = 16'h0068; B = 16'h0065; #100;
A = 16'h0068; B = 16'h0066; #100;
A = 16'h0068; B = 16'h0067; #100;
A = 16'h0068; B = 16'h0068; #100;
A = 16'h0068; B = 16'h0069; #100;
A = 16'h0068; B = 16'h006A; #100;
A = 16'h0068; B = 16'h006B; #100;
A = 16'h0068; B = 16'h006C; #100;
A = 16'h0068; B = 16'h006D; #100;
A = 16'h0068; B = 16'h006E; #100;
A = 16'h0068; B = 16'h006F; #100;
A = 16'h0068; B = 16'h0070; #100;
A = 16'h0068; B = 16'h0071; #100;
A = 16'h0068; B = 16'h0072; #100;
A = 16'h0068; B = 16'h0073; #100;
A = 16'h0068; B = 16'h0074; #100;
A = 16'h0068; B = 16'h0075; #100;
A = 16'h0068; B = 16'h0076; #100;
A = 16'h0068; B = 16'h0077; #100;
A = 16'h0068; B = 16'h0078; #100;
A = 16'h0068; B = 16'h0079; #100;
A = 16'h0068; B = 16'h007A; #100;
A = 16'h0068; B = 16'h007B; #100;
A = 16'h0068; B = 16'h007C; #100;
A = 16'h0068; B = 16'h007D; #100;
A = 16'h0068; B = 16'h007E; #100;
A = 16'h0068; B = 16'h007F; #100;
A = 16'h0068; B = 16'h0080; #100;
A = 16'h0068; B = 16'h0081; #100;
A = 16'h0068; B = 16'h0082; #100;
A = 16'h0068; B = 16'h0083; #100;
A = 16'h0068; B = 16'h0084; #100;
A = 16'h0068; B = 16'h0085; #100;
A = 16'h0068; B = 16'h0086; #100;
A = 16'h0068; B = 16'h0087; #100;
A = 16'h0068; B = 16'h0088; #100;
A = 16'h0068; B = 16'h0089; #100;
A = 16'h0068; B = 16'h008A; #100;
A = 16'h0068; B = 16'h008B; #100;
A = 16'h0068; B = 16'h008C; #100;
A = 16'h0068; B = 16'h008D; #100;
A = 16'h0068; B = 16'h008E; #100;
A = 16'h0068; B = 16'h008F; #100;
A = 16'h0068; B = 16'h0090; #100;
A = 16'h0068; B = 16'h0091; #100;
A = 16'h0068; B = 16'h0092; #100;
A = 16'h0068; B = 16'h0093; #100;
A = 16'h0068; B = 16'h0094; #100;
A = 16'h0068; B = 16'h0095; #100;
A = 16'h0068; B = 16'h0096; #100;
A = 16'h0068; B = 16'h0097; #100;
A = 16'h0068; B = 16'h0098; #100;
A = 16'h0068; B = 16'h0099; #100;
A = 16'h0068; B = 16'h009A; #100;
A = 16'h0068; B = 16'h009B; #100;
A = 16'h0068; B = 16'h009C; #100;
A = 16'h0068; B = 16'h009D; #100;
A = 16'h0068; B = 16'h009E; #100;
A = 16'h0068; B = 16'h009F; #100;
A = 16'h0068; B = 16'h00A0; #100;
A = 16'h0068; B = 16'h00A1; #100;
A = 16'h0068; B = 16'h00A2; #100;
A = 16'h0068; B = 16'h00A3; #100;
A = 16'h0068; B = 16'h00A4; #100;
A = 16'h0068; B = 16'h00A5; #100;
A = 16'h0068; B = 16'h00A6; #100;
A = 16'h0068; B = 16'h00A7; #100;
A = 16'h0068; B = 16'h00A8; #100;
A = 16'h0068; B = 16'h00A9; #100;
A = 16'h0068; B = 16'h00AA; #100;
A = 16'h0068; B = 16'h00AB; #100;
A = 16'h0068; B = 16'h00AC; #100;
A = 16'h0068; B = 16'h00AD; #100;
A = 16'h0068; B = 16'h00AE; #100;
A = 16'h0068; B = 16'h00AF; #100;
A = 16'h0068; B = 16'h00B0; #100;
A = 16'h0068; B = 16'h00B1; #100;
A = 16'h0068; B = 16'h00B2; #100;
A = 16'h0068; B = 16'h00B3; #100;
A = 16'h0068; B = 16'h00B4; #100;
A = 16'h0068; B = 16'h00B5; #100;
A = 16'h0068; B = 16'h00B6; #100;
A = 16'h0068; B = 16'h00B7; #100;
A = 16'h0068; B = 16'h00B8; #100;
A = 16'h0068; B = 16'h00B9; #100;
A = 16'h0068; B = 16'h00BA; #100;
A = 16'h0068; B = 16'h00BB; #100;
A = 16'h0068; B = 16'h00BC; #100;
A = 16'h0068; B = 16'h00BD; #100;
A = 16'h0068; B = 16'h00BE; #100;
A = 16'h0068; B = 16'h00BF; #100;
A = 16'h0068; B = 16'h00C0; #100;
A = 16'h0068; B = 16'h00C1; #100;
A = 16'h0068; B = 16'h00C2; #100;
A = 16'h0068; B = 16'h00C3; #100;
A = 16'h0068; B = 16'h00C4; #100;
A = 16'h0068; B = 16'h00C5; #100;
A = 16'h0068; B = 16'h00C6; #100;
A = 16'h0068; B = 16'h00C7; #100;
A = 16'h0068; B = 16'h00C8; #100;
A = 16'h0068; B = 16'h00C9; #100;
A = 16'h0068; B = 16'h00CA; #100;
A = 16'h0068; B = 16'h00CB; #100;
A = 16'h0068; B = 16'h00CC; #100;
A = 16'h0068; B = 16'h00CD; #100;
A = 16'h0068; B = 16'h00CE; #100;
A = 16'h0068; B = 16'h00CF; #100;
A = 16'h0068; B = 16'h00D0; #100;
A = 16'h0068; B = 16'h00D1; #100;
A = 16'h0068; B = 16'h00D2; #100;
A = 16'h0068; B = 16'h00D3; #100;
A = 16'h0068; B = 16'h00D4; #100;
A = 16'h0068; B = 16'h00D5; #100;
A = 16'h0068; B = 16'h00D6; #100;
A = 16'h0068; B = 16'h00D7; #100;
A = 16'h0068; B = 16'h00D8; #100;
A = 16'h0068; B = 16'h00D9; #100;
A = 16'h0068; B = 16'h00DA; #100;
A = 16'h0068; B = 16'h00DB; #100;
A = 16'h0068; B = 16'h00DC; #100;
A = 16'h0068; B = 16'h00DD; #100;
A = 16'h0068; B = 16'h00DE; #100;
A = 16'h0068; B = 16'h00DF; #100;
A = 16'h0068; B = 16'h00E0; #100;
A = 16'h0068; B = 16'h00E1; #100;
A = 16'h0068; B = 16'h00E2; #100;
A = 16'h0068; B = 16'h00E3; #100;
A = 16'h0068; B = 16'h00E4; #100;
A = 16'h0068; B = 16'h00E5; #100;
A = 16'h0068; B = 16'h00E6; #100;
A = 16'h0068; B = 16'h00E7; #100;
A = 16'h0068; B = 16'h00E8; #100;
A = 16'h0068; B = 16'h00E9; #100;
A = 16'h0068; B = 16'h00EA; #100;
A = 16'h0068; B = 16'h00EB; #100;
A = 16'h0068; B = 16'h00EC; #100;
A = 16'h0068; B = 16'h00ED; #100;
A = 16'h0068; B = 16'h00EE; #100;
A = 16'h0068; B = 16'h00EF; #100;
A = 16'h0068; B = 16'h00F0; #100;
A = 16'h0068; B = 16'h00F1; #100;
A = 16'h0068; B = 16'h00F2; #100;
A = 16'h0068; B = 16'h00F3; #100;
A = 16'h0068; B = 16'h00F4; #100;
A = 16'h0068; B = 16'h00F5; #100;
A = 16'h0068; B = 16'h00F6; #100;
A = 16'h0068; B = 16'h00F7; #100;
A = 16'h0068; B = 16'h00F8; #100;
A = 16'h0068; B = 16'h00F9; #100;
A = 16'h0068; B = 16'h00FA; #100;
A = 16'h0068; B = 16'h00FB; #100;
A = 16'h0068; B = 16'h00FC; #100;
A = 16'h0068; B = 16'h00FD; #100;
A = 16'h0068; B = 16'h00FE; #100;
A = 16'h0068; B = 16'h00FF; #100;
A = 16'h0069; B = 16'h000; #100;
A = 16'h0069; B = 16'h001; #100;
A = 16'h0069; B = 16'h002; #100;
A = 16'h0069; B = 16'h003; #100;
A = 16'h0069; B = 16'h004; #100;
A = 16'h0069; B = 16'h005; #100;
A = 16'h0069; B = 16'h006; #100;
A = 16'h0069; B = 16'h007; #100;
A = 16'h0069; B = 16'h008; #100;
A = 16'h0069; B = 16'h009; #100;
A = 16'h0069; B = 16'h00A; #100;
A = 16'h0069; B = 16'h00B; #100;
A = 16'h0069; B = 16'h00C; #100;
A = 16'h0069; B = 16'h00D; #100;
A = 16'h0069; B = 16'h00E; #100;
A = 16'h0069; B = 16'h00F; #100;
A = 16'h0069; B = 16'h0010; #100;
A = 16'h0069; B = 16'h0011; #100;
A = 16'h0069; B = 16'h0012; #100;
A = 16'h0069; B = 16'h0013; #100;
A = 16'h0069; B = 16'h0014; #100;
A = 16'h0069; B = 16'h0015; #100;
A = 16'h0069; B = 16'h0016; #100;
A = 16'h0069; B = 16'h0017; #100;
A = 16'h0069; B = 16'h0018; #100;
A = 16'h0069; B = 16'h0019; #100;
A = 16'h0069; B = 16'h001A; #100;
A = 16'h0069; B = 16'h001B; #100;
A = 16'h0069; B = 16'h001C; #100;
A = 16'h0069; B = 16'h001D; #100;
A = 16'h0069; B = 16'h001E; #100;
A = 16'h0069; B = 16'h001F; #100;
A = 16'h0069; B = 16'h0020; #100;
A = 16'h0069; B = 16'h0021; #100;
A = 16'h0069; B = 16'h0022; #100;
A = 16'h0069; B = 16'h0023; #100;
A = 16'h0069; B = 16'h0024; #100;
A = 16'h0069; B = 16'h0025; #100;
A = 16'h0069; B = 16'h0026; #100;
A = 16'h0069; B = 16'h0027; #100;
A = 16'h0069; B = 16'h0028; #100;
A = 16'h0069; B = 16'h0029; #100;
A = 16'h0069; B = 16'h002A; #100;
A = 16'h0069; B = 16'h002B; #100;
A = 16'h0069; B = 16'h002C; #100;
A = 16'h0069; B = 16'h002D; #100;
A = 16'h0069; B = 16'h002E; #100;
A = 16'h0069; B = 16'h002F; #100;
A = 16'h0069; B = 16'h0030; #100;
A = 16'h0069; B = 16'h0031; #100;
A = 16'h0069; B = 16'h0032; #100;
A = 16'h0069; B = 16'h0033; #100;
A = 16'h0069; B = 16'h0034; #100;
A = 16'h0069; B = 16'h0035; #100;
A = 16'h0069; B = 16'h0036; #100;
A = 16'h0069; B = 16'h0037; #100;
A = 16'h0069; B = 16'h0038; #100;
A = 16'h0069; B = 16'h0039; #100;
A = 16'h0069; B = 16'h003A; #100;
A = 16'h0069; B = 16'h003B; #100;
A = 16'h0069; B = 16'h003C; #100;
A = 16'h0069; B = 16'h003D; #100;
A = 16'h0069; B = 16'h003E; #100;
A = 16'h0069; B = 16'h003F; #100;
A = 16'h0069; B = 16'h0040; #100;
A = 16'h0069; B = 16'h0041; #100;
A = 16'h0069; B = 16'h0042; #100;
A = 16'h0069; B = 16'h0043; #100;
A = 16'h0069; B = 16'h0044; #100;
A = 16'h0069; B = 16'h0045; #100;
A = 16'h0069; B = 16'h0046; #100;
A = 16'h0069; B = 16'h0047; #100;
A = 16'h0069; B = 16'h0048; #100;
A = 16'h0069; B = 16'h0049; #100;
A = 16'h0069; B = 16'h004A; #100;
A = 16'h0069; B = 16'h004B; #100;
A = 16'h0069; B = 16'h004C; #100;
A = 16'h0069; B = 16'h004D; #100;
A = 16'h0069; B = 16'h004E; #100;
A = 16'h0069; B = 16'h004F; #100;
A = 16'h0069; B = 16'h0050; #100;
A = 16'h0069; B = 16'h0051; #100;
A = 16'h0069; B = 16'h0052; #100;
A = 16'h0069; B = 16'h0053; #100;
A = 16'h0069; B = 16'h0054; #100;
A = 16'h0069; B = 16'h0055; #100;
A = 16'h0069; B = 16'h0056; #100;
A = 16'h0069; B = 16'h0057; #100;
A = 16'h0069; B = 16'h0058; #100;
A = 16'h0069; B = 16'h0059; #100;
A = 16'h0069; B = 16'h005A; #100;
A = 16'h0069; B = 16'h005B; #100;
A = 16'h0069; B = 16'h005C; #100;
A = 16'h0069; B = 16'h005D; #100;
A = 16'h0069; B = 16'h005E; #100;
A = 16'h0069; B = 16'h005F; #100;
A = 16'h0069; B = 16'h0060; #100;
A = 16'h0069; B = 16'h0061; #100;
A = 16'h0069; B = 16'h0062; #100;
A = 16'h0069; B = 16'h0063; #100;
A = 16'h0069; B = 16'h0064; #100;
A = 16'h0069; B = 16'h0065; #100;
A = 16'h0069; B = 16'h0066; #100;
A = 16'h0069; B = 16'h0067; #100;
A = 16'h0069; B = 16'h0068; #100;
A = 16'h0069; B = 16'h0069; #100;
A = 16'h0069; B = 16'h006A; #100;
A = 16'h0069; B = 16'h006B; #100;
A = 16'h0069; B = 16'h006C; #100;
A = 16'h0069; B = 16'h006D; #100;
A = 16'h0069; B = 16'h006E; #100;
A = 16'h0069; B = 16'h006F; #100;
A = 16'h0069; B = 16'h0070; #100;
A = 16'h0069; B = 16'h0071; #100;
A = 16'h0069; B = 16'h0072; #100;
A = 16'h0069; B = 16'h0073; #100;
A = 16'h0069; B = 16'h0074; #100;
A = 16'h0069; B = 16'h0075; #100;
A = 16'h0069; B = 16'h0076; #100;
A = 16'h0069; B = 16'h0077; #100;
A = 16'h0069; B = 16'h0078; #100;
A = 16'h0069; B = 16'h0079; #100;
A = 16'h0069; B = 16'h007A; #100;
A = 16'h0069; B = 16'h007B; #100;
A = 16'h0069; B = 16'h007C; #100;
A = 16'h0069; B = 16'h007D; #100;
A = 16'h0069; B = 16'h007E; #100;
A = 16'h0069; B = 16'h007F; #100;
A = 16'h0069; B = 16'h0080; #100;
A = 16'h0069; B = 16'h0081; #100;
A = 16'h0069; B = 16'h0082; #100;
A = 16'h0069; B = 16'h0083; #100;
A = 16'h0069; B = 16'h0084; #100;
A = 16'h0069; B = 16'h0085; #100;
A = 16'h0069; B = 16'h0086; #100;
A = 16'h0069; B = 16'h0087; #100;
A = 16'h0069; B = 16'h0088; #100;
A = 16'h0069; B = 16'h0089; #100;
A = 16'h0069; B = 16'h008A; #100;
A = 16'h0069; B = 16'h008B; #100;
A = 16'h0069; B = 16'h008C; #100;
A = 16'h0069; B = 16'h008D; #100;
A = 16'h0069; B = 16'h008E; #100;
A = 16'h0069; B = 16'h008F; #100;
A = 16'h0069; B = 16'h0090; #100;
A = 16'h0069; B = 16'h0091; #100;
A = 16'h0069; B = 16'h0092; #100;
A = 16'h0069; B = 16'h0093; #100;
A = 16'h0069; B = 16'h0094; #100;
A = 16'h0069; B = 16'h0095; #100;
A = 16'h0069; B = 16'h0096; #100;
A = 16'h0069; B = 16'h0097; #100;
A = 16'h0069; B = 16'h0098; #100;
A = 16'h0069; B = 16'h0099; #100;
A = 16'h0069; B = 16'h009A; #100;
A = 16'h0069; B = 16'h009B; #100;
A = 16'h0069; B = 16'h009C; #100;
A = 16'h0069; B = 16'h009D; #100;
A = 16'h0069; B = 16'h009E; #100;
A = 16'h0069; B = 16'h009F; #100;
A = 16'h0069; B = 16'h00A0; #100;
A = 16'h0069; B = 16'h00A1; #100;
A = 16'h0069; B = 16'h00A2; #100;
A = 16'h0069; B = 16'h00A3; #100;
A = 16'h0069; B = 16'h00A4; #100;
A = 16'h0069; B = 16'h00A5; #100;
A = 16'h0069; B = 16'h00A6; #100;
A = 16'h0069; B = 16'h00A7; #100;
A = 16'h0069; B = 16'h00A8; #100;
A = 16'h0069; B = 16'h00A9; #100;
A = 16'h0069; B = 16'h00AA; #100;
A = 16'h0069; B = 16'h00AB; #100;
A = 16'h0069; B = 16'h00AC; #100;
A = 16'h0069; B = 16'h00AD; #100;
A = 16'h0069; B = 16'h00AE; #100;
A = 16'h0069; B = 16'h00AF; #100;
A = 16'h0069; B = 16'h00B0; #100;
A = 16'h0069; B = 16'h00B1; #100;
A = 16'h0069; B = 16'h00B2; #100;
A = 16'h0069; B = 16'h00B3; #100;
A = 16'h0069; B = 16'h00B4; #100;
A = 16'h0069; B = 16'h00B5; #100;
A = 16'h0069; B = 16'h00B6; #100;
A = 16'h0069; B = 16'h00B7; #100;
A = 16'h0069; B = 16'h00B8; #100;
A = 16'h0069; B = 16'h00B9; #100;
A = 16'h0069; B = 16'h00BA; #100;
A = 16'h0069; B = 16'h00BB; #100;
A = 16'h0069; B = 16'h00BC; #100;
A = 16'h0069; B = 16'h00BD; #100;
A = 16'h0069; B = 16'h00BE; #100;
A = 16'h0069; B = 16'h00BF; #100;
A = 16'h0069; B = 16'h00C0; #100;
A = 16'h0069; B = 16'h00C1; #100;
A = 16'h0069; B = 16'h00C2; #100;
A = 16'h0069; B = 16'h00C3; #100;
A = 16'h0069; B = 16'h00C4; #100;
A = 16'h0069; B = 16'h00C5; #100;
A = 16'h0069; B = 16'h00C6; #100;
A = 16'h0069; B = 16'h00C7; #100;
A = 16'h0069; B = 16'h00C8; #100;
A = 16'h0069; B = 16'h00C9; #100;
A = 16'h0069; B = 16'h00CA; #100;
A = 16'h0069; B = 16'h00CB; #100;
A = 16'h0069; B = 16'h00CC; #100;
A = 16'h0069; B = 16'h00CD; #100;
A = 16'h0069; B = 16'h00CE; #100;
A = 16'h0069; B = 16'h00CF; #100;
A = 16'h0069; B = 16'h00D0; #100;
A = 16'h0069; B = 16'h00D1; #100;
A = 16'h0069; B = 16'h00D2; #100;
A = 16'h0069; B = 16'h00D3; #100;
A = 16'h0069; B = 16'h00D4; #100;
A = 16'h0069; B = 16'h00D5; #100;
A = 16'h0069; B = 16'h00D6; #100;
A = 16'h0069; B = 16'h00D7; #100;
A = 16'h0069; B = 16'h00D8; #100;
A = 16'h0069; B = 16'h00D9; #100;
A = 16'h0069; B = 16'h00DA; #100;
A = 16'h0069; B = 16'h00DB; #100;
A = 16'h0069; B = 16'h00DC; #100;
A = 16'h0069; B = 16'h00DD; #100;
A = 16'h0069; B = 16'h00DE; #100;
A = 16'h0069; B = 16'h00DF; #100;
A = 16'h0069; B = 16'h00E0; #100;
A = 16'h0069; B = 16'h00E1; #100;
A = 16'h0069; B = 16'h00E2; #100;
A = 16'h0069; B = 16'h00E3; #100;
A = 16'h0069; B = 16'h00E4; #100;
A = 16'h0069; B = 16'h00E5; #100;
A = 16'h0069; B = 16'h00E6; #100;
A = 16'h0069; B = 16'h00E7; #100;
A = 16'h0069; B = 16'h00E8; #100;
A = 16'h0069; B = 16'h00E9; #100;
A = 16'h0069; B = 16'h00EA; #100;
A = 16'h0069; B = 16'h00EB; #100;
A = 16'h0069; B = 16'h00EC; #100;
A = 16'h0069; B = 16'h00ED; #100;
A = 16'h0069; B = 16'h00EE; #100;
A = 16'h0069; B = 16'h00EF; #100;
A = 16'h0069; B = 16'h00F0; #100;
A = 16'h0069; B = 16'h00F1; #100;
A = 16'h0069; B = 16'h00F2; #100;
A = 16'h0069; B = 16'h00F3; #100;
A = 16'h0069; B = 16'h00F4; #100;
A = 16'h0069; B = 16'h00F5; #100;
A = 16'h0069; B = 16'h00F6; #100;
A = 16'h0069; B = 16'h00F7; #100;
A = 16'h0069; B = 16'h00F8; #100;
A = 16'h0069; B = 16'h00F9; #100;
A = 16'h0069; B = 16'h00FA; #100;
A = 16'h0069; B = 16'h00FB; #100;
A = 16'h0069; B = 16'h00FC; #100;
A = 16'h0069; B = 16'h00FD; #100;
A = 16'h0069; B = 16'h00FE; #100;
A = 16'h0069; B = 16'h00FF; #100;
A = 16'h006A; B = 16'h000; #100;
A = 16'h006A; B = 16'h001; #100;
A = 16'h006A; B = 16'h002; #100;
A = 16'h006A; B = 16'h003; #100;
A = 16'h006A; B = 16'h004; #100;
A = 16'h006A; B = 16'h005; #100;
A = 16'h006A; B = 16'h006; #100;
A = 16'h006A; B = 16'h007; #100;
A = 16'h006A; B = 16'h008; #100;
A = 16'h006A; B = 16'h009; #100;
A = 16'h006A; B = 16'h00A; #100;
A = 16'h006A; B = 16'h00B; #100;
A = 16'h006A; B = 16'h00C; #100;
A = 16'h006A; B = 16'h00D; #100;
A = 16'h006A; B = 16'h00E; #100;
A = 16'h006A; B = 16'h00F; #100;
A = 16'h006A; B = 16'h0010; #100;
A = 16'h006A; B = 16'h0011; #100;
A = 16'h006A; B = 16'h0012; #100;
A = 16'h006A; B = 16'h0013; #100;
A = 16'h006A; B = 16'h0014; #100;
A = 16'h006A; B = 16'h0015; #100;
A = 16'h006A; B = 16'h0016; #100;
A = 16'h006A; B = 16'h0017; #100;
A = 16'h006A; B = 16'h0018; #100;
A = 16'h006A; B = 16'h0019; #100;
A = 16'h006A; B = 16'h001A; #100;
A = 16'h006A; B = 16'h001B; #100;
A = 16'h006A; B = 16'h001C; #100;
A = 16'h006A; B = 16'h001D; #100;
A = 16'h006A; B = 16'h001E; #100;
A = 16'h006A; B = 16'h001F; #100;
A = 16'h006A; B = 16'h0020; #100;
A = 16'h006A; B = 16'h0021; #100;
A = 16'h006A; B = 16'h0022; #100;
A = 16'h006A; B = 16'h0023; #100;
A = 16'h006A; B = 16'h0024; #100;
A = 16'h006A; B = 16'h0025; #100;
A = 16'h006A; B = 16'h0026; #100;
A = 16'h006A; B = 16'h0027; #100;
A = 16'h006A; B = 16'h0028; #100;
A = 16'h006A; B = 16'h0029; #100;
A = 16'h006A; B = 16'h002A; #100;
A = 16'h006A; B = 16'h002B; #100;
A = 16'h006A; B = 16'h002C; #100;
A = 16'h006A; B = 16'h002D; #100;
A = 16'h006A; B = 16'h002E; #100;
A = 16'h006A; B = 16'h002F; #100;
A = 16'h006A; B = 16'h0030; #100;
A = 16'h006A; B = 16'h0031; #100;
A = 16'h006A; B = 16'h0032; #100;
A = 16'h006A; B = 16'h0033; #100;
A = 16'h006A; B = 16'h0034; #100;
A = 16'h006A; B = 16'h0035; #100;
A = 16'h006A; B = 16'h0036; #100;
A = 16'h006A; B = 16'h0037; #100;
A = 16'h006A; B = 16'h0038; #100;
A = 16'h006A; B = 16'h0039; #100;
A = 16'h006A; B = 16'h003A; #100;
A = 16'h006A; B = 16'h003B; #100;
A = 16'h006A; B = 16'h003C; #100;
A = 16'h006A; B = 16'h003D; #100;
A = 16'h006A; B = 16'h003E; #100;
A = 16'h006A; B = 16'h003F; #100;
A = 16'h006A; B = 16'h0040; #100;
A = 16'h006A; B = 16'h0041; #100;
A = 16'h006A; B = 16'h0042; #100;
A = 16'h006A; B = 16'h0043; #100;
A = 16'h006A; B = 16'h0044; #100;
A = 16'h006A; B = 16'h0045; #100;
A = 16'h006A; B = 16'h0046; #100;
A = 16'h006A; B = 16'h0047; #100;
A = 16'h006A; B = 16'h0048; #100;
A = 16'h006A; B = 16'h0049; #100;
A = 16'h006A; B = 16'h004A; #100;
A = 16'h006A; B = 16'h004B; #100;
A = 16'h006A; B = 16'h004C; #100;
A = 16'h006A; B = 16'h004D; #100;
A = 16'h006A; B = 16'h004E; #100;
A = 16'h006A; B = 16'h004F; #100;
A = 16'h006A; B = 16'h0050; #100;
A = 16'h006A; B = 16'h0051; #100;
A = 16'h006A; B = 16'h0052; #100;
A = 16'h006A; B = 16'h0053; #100;
A = 16'h006A; B = 16'h0054; #100;
A = 16'h006A; B = 16'h0055; #100;
A = 16'h006A; B = 16'h0056; #100;
A = 16'h006A; B = 16'h0057; #100;
A = 16'h006A; B = 16'h0058; #100;
A = 16'h006A; B = 16'h0059; #100;
A = 16'h006A; B = 16'h005A; #100;
A = 16'h006A; B = 16'h005B; #100;
A = 16'h006A; B = 16'h005C; #100;
A = 16'h006A; B = 16'h005D; #100;
A = 16'h006A; B = 16'h005E; #100;
A = 16'h006A; B = 16'h005F; #100;
A = 16'h006A; B = 16'h0060; #100;
A = 16'h006A; B = 16'h0061; #100;
A = 16'h006A; B = 16'h0062; #100;
A = 16'h006A; B = 16'h0063; #100;
A = 16'h006A; B = 16'h0064; #100;
A = 16'h006A; B = 16'h0065; #100;
A = 16'h006A; B = 16'h0066; #100;
A = 16'h006A; B = 16'h0067; #100;
A = 16'h006A; B = 16'h0068; #100;
A = 16'h006A; B = 16'h0069; #100;
A = 16'h006A; B = 16'h006A; #100;
A = 16'h006A; B = 16'h006B; #100;
A = 16'h006A; B = 16'h006C; #100;
A = 16'h006A; B = 16'h006D; #100;
A = 16'h006A; B = 16'h006E; #100;
A = 16'h006A; B = 16'h006F; #100;
A = 16'h006A; B = 16'h0070; #100;
A = 16'h006A; B = 16'h0071; #100;
A = 16'h006A; B = 16'h0072; #100;
A = 16'h006A; B = 16'h0073; #100;
A = 16'h006A; B = 16'h0074; #100;
A = 16'h006A; B = 16'h0075; #100;
A = 16'h006A; B = 16'h0076; #100;
A = 16'h006A; B = 16'h0077; #100;
A = 16'h006A; B = 16'h0078; #100;
A = 16'h006A; B = 16'h0079; #100;
A = 16'h006A; B = 16'h007A; #100;
A = 16'h006A; B = 16'h007B; #100;
A = 16'h006A; B = 16'h007C; #100;
A = 16'h006A; B = 16'h007D; #100;
A = 16'h006A; B = 16'h007E; #100;
A = 16'h006A; B = 16'h007F; #100;
A = 16'h006A; B = 16'h0080; #100;
A = 16'h006A; B = 16'h0081; #100;
A = 16'h006A; B = 16'h0082; #100;
A = 16'h006A; B = 16'h0083; #100;
A = 16'h006A; B = 16'h0084; #100;
A = 16'h006A; B = 16'h0085; #100;
A = 16'h006A; B = 16'h0086; #100;
A = 16'h006A; B = 16'h0087; #100;
A = 16'h006A; B = 16'h0088; #100;
A = 16'h006A; B = 16'h0089; #100;
A = 16'h006A; B = 16'h008A; #100;
A = 16'h006A; B = 16'h008B; #100;
A = 16'h006A; B = 16'h008C; #100;
A = 16'h006A; B = 16'h008D; #100;
A = 16'h006A; B = 16'h008E; #100;
A = 16'h006A; B = 16'h008F; #100;
A = 16'h006A; B = 16'h0090; #100;
A = 16'h006A; B = 16'h0091; #100;
A = 16'h006A; B = 16'h0092; #100;
A = 16'h006A; B = 16'h0093; #100;
A = 16'h006A; B = 16'h0094; #100;
A = 16'h006A; B = 16'h0095; #100;
A = 16'h006A; B = 16'h0096; #100;
A = 16'h006A; B = 16'h0097; #100;
A = 16'h006A; B = 16'h0098; #100;
A = 16'h006A; B = 16'h0099; #100;
A = 16'h006A; B = 16'h009A; #100;
A = 16'h006A; B = 16'h009B; #100;
A = 16'h006A; B = 16'h009C; #100;
A = 16'h006A; B = 16'h009D; #100;
A = 16'h006A; B = 16'h009E; #100;
A = 16'h006A; B = 16'h009F; #100;
A = 16'h006A; B = 16'h00A0; #100;
A = 16'h006A; B = 16'h00A1; #100;
A = 16'h006A; B = 16'h00A2; #100;
A = 16'h006A; B = 16'h00A3; #100;
A = 16'h006A; B = 16'h00A4; #100;
A = 16'h006A; B = 16'h00A5; #100;
A = 16'h006A; B = 16'h00A6; #100;
A = 16'h006A; B = 16'h00A7; #100;
A = 16'h006A; B = 16'h00A8; #100;
A = 16'h006A; B = 16'h00A9; #100;
A = 16'h006A; B = 16'h00AA; #100;
A = 16'h006A; B = 16'h00AB; #100;
A = 16'h006A; B = 16'h00AC; #100;
A = 16'h006A; B = 16'h00AD; #100;
A = 16'h006A; B = 16'h00AE; #100;
A = 16'h006A; B = 16'h00AF; #100;
A = 16'h006A; B = 16'h00B0; #100;
A = 16'h006A; B = 16'h00B1; #100;
A = 16'h006A; B = 16'h00B2; #100;
A = 16'h006A; B = 16'h00B3; #100;
A = 16'h006A; B = 16'h00B4; #100;
A = 16'h006A; B = 16'h00B5; #100;
A = 16'h006A; B = 16'h00B6; #100;
A = 16'h006A; B = 16'h00B7; #100;
A = 16'h006A; B = 16'h00B8; #100;
A = 16'h006A; B = 16'h00B9; #100;
A = 16'h006A; B = 16'h00BA; #100;
A = 16'h006A; B = 16'h00BB; #100;
A = 16'h006A; B = 16'h00BC; #100;
A = 16'h006A; B = 16'h00BD; #100;
A = 16'h006A; B = 16'h00BE; #100;
A = 16'h006A; B = 16'h00BF; #100;
A = 16'h006A; B = 16'h00C0; #100;
A = 16'h006A; B = 16'h00C1; #100;
A = 16'h006A; B = 16'h00C2; #100;
A = 16'h006A; B = 16'h00C3; #100;
A = 16'h006A; B = 16'h00C4; #100;
A = 16'h006A; B = 16'h00C5; #100;
A = 16'h006A; B = 16'h00C6; #100;
A = 16'h006A; B = 16'h00C7; #100;
A = 16'h006A; B = 16'h00C8; #100;
A = 16'h006A; B = 16'h00C9; #100;
A = 16'h006A; B = 16'h00CA; #100;
A = 16'h006A; B = 16'h00CB; #100;
A = 16'h006A; B = 16'h00CC; #100;
A = 16'h006A; B = 16'h00CD; #100;
A = 16'h006A; B = 16'h00CE; #100;
A = 16'h006A; B = 16'h00CF; #100;
A = 16'h006A; B = 16'h00D0; #100;
A = 16'h006A; B = 16'h00D1; #100;
A = 16'h006A; B = 16'h00D2; #100;
A = 16'h006A; B = 16'h00D3; #100;
A = 16'h006A; B = 16'h00D4; #100;
A = 16'h006A; B = 16'h00D5; #100;
A = 16'h006A; B = 16'h00D6; #100;
A = 16'h006A; B = 16'h00D7; #100;
A = 16'h006A; B = 16'h00D8; #100;
A = 16'h006A; B = 16'h00D9; #100;
A = 16'h006A; B = 16'h00DA; #100;
A = 16'h006A; B = 16'h00DB; #100;
A = 16'h006A; B = 16'h00DC; #100;
A = 16'h006A; B = 16'h00DD; #100;
A = 16'h006A; B = 16'h00DE; #100;
A = 16'h006A; B = 16'h00DF; #100;
A = 16'h006A; B = 16'h00E0; #100;
A = 16'h006A; B = 16'h00E1; #100;
A = 16'h006A; B = 16'h00E2; #100;
A = 16'h006A; B = 16'h00E3; #100;
A = 16'h006A; B = 16'h00E4; #100;
A = 16'h006A; B = 16'h00E5; #100;
A = 16'h006A; B = 16'h00E6; #100;
A = 16'h006A; B = 16'h00E7; #100;
A = 16'h006A; B = 16'h00E8; #100;
A = 16'h006A; B = 16'h00E9; #100;
A = 16'h006A; B = 16'h00EA; #100;
A = 16'h006A; B = 16'h00EB; #100;
A = 16'h006A; B = 16'h00EC; #100;
A = 16'h006A; B = 16'h00ED; #100;
A = 16'h006A; B = 16'h00EE; #100;
A = 16'h006A; B = 16'h00EF; #100;
A = 16'h006A; B = 16'h00F0; #100;
A = 16'h006A; B = 16'h00F1; #100;
A = 16'h006A; B = 16'h00F2; #100;
A = 16'h006A; B = 16'h00F3; #100;
A = 16'h006A; B = 16'h00F4; #100;
A = 16'h006A; B = 16'h00F5; #100;
A = 16'h006A; B = 16'h00F6; #100;
A = 16'h006A; B = 16'h00F7; #100;
A = 16'h006A; B = 16'h00F8; #100;
A = 16'h006A; B = 16'h00F9; #100;
A = 16'h006A; B = 16'h00FA; #100;
A = 16'h006A; B = 16'h00FB; #100;
A = 16'h006A; B = 16'h00FC; #100;
A = 16'h006A; B = 16'h00FD; #100;
A = 16'h006A; B = 16'h00FE; #100;
A = 16'h006A; B = 16'h00FF; #100;
A = 16'h006B; B = 16'h000; #100;
A = 16'h006B; B = 16'h001; #100;
A = 16'h006B; B = 16'h002; #100;
A = 16'h006B; B = 16'h003; #100;
A = 16'h006B; B = 16'h004; #100;
A = 16'h006B; B = 16'h005; #100;
A = 16'h006B; B = 16'h006; #100;
A = 16'h006B; B = 16'h007; #100;
A = 16'h006B; B = 16'h008; #100;
A = 16'h006B; B = 16'h009; #100;
A = 16'h006B; B = 16'h00A; #100;
A = 16'h006B; B = 16'h00B; #100;
A = 16'h006B; B = 16'h00C; #100;
A = 16'h006B; B = 16'h00D; #100;
A = 16'h006B; B = 16'h00E; #100;
A = 16'h006B; B = 16'h00F; #100;
A = 16'h006B; B = 16'h0010; #100;
A = 16'h006B; B = 16'h0011; #100;
A = 16'h006B; B = 16'h0012; #100;
A = 16'h006B; B = 16'h0013; #100;
A = 16'h006B; B = 16'h0014; #100;
A = 16'h006B; B = 16'h0015; #100;
A = 16'h006B; B = 16'h0016; #100;
A = 16'h006B; B = 16'h0017; #100;
A = 16'h006B; B = 16'h0018; #100;
A = 16'h006B; B = 16'h0019; #100;
A = 16'h006B; B = 16'h001A; #100;
A = 16'h006B; B = 16'h001B; #100;
A = 16'h006B; B = 16'h001C; #100;
A = 16'h006B; B = 16'h001D; #100;
A = 16'h006B; B = 16'h001E; #100;
A = 16'h006B; B = 16'h001F; #100;
A = 16'h006B; B = 16'h0020; #100;
A = 16'h006B; B = 16'h0021; #100;
A = 16'h006B; B = 16'h0022; #100;
A = 16'h006B; B = 16'h0023; #100;
A = 16'h006B; B = 16'h0024; #100;
A = 16'h006B; B = 16'h0025; #100;
A = 16'h006B; B = 16'h0026; #100;
A = 16'h006B; B = 16'h0027; #100;
A = 16'h006B; B = 16'h0028; #100;
A = 16'h006B; B = 16'h0029; #100;
A = 16'h006B; B = 16'h002A; #100;
A = 16'h006B; B = 16'h002B; #100;
A = 16'h006B; B = 16'h002C; #100;
A = 16'h006B; B = 16'h002D; #100;
A = 16'h006B; B = 16'h002E; #100;
A = 16'h006B; B = 16'h002F; #100;
A = 16'h006B; B = 16'h0030; #100;
A = 16'h006B; B = 16'h0031; #100;
A = 16'h006B; B = 16'h0032; #100;
A = 16'h006B; B = 16'h0033; #100;
A = 16'h006B; B = 16'h0034; #100;
A = 16'h006B; B = 16'h0035; #100;
A = 16'h006B; B = 16'h0036; #100;
A = 16'h006B; B = 16'h0037; #100;
A = 16'h006B; B = 16'h0038; #100;
A = 16'h006B; B = 16'h0039; #100;
A = 16'h006B; B = 16'h003A; #100;
A = 16'h006B; B = 16'h003B; #100;
A = 16'h006B; B = 16'h003C; #100;
A = 16'h006B; B = 16'h003D; #100;
A = 16'h006B; B = 16'h003E; #100;
A = 16'h006B; B = 16'h003F; #100;
A = 16'h006B; B = 16'h0040; #100;
A = 16'h006B; B = 16'h0041; #100;
A = 16'h006B; B = 16'h0042; #100;
A = 16'h006B; B = 16'h0043; #100;
A = 16'h006B; B = 16'h0044; #100;
A = 16'h006B; B = 16'h0045; #100;
A = 16'h006B; B = 16'h0046; #100;
A = 16'h006B; B = 16'h0047; #100;
A = 16'h006B; B = 16'h0048; #100;
A = 16'h006B; B = 16'h0049; #100;
A = 16'h006B; B = 16'h004A; #100;
A = 16'h006B; B = 16'h004B; #100;
A = 16'h006B; B = 16'h004C; #100;
A = 16'h006B; B = 16'h004D; #100;
A = 16'h006B; B = 16'h004E; #100;
A = 16'h006B; B = 16'h004F; #100;
A = 16'h006B; B = 16'h0050; #100;
A = 16'h006B; B = 16'h0051; #100;
A = 16'h006B; B = 16'h0052; #100;
A = 16'h006B; B = 16'h0053; #100;
A = 16'h006B; B = 16'h0054; #100;
A = 16'h006B; B = 16'h0055; #100;
A = 16'h006B; B = 16'h0056; #100;
A = 16'h006B; B = 16'h0057; #100;
A = 16'h006B; B = 16'h0058; #100;
A = 16'h006B; B = 16'h0059; #100;
A = 16'h006B; B = 16'h005A; #100;
A = 16'h006B; B = 16'h005B; #100;
A = 16'h006B; B = 16'h005C; #100;
A = 16'h006B; B = 16'h005D; #100;
A = 16'h006B; B = 16'h005E; #100;
A = 16'h006B; B = 16'h005F; #100;
A = 16'h006B; B = 16'h0060; #100;
A = 16'h006B; B = 16'h0061; #100;
A = 16'h006B; B = 16'h0062; #100;
A = 16'h006B; B = 16'h0063; #100;
A = 16'h006B; B = 16'h0064; #100;
A = 16'h006B; B = 16'h0065; #100;
A = 16'h006B; B = 16'h0066; #100;
A = 16'h006B; B = 16'h0067; #100;
A = 16'h006B; B = 16'h0068; #100;
A = 16'h006B; B = 16'h0069; #100;
A = 16'h006B; B = 16'h006A; #100;
A = 16'h006B; B = 16'h006B; #100;
A = 16'h006B; B = 16'h006C; #100;
A = 16'h006B; B = 16'h006D; #100;
A = 16'h006B; B = 16'h006E; #100;
A = 16'h006B; B = 16'h006F; #100;
A = 16'h006B; B = 16'h0070; #100;
A = 16'h006B; B = 16'h0071; #100;
A = 16'h006B; B = 16'h0072; #100;
A = 16'h006B; B = 16'h0073; #100;
A = 16'h006B; B = 16'h0074; #100;
A = 16'h006B; B = 16'h0075; #100;
A = 16'h006B; B = 16'h0076; #100;
A = 16'h006B; B = 16'h0077; #100;
A = 16'h006B; B = 16'h0078; #100;
A = 16'h006B; B = 16'h0079; #100;
A = 16'h006B; B = 16'h007A; #100;
A = 16'h006B; B = 16'h007B; #100;
A = 16'h006B; B = 16'h007C; #100;
A = 16'h006B; B = 16'h007D; #100;
A = 16'h006B; B = 16'h007E; #100;
A = 16'h006B; B = 16'h007F; #100;
A = 16'h006B; B = 16'h0080; #100;
A = 16'h006B; B = 16'h0081; #100;
A = 16'h006B; B = 16'h0082; #100;
A = 16'h006B; B = 16'h0083; #100;
A = 16'h006B; B = 16'h0084; #100;
A = 16'h006B; B = 16'h0085; #100;
A = 16'h006B; B = 16'h0086; #100;
A = 16'h006B; B = 16'h0087; #100;
A = 16'h006B; B = 16'h0088; #100;
A = 16'h006B; B = 16'h0089; #100;
A = 16'h006B; B = 16'h008A; #100;
A = 16'h006B; B = 16'h008B; #100;
A = 16'h006B; B = 16'h008C; #100;
A = 16'h006B; B = 16'h008D; #100;
A = 16'h006B; B = 16'h008E; #100;
A = 16'h006B; B = 16'h008F; #100;
A = 16'h006B; B = 16'h0090; #100;
A = 16'h006B; B = 16'h0091; #100;
A = 16'h006B; B = 16'h0092; #100;
A = 16'h006B; B = 16'h0093; #100;
A = 16'h006B; B = 16'h0094; #100;
A = 16'h006B; B = 16'h0095; #100;
A = 16'h006B; B = 16'h0096; #100;
A = 16'h006B; B = 16'h0097; #100;
A = 16'h006B; B = 16'h0098; #100;
A = 16'h006B; B = 16'h0099; #100;
A = 16'h006B; B = 16'h009A; #100;
A = 16'h006B; B = 16'h009B; #100;
A = 16'h006B; B = 16'h009C; #100;
A = 16'h006B; B = 16'h009D; #100;
A = 16'h006B; B = 16'h009E; #100;
A = 16'h006B; B = 16'h009F; #100;
A = 16'h006B; B = 16'h00A0; #100;
A = 16'h006B; B = 16'h00A1; #100;
A = 16'h006B; B = 16'h00A2; #100;
A = 16'h006B; B = 16'h00A3; #100;
A = 16'h006B; B = 16'h00A4; #100;
A = 16'h006B; B = 16'h00A5; #100;
A = 16'h006B; B = 16'h00A6; #100;
A = 16'h006B; B = 16'h00A7; #100;
A = 16'h006B; B = 16'h00A8; #100;
A = 16'h006B; B = 16'h00A9; #100;
A = 16'h006B; B = 16'h00AA; #100;
A = 16'h006B; B = 16'h00AB; #100;
A = 16'h006B; B = 16'h00AC; #100;
A = 16'h006B; B = 16'h00AD; #100;
A = 16'h006B; B = 16'h00AE; #100;
A = 16'h006B; B = 16'h00AF; #100;
A = 16'h006B; B = 16'h00B0; #100;
A = 16'h006B; B = 16'h00B1; #100;
A = 16'h006B; B = 16'h00B2; #100;
A = 16'h006B; B = 16'h00B3; #100;
A = 16'h006B; B = 16'h00B4; #100;
A = 16'h006B; B = 16'h00B5; #100;
A = 16'h006B; B = 16'h00B6; #100;
A = 16'h006B; B = 16'h00B7; #100;
A = 16'h006B; B = 16'h00B8; #100;
A = 16'h006B; B = 16'h00B9; #100;
A = 16'h006B; B = 16'h00BA; #100;
A = 16'h006B; B = 16'h00BB; #100;
A = 16'h006B; B = 16'h00BC; #100;
A = 16'h006B; B = 16'h00BD; #100;
A = 16'h006B; B = 16'h00BE; #100;
A = 16'h006B; B = 16'h00BF; #100;
A = 16'h006B; B = 16'h00C0; #100;
A = 16'h006B; B = 16'h00C1; #100;
A = 16'h006B; B = 16'h00C2; #100;
A = 16'h006B; B = 16'h00C3; #100;
A = 16'h006B; B = 16'h00C4; #100;
A = 16'h006B; B = 16'h00C5; #100;
A = 16'h006B; B = 16'h00C6; #100;
A = 16'h006B; B = 16'h00C7; #100;
A = 16'h006B; B = 16'h00C8; #100;
A = 16'h006B; B = 16'h00C9; #100;
A = 16'h006B; B = 16'h00CA; #100;
A = 16'h006B; B = 16'h00CB; #100;
A = 16'h006B; B = 16'h00CC; #100;
A = 16'h006B; B = 16'h00CD; #100;
A = 16'h006B; B = 16'h00CE; #100;
A = 16'h006B; B = 16'h00CF; #100;
A = 16'h006B; B = 16'h00D0; #100;
A = 16'h006B; B = 16'h00D1; #100;
A = 16'h006B; B = 16'h00D2; #100;
A = 16'h006B; B = 16'h00D3; #100;
A = 16'h006B; B = 16'h00D4; #100;
A = 16'h006B; B = 16'h00D5; #100;
A = 16'h006B; B = 16'h00D6; #100;
A = 16'h006B; B = 16'h00D7; #100;
A = 16'h006B; B = 16'h00D8; #100;
A = 16'h006B; B = 16'h00D9; #100;
A = 16'h006B; B = 16'h00DA; #100;
A = 16'h006B; B = 16'h00DB; #100;
A = 16'h006B; B = 16'h00DC; #100;
A = 16'h006B; B = 16'h00DD; #100;
A = 16'h006B; B = 16'h00DE; #100;
A = 16'h006B; B = 16'h00DF; #100;
A = 16'h006B; B = 16'h00E0; #100;
A = 16'h006B; B = 16'h00E1; #100;
A = 16'h006B; B = 16'h00E2; #100;
A = 16'h006B; B = 16'h00E3; #100;
A = 16'h006B; B = 16'h00E4; #100;
A = 16'h006B; B = 16'h00E5; #100;
A = 16'h006B; B = 16'h00E6; #100;
A = 16'h006B; B = 16'h00E7; #100;
A = 16'h006B; B = 16'h00E8; #100;
A = 16'h006B; B = 16'h00E9; #100;
A = 16'h006B; B = 16'h00EA; #100;
A = 16'h006B; B = 16'h00EB; #100;
A = 16'h006B; B = 16'h00EC; #100;
A = 16'h006B; B = 16'h00ED; #100;
A = 16'h006B; B = 16'h00EE; #100;
A = 16'h006B; B = 16'h00EF; #100;
A = 16'h006B; B = 16'h00F0; #100;
A = 16'h006B; B = 16'h00F1; #100;
A = 16'h006B; B = 16'h00F2; #100;
A = 16'h006B; B = 16'h00F3; #100;
A = 16'h006B; B = 16'h00F4; #100;
A = 16'h006B; B = 16'h00F5; #100;
A = 16'h006B; B = 16'h00F6; #100;
A = 16'h006B; B = 16'h00F7; #100;
A = 16'h006B; B = 16'h00F8; #100;
A = 16'h006B; B = 16'h00F9; #100;
A = 16'h006B; B = 16'h00FA; #100;
A = 16'h006B; B = 16'h00FB; #100;
A = 16'h006B; B = 16'h00FC; #100;
A = 16'h006B; B = 16'h00FD; #100;
A = 16'h006B; B = 16'h00FE; #100;
A = 16'h006B; B = 16'h00FF; #100;
A = 16'h006C; B = 16'h000; #100;
A = 16'h006C; B = 16'h001; #100;
A = 16'h006C; B = 16'h002; #100;
A = 16'h006C; B = 16'h003; #100;
A = 16'h006C; B = 16'h004; #100;
A = 16'h006C; B = 16'h005; #100;
A = 16'h006C; B = 16'h006; #100;
A = 16'h006C; B = 16'h007; #100;
A = 16'h006C; B = 16'h008; #100;
A = 16'h006C; B = 16'h009; #100;
A = 16'h006C; B = 16'h00A; #100;
A = 16'h006C; B = 16'h00B; #100;
A = 16'h006C; B = 16'h00C; #100;
A = 16'h006C; B = 16'h00D; #100;
A = 16'h006C; B = 16'h00E; #100;
A = 16'h006C; B = 16'h00F; #100;
A = 16'h006C; B = 16'h0010; #100;
A = 16'h006C; B = 16'h0011; #100;
A = 16'h006C; B = 16'h0012; #100;
A = 16'h006C; B = 16'h0013; #100;
A = 16'h006C; B = 16'h0014; #100;
A = 16'h006C; B = 16'h0015; #100;
A = 16'h006C; B = 16'h0016; #100;
A = 16'h006C; B = 16'h0017; #100;
A = 16'h006C; B = 16'h0018; #100;
A = 16'h006C; B = 16'h0019; #100;
A = 16'h006C; B = 16'h001A; #100;
A = 16'h006C; B = 16'h001B; #100;
A = 16'h006C; B = 16'h001C; #100;
A = 16'h006C; B = 16'h001D; #100;
A = 16'h006C; B = 16'h001E; #100;
A = 16'h006C; B = 16'h001F; #100;
A = 16'h006C; B = 16'h0020; #100;
A = 16'h006C; B = 16'h0021; #100;
A = 16'h006C; B = 16'h0022; #100;
A = 16'h006C; B = 16'h0023; #100;
A = 16'h006C; B = 16'h0024; #100;
A = 16'h006C; B = 16'h0025; #100;
A = 16'h006C; B = 16'h0026; #100;
A = 16'h006C; B = 16'h0027; #100;
A = 16'h006C; B = 16'h0028; #100;
A = 16'h006C; B = 16'h0029; #100;
A = 16'h006C; B = 16'h002A; #100;
A = 16'h006C; B = 16'h002B; #100;
A = 16'h006C; B = 16'h002C; #100;
A = 16'h006C; B = 16'h002D; #100;
A = 16'h006C; B = 16'h002E; #100;
A = 16'h006C; B = 16'h002F; #100;
A = 16'h006C; B = 16'h0030; #100;
A = 16'h006C; B = 16'h0031; #100;
A = 16'h006C; B = 16'h0032; #100;
A = 16'h006C; B = 16'h0033; #100;
A = 16'h006C; B = 16'h0034; #100;
A = 16'h006C; B = 16'h0035; #100;
A = 16'h006C; B = 16'h0036; #100;
A = 16'h006C; B = 16'h0037; #100;
A = 16'h006C; B = 16'h0038; #100;
A = 16'h006C; B = 16'h0039; #100;
A = 16'h006C; B = 16'h003A; #100;
A = 16'h006C; B = 16'h003B; #100;
A = 16'h006C; B = 16'h003C; #100;
A = 16'h006C; B = 16'h003D; #100;
A = 16'h006C; B = 16'h003E; #100;
A = 16'h006C; B = 16'h003F; #100;
A = 16'h006C; B = 16'h0040; #100;
A = 16'h006C; B = 16'h0041; #100;
A = 16'h006C; B = 16'h0042; #100;
A = 16'h006C; B = 16'h0043; #100;
A = 16'h006C; B = 16'h0044; #100;
A = 16'h006C; B = 16'h0045; #100;
A = 16'h006C; B = 16'h0046; #100;
A = 16'h006C; B = 16'h0047; #100;
A = 16'h006C; B = 16'h0048; #100;
A = 16'h006C; B = 16'h0049; #100;
A = 16'h006C; B = 16'h004A; #100;
A = 16'h006C; B = 16'h004B; #100;
A = 16'h006C; B = 16'h004C; #100;
A = 16'h006C; B = 16'h004D; #100;
A = 16'h006C; B = 16'h004E; #100;
A = 16'h006C; B = 16'h004F; #100;
A = 16'h006C; B = 16'h0050; #100;
A = 16'h006C; B = 16'h0051; #100;
A = 16'h006C; B = 16'h0052; #100;
A = 16'h006C; B = 16'h0053; #100;
A = 16'h006C; B = 16'h0054; #100;
A = 16'h006C; B = 16'h0055; #100;
A = 16'h006C; B = 16'h0056; #100;
A = 16'h006C; B = 16'h0057; #100;
A = 16'h006C; B = 16'h0058; #100;
A = 16'h006C; B = 16'h0059; #100;
A = 16'h006C; B = 16'h005A; #100;
A = 16'h006C; B = 16'h005B; #100;
A = 16'h006C; B = 16'h005C; #100;
A = 16'h006C; B = 16'h005D; #100;
A = 16'h006C; B = 16'h005E; #100;
A = 16'h006C; B = 16'h005F; #100;
A = 16'h006C; B = 16'h0060; #100;
A = 16'h006C; B = 16'h0061; #100;
A = 16'h006C; B = 16'h0062; #100;
A = 16'h006C; B = 16'h0063; #100;
A = 16'h006C; B = 16'h0064; #100;
A = 16'h006C; B = 16'h0065; #100;
A = 16'h006C; B = 16'h0066; #100;
A = 16'h006C; B = 16'h0067; #100;
A = 16'h006C; B = 16'h0068; #100;
A = 16'h006C; B = 16'h0069; #100;
A = 16'h006C; B = 16'h006A; #100;
A = 16'h006C; B = 16'h006B; #100;
A = 16'h006C; B = 16'h006C; #100;
A = 16'h006C; B = 16'h006D; #100;
A = 16'h006C; B = 16'h006E; #100;
A = 16'h006C; B = 16'h006F; #100;
A = 16'h006C; B = 16'h0070; #100;
A = 16'h006C; B = 16'h0071; #100;
A = 16'h006C; B = 16'h0072; #100;
A = 16'h006C; B = 16'h0073; #100;
A = 16'h006C; B = 16'h0074; #100;
A = 16'h006C; B = 16'h0075; #100;
A = 16'h006C; B = 16'h0076; #100;
A = 16'h006C; B = 16'h0077; #100;
A = 16'h006C; B = 16'h0078; #100;
A = 16'h006C; B = 16'h0079; #100;
A = 16'h006C; B = 16'h007A; #100;
A = 16'h006C; B = 16'h007B; #100;
A = 16'h006C; B = 16'h007C; #100;
A = 16'h006C; B = 16'h007D; #100;
A = 16'h006C; B = 16'h007E; #100;
A = 16'h006C; B = 16'h007F; #100;
A = 16'h006C; B = 16'h0080; #100;
A = 16'h006C; B = 16'h0081; #100;
A = 16'h006C; B = 16'h0082; #100;
A = 16'h006C; B = 16'h0083; #100;
A = 16'h006C; B = 16'h0084; #100;
A = 16'h006C; B = 16'h0085; #100;
A = 16'h006C; B = 16'h0086; #100;
A = 16'h006C; B = 16'h0087; #100;
A = 16'h006C; B = 16'h0088; #100;
A = 16'h006C; B = 16'h0089; #100;
A = 16'h006C; B = 16'h008A; #100;
A = 16'h006C; B = 16'h008B; #100;
A = 16'h006C; B = 16'h008C; #100;
A = 16'h006C; B = 16'h008D; #100;
A = 16'h006C; B = 16'h008E; #100;
A = 16'h006C; B = 16'h008F; #100;
A = 16'h006C; B = 16'h0090; #100;
A = 16'h006C; B = 16'h0091; #100;
A = 16'h006C; B = 16'h0092; #100;
A = 16'h006C; B = 16'h0093; #100;
A = 16'h006C; B = 16'h0094; #100;
A = 16'h006C; B = 16'h0095; #100;
A = 16'h006C; B = 16'h0096; #100;
A = 16'h006C; B = 16'h0097; #100;
A = 16'h006C; B = 16'h0098; #100;
A = 16'h006C; B = 16'h0099; #100;
A = 16'h006C; B = 16'h009A; #100;
A = 16'h006C; B = 16'h009B; #100;
A = 16'h006C; B = 16'h009C; #100;
A = 16'h006C; B = 16'h009D; #100;
A = 16'h006C; B = 16'h009E; #100;
A = 16'h006C; B = 16'h009F; #100;
A = 16'h006C; B = 16'h00A0; #100;
A = 16'h006C; B = 16'h00A1; #100;
A = 16'h006C; B = 16'h00A2; #100;
A = 16'h006C; B = 16'h00A3; #100;
A = 16'h006C; B = 16'h00A4; #100;
A = 16'h006C; B = 16'h00A5; #100;
A = 16'h006C; B = 16'h00A6; #100;
A = 16'h006C; B = 16'h00A7; #100;
A = 16'h006C; B = 16'h00A8; #100;
A = 16'h006C; B = 16'h00A9; #100;
A = 16'h006C; B = 16'h00AA; #100;
A = 16'h006C; B = 16'h00AB; #100;
A = 16'h006C; B = 16'h00AC; #100;
A = 16'h006C; B = 16'h00AD; #100;
A = 16'h006C; B = 16'h00AE; #100;
A = 16'h006C; B = 16'h00AF; #100;
A = 16'h006C; B = 16'h00B0; #100;
A = 16'h006C; B = 16'h00B1; #100;
A = 16'h006C; B = 16'h00B2; #100;
A = 16'h006C; B = 16'h00B3; #100;
A = 16'h006C; B = 16'h00B4; #100;
A = 16'h006C; B = 16'h00B5; #100;
A = 16'h006C; B = 16'h00B6; #100;
A = 16'h006C; B = 16'h00B7; #100;
A = 16'h006C; B = 16'h00B8; #100;
A = 16'h006C; B = 16'h00B9; #100;
A = 16'h006C; B = 16'h00BA; #100;
A = 16'h006C; B = 16'h00BB; #100;
A = 16'h006C; B = 16'h00BC; #100;
A = 16'h006C; B = 16'h00BD; #100;
A = 16'h006C; B = 16'h00BE; #100;
A = 16'h006C; B = 16'h00BF; #100;
A = 16'h006C; B = 16'h00C0; #100;
A = 16'h006C; B = 16'h00C1; #100;
A = 16'h006C; B = 16'h00C2; #100;
A = 16'h006C; B = 16'h00C3; #100;
A = 16'h006C; B = 16'h00C4; #100;
A = 16'h006C; B = 16'h00C5; #100;
A = 16'h006C; B = 16'h00C6; #100;
A = 16'h006C; B = 16'h00C7; #100;
A = 16'h006C; B = 16'h00C8; #100;
A = 16'h006C; B = 16'h00C9; #100;
A = 16'h006C; B = 16'h00CA; #100;
A = 16'h006C; B = 16'h00CB; #100;
A = 16'h006C; B = 16'h00CC; #100;
A = 16'h006C; B = 16'h00CD; #100;
A = 16'h006C; B = 16'h00CE; #100;
A = 16'h006C; B = 16'h00CF; #100;
A = 16'h006C; B = 16'h00D0; #100;
A = 16'h006C; B = 16'h00D1; #100;
A = 16'h006C; B = 16'h00D2; #100;
A = 16'h006C; B = 16'h00D3; #100;
A = 16'h006C; B = 16'h00D4; #100;
A = 16'h006C; B = 16'h00D5; #100;
A = 16'h006C; B = 16'h00D6; #100;
A = 16'h006C; B = 16'h00D7; #100;
A = 16'h006C; B = 16'h00D8; #100;
A = 16'h006C; B = 16'h00D9; #100;
A = 16'h006C; B = 16'h00DA; #100;
A = 16'h006C; B = 16'h00DB; #100;
A = 16'h006C; B = 16'h00DC; #100;
A = 16'h006C; B = 16'h00DD; #100;
A = 16'h006C; B = 16'h00DE; #100;
A = 16'h006C; B = 16'h00DF; #100;
A = 16'h006C; B = 16'h00E0; #100;
A = 16'h006C; B = 16'h00E1; #100;
A = 16'h006C; B = 16'h00E2; #100;
A = 16'h006C; B = 16'h00E3; #100;
A = 16'h006C; B = 16'h00E4; #100;
A = 16'h006C; B = 16'h00E5; #100;
A = 16'h006C; B = 16'h00E6; #100;
A = 16'h006C; B = 16'h00E7; #100;
A = 16'h006C; B = 16'h00E8; #100;
A = 16'h006C; B = 16'h00E9; #100;
A = 16'h006C; B = 16'h00EA; #100;
A = 16'h006C; B = 16'h00EB; #100;
A = 16'h006C; B = 16'h00EC; #100;
A = 16'h006C; B = 16'h00ED; #100;
A = 16'h006C; B = 16'h00EE; #100;
A = 16'h006C; B = 16'h00EF; #100;
A = 16'h006C; B = 16'h00F0; #100;
A = 16'h006C; B = 16'h00F1; #100;
A = 16'h006C; B = 16'h00F2; #100;
A = 16'h006C; B = 16'h00F3; #100;
A = 16'h006C; B = 16'h00F4; #100;
A = 16'h006C; B = 16'h00F5; #100;
A = 16'h006C; B = 16'h00F6; #100;
A = 16'h006C; B = 16'h00F7; #100;
A = 16'h006C; B = 16'h00F8; #100;
A = 16'h006C; B = 16'h00F9; #100;
A = 16'h006C; B = 16'h00FA; #100;
A = 16'h006C; B = 16'h00FB; #100;
A = 16'h006C; B = 16'h00FC; #100;
A = 16'h006C; B = 16'h00FD; #100;
A = 16'h006C; B = 16'h00FE; #100;
A = 16'h006C; B = 16'h00FF; #100;
A = 16'h006D; B = 16'h000; #100;
A = 16'h006D; B = 16'h001; #100;
A = 16'h006D; B = 16'h002; #100;
A = 16'h006D; B = 16'h003; #100;
A = 16'h006D; B = 16'h004; #100;
A = 16'h006D; B = 16'h005; #100;
A = 16'h006D; B = 16'h006; #100;
A = 16'h006D; B = 16'h007; #100;
A = 16'h006D; B = 16'h008; #100;
A = 16'h006D; B = 16'h009; #100;
A = 16'h006D; B = 16'h00A; #100;
A = 16'h006D; B = 16'h00B; #100;
A = 16'h006D; B = 16'h00C; #100;
A = 16'h006D; B = 16'h00D; #100;
A = 16'h006D; B = 16'h00E; #100;
A = 16'h006D; B = 16'h00F; #100;
A = 16'h006D; B = 16'h0010; #100;
A = 16'h006D; B = 16'h0011; #100;
A = 16'h006D; B = 16'h0012; #100;
A = 16'h006D; B = 16'h0013; #100;
A = 16'h006D; B = 16'h0014; #100;
A = 16'h006D; B = 16'h0015; #100;
A = 16'h006D; B = 16'h0016; #100;
A = 16'h006D; B = 16'h0017; #100;
A = 16'h006D; B = 16'h0018; #100;
A = 16'h006D; B = 16'h0019; #100;
A = 16'h006D; B = 16'h001A; #100;
A = 16'h006D; B = 16'h001B; #100;
A = 16'h006D; B = 16'h001C; #100;
A = 16'h006D; B = 16'h001D; #100;
A = 16'h006D; B = 16'h001E; #100;
A = 16'h006D; B = 16'h001F; #100;
A = 16'h006D; B = 16'h0020; #100;
A = 16'h006D; B = 16'h0021; #100;
A = 16'h006D; B = 16'h0022; #100;
A = 16'h006D; B = 16'h0023; #100;
A = 16'h006D; B = 16'h0024; #100;
A = 16'h006D; B = 16'h0025; #100;
A = 16'h006D; B = 16'h0026; #100;
A = 16'h006D; B = 16'h0027; #100;
A = 16'h006D; B = 16'h0028; #100;
A = 16'h006D; B = 16'h0029; #100;
A = 16'h006D; B = 16'h002A; #100;
A = 16'h006D; B = 16'h002B; #100;
A = 16'h006D; B = 16'h002C; #100;
A = 16'h006D; B = 16'h002D; #100;
A = 16'h006D; B = 16'h002E; #100;
A = 16'h006D; B = 16'h002F; #100;
A = 16'h006D; B = 16'h0030; #100;
A = 16'h006D; B = 16'h0031; #100;
A = 16'h006D; B = 16'h0032; #100;
A = 16'h006D; B = 16'h0033; #100;
A = 16'h006D; B = 16'h0034; #100;
A = 16'h006D; B = 16'h0035; #100;
A = 16'h006D; B = 16'h0036; #100;
A = 16'h006D; B = 16'h0037; #100;
A = 16'h006D; B = 16'h0038; #100;
A = 16'h006D; B = 16'h0039; #100;
A = 16'h006D; B = 16'h003A; #100;
A = 16'h006D; B = 16'h003B; #100;
A = 16'h006D; B = 16'h003C; #100;
A = 16'h006D; B = 16'h003D; #100;
A = 16'h006D; B = 16'h003E; #100;
A = 16'h006D; B = 16'h003F; #100;
A = 16'h006D; B = 16'h0040; #100;
A = 16'h006D; B = 16'h0041; #100;
A = 16'h006D; B = 16'h0042; #100;
A = 16'h006D; B = 16'h0043; #100;
A = 16'h006D; B = 16'h0044; #100;
A = 16'h006D; B = 16'h0045; #100;
A = 16'h006D; B = 16'h0046; #100;
A = 16'h006D; B = 16'h0047; #100;
A = 16'h006D; B = 16'h0048; #100;
A = 16'h006D; B = 16'h0049; #100;
A = 16'h006D; B = 16'h004A; #100;
A = 16'h006D; B = 16'h004B; #100;
A = 16'h006D; B = 16'h004C; #100;
A = 16'h006D; B = 16'h004D; #100;
A = 16'h006D; B = 16'h004E; #100;
A = 16'h006D; B = 16'h004F; #100;
A = 16'h006D; B = 16'h0050; #100;
A = 16'h006D; B = 16'h0051; #100;
A = 16'h006D; B = 16'h0052; #100;
A = 16'h006D; B = 16'h0053; #100;
A = 16'h006D; B = 16'h0054; #100;
A = 16'h006D; B = 16'h0055; #100;
A = 16'h006D; B = 16'h0056; #100;
A = 16'h006D; B = 16'h0057; #100;
A = 16'h006D; B = 16'h0058; #100;
A = 16'h006D; B = 16'h0059; #100;
A = 16'h006D; B = 16'h005A; #100;
A = 16'h006D; B = 16'h005B; #100;
A = 16'h006D; B = 16'h005C; #100;
A = 16'h006D; B = 16'h005D; #100;
A = 16'h006D; B = 16'h005E; #100;
A = 16'h006D; B = 16'h005F; #100;
A = 16'h006D; B = 16'h0060; #100;
A = 16'h006D; B = 16'h0061; #100;
A = 16'h006D; B = 16'h0062; #100;
A = 16'h006D; B = 16'h0063; #100;
A = 16'h006D; B = 16'h0064; #100;
A = 16'h006D; B = 16'h0065; #100;
A = 16'h006D; B = 16'h0066; #100;
A = 16'h006D; B = 16'h0067; #100;
A = 16'h006D; B = 16'h0068; #100;
A = 16'h006D; B = 16'h0069; #100;
A = 16'h006D; B = 16'h006A; #100;
A = 16'h006D; B = 16'h006B; #100;
A = 16'h006D; B = 16'h006C; #100;
A = 16'h006D; B = 16'h006D; #100;
A = 16'h006D; B = 16'h006E; #100;
A = 16'h006D; B = 16'h006F; #100;
A = 16'h006D; B = 16'h0070; #100;
A = 16'h006D; B = 16'h0071; #100;
A = 16'h006D; B = 16'h0072; #100;
A = 16'h006D; B = 16'h0073; #100;
A = 16'h006D; B = 16'h0074; #100;
A = 16'h006D; B = 16'h0075; #100;
A = 16'h006D; B = 16'h0076; #100;
A = 16'h006D; B = 16'h0077; #100;
A = 16'h006D; B = 16'h0078; #100;
A = 16'h006D; B = 16'h0079; #100;
A = 16'h006D; B = 16'h007A; #100;
A = 16'h006D; B = 16'h007B; #100;
A = 16'h006D; B = 16'h007C; #100;
A = 16'h006D; B = 16'h007D; #100;
A = 16'h006D; B = 16'h007E; #100;
A = 16'h006D; B = 16'h007F; #100;
A = 16'h006D; B = 16'h0080; #100;
A = 16'h006D; B = 16'h0081; #100;
A = 16'h006D; B = 16'h0082; #100;
A = 16'h006D; B = 16'h0083; #100;
A = 16'h006D; B = 16'h0084; #100;
A = 16'h006D; B = 16'h0085; #100;
A = 16'h006D; B = 16'h0086; #100;
A = 16'h006D; B = 16'h0087; #100;
A = 16'h006D; B = 16'h0088; #100;
A = 16'h006D; B = 16'h0089; #100;
A = 16'h006D; B = 16'h008A; #100;
A = 16'h006D; B = 16'h008B; #100;
A = 16'h006D; B = 16'h008C; #100;
A = 16'h006D; B = 16'h008D; #100;
A = 16'h006D; B = 16'h008E; #100;
A = 16'h006D; B = 16'h008F; #100;
A = 16'h006D; B = 16'h0090; #100;
A = 16'h006D; B = 16'h0091; #100;
A = 16'h006D; B = 16'h0092; #100;
A = 16'h006D; B = 16'h0093; #100;
A = 16'h006D; B = 16'h0094; #100;
A = 16'h006D; B = 16'h0095; #100;
A = 16'h006D; B = 16'h0096; #100;
A = 16'h006D; B = 16'h0097; #100;
A = 16'h006D; B = 16'h0098; #100;
A = 16'h006D; B = 16'h0099; #100;
A = 16'h006D; B = 16'h009A; #100;
A = 16'h006D; B = 16'h009B; #100;
A = 16'h006D; B = 16'h009C; #100;
A = 16'h006D; B = 16'h009D; #100;
A = 16'h006D; B = 16'h009E; #100;
A = 16'h006D; B = 16'h009F; #100;
A = 16'h006D; B = 16'h00A0; #100;
A = 16'h006D; B = 16'h00A1; #100;
A = 16'h006D; B = 16'h00A2; #100;
A = 16'h006D; B = 16'h00A3; #100;
A = 16'h006D; B = 16'h00A4; #100;
A = 16'h006D; B = 16'h00A5; #100;
A = 16'h006D; B = 16'h00A6; #100;
A = 16'h006D; B = 16'h00A7; #100;
A = 16'h006D; B = 16'h00A8; #100;
A = 16'h006D; B = 16'h00A9; #100;
A = 16'h006D; B = 16'h00AA; #100;
A = 16'h006D; B = 16'h00AB; #100;
A = 16'h006D; B = 16'h00AC; #100;
A = 16'h006D; B = 16'h00AD; #100;
A = 16'h006D; B = 16'h00AE; #100;
A = 16'h006D; B = 16'h00AF; #100;
A = 16'h006D; B = 16'h00B0; #100;
A = 16'h006D; B = 16'h00B1; #100;
A = 16'h006D; B = 16'h00B2; #100;
A = 16'h006D; B = 16'h00B3; #100;
A = 16'h006D; B = 16'h00B4; #100;
A = 16'h006D; B = 16'h00B5; #100;
A = 16'h006D; B = 16'h00B6; #100;
A = 16'h006D; B = 16'h00B7; #100;
A = 16'h006D; B = 16'h00B8; #100;
A = 16'h006D; B = 16'h00B9; #100;
A = 16'h006D; B = 16'h00BA; #100;
A = 16'h006D; B = 16'h00BB; #100;
A = 16'h006D; B = 16'h00BC; #100;
A = 16'h006D; B = 16'h00BD; #100;
A = 16'h006D; B = 16'h00BE; #100;
A = 16'h006D; B = 16'h00BF; #100;
A = 16'h006D; B = 16'h00C0; #100;
A = 16'h006D; B = 16'h00C1; #100;
A = 16'h006D; B = 16'h00C2; #100;
A = 16'h006D; B = 16'h00C3; #100;
A = 16'h006D; B = 16'h00C4; #100;
A = 16'h006D; B = 16'h00C5; #100;
A = 16'h006D; B = 16'h00C6; #100;
A = 16'h006D; B = 16'h00C7; #100;
A = 16'h006D; B = 16'h00C8; #100;
A = 16'h006D; B = 16'h00C9; #100;
A = 16'h006D; B = 16'h00CA; #100;
A = 16'h006D; B = 16'h00CB; #100;
A = 16'h006D; B = 16'h00CC; #100;
A = 16'h006D; B = 16'h00CD; #100;
A = 16'h006D; B = 16'h00CE; #100;
A = 16'h006D; B = 16'h00CF; #100;
A = 16'h006D; B = 16'h00D0; #100;
A = 16'h006D; B = 16'h00D1; #100;
A = 16'h006D; B = 16'h00D2; #100;
A = 16'h006D; B = 16'h00D3; #100;
A = 16'h006D; B = 16'h00D4; #100;
A = 16'h006D; B = 16'h00D5; #100;
A = 16'h006D; B = 16'h00D6; #100;
A = 16'h006D; B = 16'h00D7; #100;
A = 16'h006D; B = 16'h00D8; #100;
A = 16'h006D; B = 16'h00D9; #100;
A = 16'h006D; B = 16'h00DA; #100;
A = 16'h006D; B = 16'h00DB; #100;
A = 16'h006D; B = 16'h00DC; #100;
A = 16'h006D; B = 16'h00DD; #100;
A = 16'h006D; B = 16'h00DE; #100;
A = 16'h006D; B = 16'h00DF; #100;
A = 16'h006D; B = 16'h00E0; #100;
A = 16'h006D; B = 16'h00E1; #100;
A = 16'h006D; B = 16'h00E2; #100;
A = 16'h006D; B = 16'h00E3; #100;
A = 16'h006D; B = 16'h00E4; #100;
A = 16'h006D; B = 16'h00E5; #100;
A = 16'h006D; B = 16'h00E6; #100;
A = 16'h006D; B = 16'h00E7; #100;
A = 16'h006D; B = 16'h00E8; #100;
A = 16'h006D; B = 16'h00E9; #100;
A = 16'h006D; B = 16'h00EA; #100;
A = 16'h006D; B = 16'h00EB; #100;
A = 16'h006D; B = 16'h00EC; #100;
A = 16'h006D; B = 16'h00ED; #100;
A = 16'h006D; B = 16'h00EE; #100;
A = 16'h006D; B = 16'h00EF; #100;
A = 16'h006D; B = 16'h00F0; #100;
A = 16'h006D; B = 16'h00F1; #100;
A = 16'h006D; B = 16'h00F2; #100;
A = 16'h006D; B = 16'h00F3; #100;
A = 16'h006D; B = 16'h00F4; #100;
A = 16'h006D; B = 16'h00F5; #100;
A = 16'h006D; B = 16'h00F6; #100;
A = 16'h006D; B = 16'h00F7; #100;
A = 16'h006D; B = 16'h00F8; #100;
A = 16'h006D; B = 16'h00F9; #100;
A = 16'h006D; B = 16'h00FA; #100;
A = 16'h006D; B = 16'h00FB; #100;
A = 16'h006D; B = 16'h00FC; #100;
A = 16'h006D; B = 16'h00FD; #100;
A = 16'h006D; B = 16'h00FE; #100;
A = 16'h006D; B = 16'h00FF; #100;
A = 16'h006E; B = 16'h000; #100;
A = 16'h006E; B = 16'h001; #100;
A = 16'h006E; B = 16'h002; #100;
A = 16'h006E; B = 16'h003; #100;
A = 16'h006E; B = 16'h004; #100;
A = 16'h006E; B = 16'h005; #100;
A = 16'h006E; B = 16'h006; #100;
A = 16'h006E; B = 16'h007; #100;
A = 16'h006E; B = 16'h008; #100;
A = 16'h006E; B = 16'h009; #100;
A = 16'h006E; B = 16'h00A; #100;
A = 16'h006E; B = 16'h00B; #100;
A = 16'h006E; B = 16'h00C; #100;
A = 16'h006E; B = 16'h00D; #100;
A = 16'h006E; B = 16'h00E; #100;
A = 16'h006E; B = 16'h00F; #100;
A = 16'h006E; B = 16'h0010; #100;
A = 16'h006E; B = 16'h0011; #100;
A = 16'h006E; B = 16'h0012; #100;
A = 16'h006E; B = 16'h0013; #100;
A = 16'h006E; B = 16'h0014; #100;
A = 16'h006E; B = 16'h0015; #100;
A = 16'h006E; B = 16'h0016; #100;
A = 16'h006E; B = 16'h0017; #100;
A = 16'h006E; B = 16'h0018; #100;
A = 16'h006E; B = 16'h0019; #100;
A = 16'h006E; B = 16'h001A; #100;
A = 16'h006E; B = 16'h001B; #100;
A = 16'h006E; B = 16'h001C; #100;
A = 16'h006E; B = 16'h001D; #100;
A = 16'h006E; B = 16'h001E; #100;
A = 16'h006E; B = 16'h001F; #100;
A = 16'h006E; B = 16'h0020; #100;
A = 16'h006E; B = 16'h0021; #100;
A = 16'h006E; B = 16'h0022; #100;
A = 16'h006E; B = 16'h0023; #100;
A = 16'h006E; B = 16'h0024; #100;
A = 16'h006E; B = 16'h0025; #100;
A = 16'h006E; B = 16'h0026; #100;
A = 16'h006E; B = 16'h0027; #100;
A = 16'h006E; B = 16'h0028; #100;
A = 16'h006E; B = 16'h0029; #100;
A = 16'h006E; B = 16'h002A; #100;
A = 16'h006E; B = 16'h002B; #100;
A = 16'h006E; B = 16'h002C; #100;
A = 16'h006E; B = 16'h002D; #100;
A = 16'h006E; B = 16'h002E; #100;
A = 16'h006E; B = 16'h002F; #100;
A = 16'h006E; B = 16'h0030; #100;
A = 16'h006E; B = 16'h0031; #100;
A = 16'h006E; B = 16'h0032; #100;
A = 16'h006E; B = 16'h0033; #100;
A = 16'h006E; B = 16'h0034; #100;
A = 16'h006E; B = 16'h0035; #100;
A = 16'h006E; B = 16'h0036; #100;
A = 16'h006E; B = 16'h0037; #100;
A = 16'h006E; B = 16'h0038; #100;
A = 16'h006E; B = 16'h0039; #100;
A = 16'h006E; B = 16'h003A; #100;
A = 16'h006E; B = 16'h003B; #100;
A = 16'h006E; B = 16'h003C; #100;
A = 16'h006E; B = 16'h003D; #100;
A = 16'h006E; B = 16'h003E; #100;
A = 16'h006E; B = 16'h003F; #100;
A = 16'h006E; B = 16'h0040; #100;
A = 16'h006E; B = 16'h0041; #100;
A = 16'h006E; B = 16'h0042; #100;
A = 16'h006E; B = 16'h0043; #100;
A = 16'h006E; B = 16'h0044; #100;
A = 16'h006E; B = 16'h0045; #100;
A = 16'h006E; B = 16'h0046; #100;
A = 16'h006E; B = 16'h0047; #100;
A = 16'h006E; B = 16'h0048; #100;
A = 16'h006E; B = 16'h0049; #100;
A = 16'h006E; B = 16'h004A; #100;
A = 16'h006E; B = 16'h004B; #100;
A = 16'h006E; B = 16'h004C; #100;
A = 16'h006E; B = 16'h004D; #100;
A = 16'h006E; B = 16'h004E; #100;
A = 16'h006E; B = 16'h004F; #100;
A = 16'h006E; B = 16'h0050; #100;
A = 16'h006E; B = 16'h0051; #100;
A = 16'h006E; B = 16'h0052; #100;
A = 16'h006E; B = 16'h0053; #100;
A = 16'h006E; B = 16'h0054; #100;
A = 16'h006E; B = 16'h0055; #100;
A = 16'h006E; B = 16'h0056; #100;
A = 16'h006E; B = 16'h0057; #100;
A = 16'h006E; B = 16'h0058; #100;
A = 16'h006E; B = 16'h0059; #100;
A = 16'h006E; B = 16'h005A; #100;
A = 16'h006E; B = 16'h005B; #100;
A = 16'h006E; B = 16'h005C; #100;
A = 16'h006E; B = 16'h005D; #100;
A = 16'h006E; B = 16'h005E; #100;
A = 16'h006E; B = 16'h005F; #100;
A = 16'h006E; B = 16'h0060; #100;
A = 16'h006E; B = 16'h0061; #100;
A = 16'h006E; B = 16'h0062; #100;
A = 16'h006E; B = 16'h0063; #100;
A = 16'h006E; B = 16'h0064; #100;
A = 16'h006E; B = 16'h0065; #100;
A = 16'h006E; B = 16'h0066; #100;
A = 16'h006E; B = 16'h0067; #100;
A = 16'h006E; B = 16'h0068; #100;
A = 16'h006E; B = 16'h0069; #100;
A = 16'h006E; B = 16'h006A; #100;
A = 16'h006E; B = 16'h006B; #100;
A = 16'h006E; B = 16'h006C; #100;
A = 16'h006E; B = 16'h006D; #100;
A = 16'h006E; B = 16'h006E; #100;
A = 16'h006E; B = 16'h006F; #100;
A = 16'h006E; B = 16'h0070; #100;
A = 16'h006E; B = 16'h0071; #100;
A = 16'h006E; B = 16'h0072; #100;
A = 16'h006E; B = 16'h0073; #100;
A = 16'h006E; B = 16'h0074; #100;
A = 16'h006E; B = 16'h0075; #100;
A = 16'h006E; B = 16'h0076; #100;
A = 16'h006E; B = 16'h0077; #100;
A = 16'h006E; B = 16'h0078; #100;
A = 16'h006E; B = 16'h0079; #100;
A = 16'h006E; B = 16'h007A; #100;
A = 16'h006E; B = 16'h007B; #100;
A = 16'h006E; B = 16'h007C; #100;
A = 16'h006E; B = 16'h007D; #100;
A = 16'h006E; B = 16'h007E; #100;
A = 16'h006E; B = 16'h007F; #100;
A = 16'h006E; B = 16'h0080; #100;
A = 16'h006E; B = 16'h0081; #100;
A = 16'h006E; B = 16'h0082; #100;
A = 16'h006E; B = 16'h0083; #100;
A = 16'h006E; B = 16'h0084; #100;
A = 16'h006E; B = 16'h0085; #100;
A = 16'h006E; B = 16'h0086; #100;
A = 16'h006E; B = 16'h0087; #100;
A = 16'h006E; B = 16'h0088; #100;
A = 16'h006E; B = 16'h0089; #100;
A = 16'h006E; B = 16'h008A; #100;
A = 16'h006E; B = 16'h008B; #100;
A = 16'h006E; B = 16'h008C; #100;
A = 16'h006E; B = 16'h008D; #100;
A = 16'h006E; B = 16'h008E; #100;
A = 16'h006E; B = 16'h008F; #100;
A = 16'h006E; B = 16'h0090; #100;
A = 16'h006E; B = 16'h0091; #100;
A = 16'h006E; B = 16'h0092; #100;
A = 16'h006E; B = 16'h0093; #100;
A = 16'h006E; B = 16'h0094; #100;
A = 16'h006E; B = 16'h0095; #100;
A = 16'h006E; B = 16'h0096; #100;
A = 16'h006E; B = 16'h0097; #100;
A = 16'h006E; B = 16'h0098; #100;
A = 16'h006E; B = 16'h0099; #100;
A = 16'h006E; B = 16'h009A; #100;
A = 16'h006E; B = 16'h009B; #100;
A = 16'h006E; B = 16'h009C; #100;
A = 16'h006E; B = 16'h009D; #100;
A = 16'h006E; B = 16'h009E; #100;
A = 16'h006E; B = 16'h009F; #100;
A = 16'h006E; B = 16'h00A0; #100;
A = 16'h006E; B = 16'h00A1; #100;
A = 16'h006E; B = 16'h00A2; #100;
A = 16'h006E; B = 16'h00A3; #100;
A = 16'h006E; B = 16'h00A4; #100;
A = 16'h006E; B = 16'h00A5; #100;
A = 16'h006E; B = 16'h00A6; #100;
A = 16'h006E; B = 16'h00A7; #100;
A = 16'h006E; B = 16'h00A8; #100;
A = 16'h006E; B = 16'h00A9; #100;
A = 16'h006E; B = 16'h00AA; #100;
A = 16'h006E; B = 16'h00AB; #100;
A = 16'h006E; B = 16'h00AC; #100;
A = 16'h006E; B = 16'h00AD; #100;
A = 16'h006E; B = 16'h00AE; #100;
A = 16'h006E; B = 16'h00AF; #100;
A = 16'h006E; B = 16'h00B0; #100;
A = 16'h006E; B = 16'h00B1; #100;
A = 16'h006E; B = 16'h00B2; #100;
A = 16'h006E; B = 16'h00B3; #100;
A = 16'h006E; B = 16'h00B4; #100;
A = 16'h006E; B = 16'h00B5; #100;
A = 16'h006E; B = 16'h00B6; #100;
A = 16'h006E; B = 16'h00B7; #100;
A = 16'h006E; B = 16'h00B8; #100;
A = 16'h006E; B = 16'h00B9; #100;
A = 16'h006E; B = 16'h00BA; #100;
A = 16'h006E; B = 16'h00BB; #100;
A = 16'h006E; B = 16'h00BC; #100;
A = 16'h006E; B = 16'h00BD; #100;
A = 16'h006E; B = 16'h00BE; #100;
A = 16'h006E; B = 16'h00BF; #100;
A = 16'h006E; B = 16'h00C0; #100;
A = 16'h006E; B = 16'h00C1; #100;
A = 16'h006E; B = 16'h00C2; #100;
A = 16'h006E; B = 16'h00C3; #100;
A = 16'h006E; B = 16'h00C4; #100;
A = 16'h006E; B = 16'h00C5; #100;
A = 16'h006E; B = 16'h00C6; #100;
A = 16'h006E; B = 16'h00C7; #100;
A = 16'h006E; B = 16'h00C8; #100;
A = 16'h006E; B = 16'h00C9; #100;
A = 16'h006E; B = 16'h00CA; #100;
A = 16'h006E; B = 16'h00CB; #100;
A = 16'h006E; B = 16'h00CC; #100;
A = 16'h006E; B = 16'h00CD; #100;
A = 16'h006E; B = 16'h00CE; #100;
A = 16'h006E; B = 16'h00CF; #100;
A = 16'h006E; B = 16'h00D0; #100;
A = 16'h006E; B = 16'h00D1; #100;
A = 16'h006E; B = 16'h00D2; #100;
A = 16'h006E; B = 16'h00D3; #100;
A = 16'h006E; B = 16'h00D4; #100;
A = 16'h006E; B = 16'h00D5; #100;
A = 16'h006E; B = 16'h00D6; #100;
A = 16'h006E; B = 16'h00D7; #100;
A = 16'h006E; B = 16'h00D8; #100;
A = 16'h006E; B = 16'h00D9; #100;
A = 16'h006E; B = 16'h00DA; #100;
A = 16'h006E; B = 16'h00DB; #100;
A = 16'h006E; B = 16'h00DC; #100;
A = 16'h006E; B = 16'h00DD; #100;
A = 16'h006E; B = 16'h00DE; #100;
A = 16'h006E; B = 16'h00DF; #100;
A = 16'h006E; B = 16'h00E0; #100;
A = 16'h006E; B = 16'h00E1; #100;
A = 16'h006E; B = 16'h00E2; #100;
A = 16'h006E; B = 16'h00E3; #100;
A = 16'h006E; B = 16'h00E4; #100;
A = 16'h006E; B = 16'h00E5; #100;
A = 16'h006E; B = 16'h00E6; #100;
A = 16'h006E; B = 16'h00E7; #100;
A = 16'h006E; B = 16'h00E8; #100;
A = 16'h006E; B = 16'h00E9; #100;
A = 16'h006E; B = 16'h00EA; #100;
A = 16'h006E; B = 16'h00EB; #100;
A = 16'h006E; B = 16'h00EC; #100;
A = 16'h006E; B = 16'h00ED; #100;
A = 16'h006E; B = 16'h00EE; #100;
A = 16'h006E; B = 16'h00EF; #100;
A = 16'h006E; B = 16'h00F0; #100;
A = 16'h006E; B = 16'h00F1; #100;
A = 16'h006E; B = 16'h00F2; #100;
A = 16'h006E; B = 16'h00F3; #100;
A = 16'h006E; B = 16'h00F4; #100;
A = 16'h006E; B = 16'h00F5; #100;
A = 16'h006E; B = 16'h00F6; #100;
A = 16'h006E; B = 16'h00F7; #100;
A = 16'h006E; B = 16'h00F8; #100;
A = 16'h006E; B = 16'h00F9; #100;
A = 16'h006E; B = 16'h00FA; #100;
A = 16'h006E; B = 16'h00FB; #100;
A = 16'h006E; B = 16'h00FC; #100;
A = 16'h006E; B = 16'h00FD; #100;
A = 16'h006E; B = 16'h00FE; #100;
A = 16'h006E; B = 16'h00FF; #100;
A = 16'h006F; B = 16'h000; #100;
A = 16'h006F; B = 16'h001; #100;
A = 16'h006F; B = 16'h002; #100;
A = 16'h006F; B = 16'h003; #100;
A = 16'h006F; B = 16'h004; #100;
A = 16'h006F; B = 16'h005; #100;
A = 16'h006F; B = 16'h006; #100;
A = 16'h006F; B = 16'h007; #100;
A = 16'h006F; B = 16'h008; #100;
A = 16'h006F; B = 16'h009; #100;
A = 16'h006F; B = 16'h00A; #100;
A = 16'h006F; B = 16'h00B; #100;
A = 16'h006F; B = 16'h00C; #100;
A = 16'h006F; B = 16'h00D; #100;
A = 16'h006F; B = 16'h00E; #100;
A = 16'h006F; B = 16'h00F; #100;
A = 16'h006F; B = 16'h0010; #100;
A = 16'h006F; B = 16'h0011; #100;
A = 16'h006F; B = 16'h0012; #100;
A = 16'h006F; B = 16'h0013; #100;
A = 16'h006F; B = 16'h0014; #100;
A = 16'h006F; B = 16'h0015; #100;
A = 16'h006F; B = 16'h0016; #100;
A = 16'h006F; B = 16'h0017; #100;
A = 16'h006F; B = 16'h0018; #100;
A = 16'h006F; B = 16'h0019; #100;
A = 16'h006F; B = 16'h001A; #100;
A = 16'h006F; B = 16'h001B; #100;
A = 16'h006F; B = 16'h001C; #100;
A = 16'h006F; B = 16'h001D; #100;
A = 16'h006F; B = 16'h001E; #100;
A = 16'h006F; B = 16'h001F; #100;
A = 16'h006F; B = 16'h0020; #100;
A = 16'h006F; B = 16'h0021; #100;
A = 16'h006F; B = 16'h0022; #100;
A = 16'h006F; B = 16'h0023; #100;
A = 16'h006F; B = 16'h0024; #100;
A = 16'h006F; B = 16'h0025; #100;
A = 16'h006F; B = 16'h0026; #100;
A = 16'h006F; B = 16'h0027; #100;
A = 16'h006F; B = 16'h0028; #100;
A = 16'h006F; B = 16'h0029; #100;
A = 16'h006F; B = 16'h002A; #100;
A = 16'h006F; B = 16'h002B; #100;
A = 16'h006F; B = 16'h002C; #100;
A = 16'h006F; B = 16'h002D; #100;
A = 16'h006F; B = 16'h002E; #100;
A = 16'h006F; B = 16'h002F; #100;
A = 16'h006F; B = 16'h0030; #100;
A = 16'h006F; B = 16'h0031; #100;
A = 16'h006F; B = 16'h0032; #100;
A = 16'h006F; B = 16'h0033; #100;
A = 16'h006F; B = 16'h0034; #100;
A = 16'h006F; B = 16'h0035; #100;
A = 16'h006F; B = 16'h0036; #100;
A = 16'h006F; B = 16'h0037; #100;
A = 16'h006F; B = 16'h0038; #100;
A = 16'h006F; B = 16'h0039; #100;
A = 16'h006F; B = 16'h003A; #100;
A = 16'h006F; B = 16'h003B; #100;
A = 16'h006F; B = 16'h003C; #100;
A = 16'h006F; B = 16'h003D; #100;
A = 16'h006F; B = 16'h003E; #100;
A = 16'h006F; B = 16'h003F; #100;
A = 16'h006F; B = 16'h0040; #100;
A = 16'h006F; B = 16'h0041; #100;
A = 16'h006F; B = 16'h0042; #100;
A = 16'h006F; B = 16'h0043; #100;
A = 16'h006F; B = 16'h0044; #100;
A = 16'h006F; B = 16'h0045; #100;
A = 16'h006F; B = 16'h0046; #100;
A = 16'h006F; B = 16'h0047; #100;
A = 16'h006F; B = 16'h0048; #100;
A = 16'h006F; B = 16'h0049; #100;
A = 16'h006F; B = 16'h004A; #100;
A = 16'h006F; B = 16'h004B; #100;
A = 16'h006F; B = 16'h004C; #100;
A = 16'h006F; B = 16'h004D; #100;
A = 16'h006F; B = 16'h004E; #100;
A = 16'h006F; B = 16'h004F; #100;
A = 16'h006F; B = 16'h0050; #100;
A = 16'h006F; B = 16'h0051; #100;
A = 16'h006F; B = 16'h0052; #100;
A = 16'h006F; B = 16'h0053; #100;
A = 16'h006F; B = 16'h0054; #100;
A = 16'h006F; B = 16'h0055; #100;
A = 16'h006F; B = 16'h0056; #100;
A = 16'h006F; B = 16'h0057; #100;
A = 16'h006F; B = 16'h0058; #100;
A = 16'h006F; B = 16'h0059; #100;
A = 16'h006F; B = 16'h005A; #100;
A = 16'h006F; B = 16'h005B; #100;
A = 16'h006F; B = 16'h005C; #100;
A = 16'h006F; B = 16'h005D; #100;
A = 16'h006F; B = 16'h005E; #100;
A = 16'h006F; B = 16'h005F; #100;
A = 16'h006F; B = 16'h0060; #100;
A = 16'h006F; B = 16'h0061; #100;
A = 16'h006F; B = 16'h0062; #100;
A = 16'h006F; B = 16'h0063; #100;
A = 16'h006F; B = 16'h0064; #100;
A = 16'h006F; B = 16'h0065; #100;
A = 16'h006F; B = 16'h0066; #100;
A = 16'h006F; B = 16'h0067; #100;
A = 16'h006F; B = 16'h0068; #100;
A = 16'h006F; B = 16'h0069; #100;
A = 16'h006F; B = 16'h006A; #100;
A = 16'h006F; B = 16'h006B; #100;
A = 16'h006F; B = 16'h006C; #100;
A = 16'h006F; B = 16'h006D; #100;
A = 16'h006F; B = 16'h006E; #100;
A = 16'h006F; B = 16'h006F; #100;
A = 16'h006F; B = 16'h0070; #100;
A = 16'h006F; B = 16'h0071; #100;
A = 16'h006F; B = 16'h0072; #100;
A = 16'h006F; B = 16'h0073; #100;
A = 16'h006F; B = 16'h0074; #100;
A = 16'h006F; B = 16'h0075; #100;
A = 16'h006F; B = 16'h0076; #100;
A = 16'h006F; B = 16'h0077; #100;
A = 16'h006F; B = 16'h0078; #100;
A = 16'h006F; B = 16'h0079; #100;
A = 16'h006F; B = 16'h007A; #100;
A = 16'h006F; B = 16'h007B; #100;
A = 16'h006F; B = 16'h007C; #100;
A = 16'h006F; B = 16'h007D; #100;
A = 16'h006F; B = 16'h007E; #100;
A = 16'h006F; B = 16'h007F; #100;
A = 16'h006F; B = 16'h0080; #100;
A = 16'h006F; B = 16'h0081; #100;
A = 16'h006F; B = 16'h0082; #100;
A = 16'h006F; B = 16'h0083; #100;
A = 16'h006F; B = 16'h0084; #100;
A = 16'h006F; B = 16'h0085; #100;
A = 16'h006F; B = 16'h0086; #100;
A = 16'h006F; B = 16'h0087; #100;
A = 16'h006F; B = 16'h0088; #100;
A = 16'h006F; B = 16'h0089; #100;
A = 16'h006F; B = 16'h008A; #100;
A = 16'h006F; B = 16'h008B; #100;
A = 16'h006F; B = 16'h008C; #100;
A = 16'h006F; B = 16'h008D; #100;
A = 16'h006F; B = 16'h008E; #100;
A = 16'h006F; B = 16'h008F; #100;
A = 16'h006F; B = 16'h0090; #100;
A = 16'h006F; B = 16'h0091; #100;
A = 16'h006F; B = 16'h0092; #100;
A = 16'h006F; B = 16'h0093; #100;
A = 16'h006F; B = 16'h0094; #100;
A = 16'h006F; B = 16'h0095; #100;
A = 16'h006F; B = 16'h0096; #100;
A = 16'h006F; B = 16'h0097; #100;
A = 16'h006F; B = 16'h0098; #100;
A = 16'h006F; B = 16'h0099; #100;
A = 16'h006F; B = 16'h009A; #100;
A = 16'h006F; B = 16'h009B; #100;
A = 16'h006F; B = 16'h009C; #100;
A = 16'h006F; B = 16'h009D; #100;
A = 16'h006F; B = 16'h009E; #100;
A = 16'h006F; B = 16'h009F; #100;
A = 16'h006F; B = 16'h00A0; #100;
A = 16'h006F; B = 16'h00A1; #100;
A = 16'h006F; B = 16'h00A2; #100;
A = 16'h006F; B = 16'h00A3; #100;
A = 16'h006F; B = 16'h00A4; #100;
A = 16'h006F; B = 16'h00A5; #100;
A = 16'h006F; B = 16'h00A6; #100;
A = 16'h006F; B = 16'h00A7; #100;
A = 16'h006F; B = 16'h00A8; #100;
A = 16'h006F; B = 16'h00A9; #100;
A = 16'h006F; B = 16'h00AA; #100;
A = 16'h006F; B = 16'h00AB; #100;
A = 16'h006F; B = 16'h00AC; #100;
A = 16'h006F; B = 16'h00AD; #100;
A = 16'h006F; B = 16'h00AE; #100;
A = 16'h006F; B = 16'h00AF; #100;
A = 16'h006F; B = 16'h00B0; #100;
A = 16'h006F; B = 16'h00B1; #100;
A = 16'h006F; B = 16'h00B2; #100;
A = 16'h006F; B = 16'h00B3; #100;
A = 16'h006F; B = 16'h00B4; #100;
A = 16'h006F; B = 16'h00B5; #100;
A = 16'h006F; B = 16'h00B6; #100;
A = 16'h006F; B = 16'h00B7; #100;
A = 16'h006F; B = 16'h00B8; #100;
A = 16'h006F; B = 16'h00B9; #100;
A = 16'h006F; B = 16'h00BA; #100;
A = 16'h006F; B = 16'h00BB; #100;
A = 16'h006F; B = 16'h00BC; #100;
A = 16'h006F; B = 16'h00BD; #100;
A = 16'h006F; B = 16'h00BE; #100;
A = 16'h006F; B = 16'h00BF; #100;
A = 16'h006F; B = 16'h00C0; #100;
A = 16'h006F; B = 16'h00C1; #100;
A = 16'h006F; B = 16'h00C2; #100;
A = 16'h006F; B = 16'h00C3; #100;
A = 16'h006F; B = 16'h00C4; #100;
A = 16'h006F; B = 16'h00C5; #100;
A = 16'h006F; B = 16'h00C6; #100;
A = 16'h006F; B = 16'h00C7; #100;
A = 16'h006F; B = 16'h00C8; #100;
A = 16'h006F; B = 16'h00C9; #100;
A = 16'h006F; B = 16'h00CA; #100;
A = 16'h006F; B = 16'h00CB; #100;
A = 16'h006F; B = 16'h00CC; #100;
A = 16'h006F; B = 16'h00CD; #100;
A = 16'h006F; B = 16'h00CE; #100;
A = 16'h006F; B = 16'h00CF; #100;
A = 16'h006F; B = 16'h00D0; #100;
A = 16'h006F; B = 16'h00D1; #100;
A = 16'h006F; B = 16'h00D2; #100;
A = 16'h006F; B = 16'h00D3; #100;
A = 16'h006F; B = 16'h00D4; #100;
A = 16'h006F; B = 16'h00D5; #100;
A = 16'h006F; B = 16'h00D6; #100;
A = 16'h006F; B = 16'h00D7; #100;
A = 16'h006F; B = 16'h00D8; #100;
A = 16'h006F; B = 16'h00D9; #100;
A = 16'h006F; B = 16'h00DA; #100;
A = 16'h006F; B = 16'h00DB; #100;
A = 16'h006F; B = 16'h00DC; #100;
A = 16'h006F; B = 16'h00DD; #100;
A = 16'h006F; B = 16'h00DE; #100;
A = 16'h006F; B = 16'h00DF; #100;
A = 16'h006F; B = 16'h00E0; #100;
A = 16'h006F; B = 16'h00E1; #100;
A = 16'h006F; B = 16'h00E2; #100;
A = 16'h006F; B = 16'h00E3; #100;
A = 16'h006F; B = 16'h00E4; #100;
A = 16'h006F; B = 16'h00E5; #100;
A = 16'h006F; B = 16'h00E6; #100;
A = 16'h006F; B = 16'h00E7; #100;
A = 16'h006F; B = 16'h00E8; #100;
A = 16'h006F; B = 16'h00E9; #100;
A = 16'h006F; B = 16'h00EA; #100;
A = 16'h006F; B = 16'h00EB; #100;
A = 16'h006F; B = 16'h00EC; #100;
A = 16'h006F; B = 16'h00ED; #100;
A = 16'h006F; B = 16'h00EE; #100;
A = 16'h006F; B = 16'h00EF; #100;
A = 16'h006F; B = 16'h00F0; #100;
A = 16'h006F; B = 16'h00F1; #100;
A = 16'h006F; B = 16'h00F2; #100;
A = 16'h006F; B = 16'h00F3; #100;
A = 16'h006F; B = 16'h00F4; #100;
A = 16'h006F; B = 16'h00F5; #100;
A = 16'h006F; B = 16'h00F6; #100;
A = 16'h006F; B = 16'h00F7; #100;
A = 16'h006F; B = 16'h00F8; #100;
A = 16'h006F; B = 16'h00F9; #100;
A = 16'h006F; B = 16'h00FA; #100;
A = 16'h006F; B = 16'h00FB; #100;
A = 16'h006F; B = 16'h00FC; #100;
A = 16'h006F; B = 16'h00FD; #100;
A = 16'h006F; B = 16'h00FE; #100;
A = 16'h006F; B = 16'h00FF; #100;
A = 16'h0070; B = 16'h000; #100;
A = 16'h0070; B = 16'h001; #100;
A = 16'h0070; B = 16'h002; #100;
A = 16'h0070; B = 16'h003; #100;
A = 16'h0070; B = 16'h004; #100;
A = 16'h0070; B = 16'h005; #100;
A = 16'h0070; B = 16'h006; #100;
A = 16'h0070; B = 16'h007; #100;
A = 16'h0070; B = 16'h008; #100;
A = 16'h0070; B = 16'h009; #100;
A = 16'h0070; B = 16'h00A; #100;
A = 16'h0070; B = 16'h00B; #100;
A = 16'h0070; B = 16'h00C; #100;
A = 16'h0070; B = 16'h00D; #100;
A = 16'h0070; B = 16'h00E; #100;
A = 16'h0070; B = 16'h00F; #100;
A = 16'h0070; B = 16'h0010; #100;
A = 16'h0070; B = 16'h0011; #100;
A = 16'h0070; B = 16'h0012; #100;
A = 16'h0070; B = 16'h0013; #100;
A = 16'h0070; B = 16'h0014; #100;
A = 16'h0070; B = 16'h0015; #100;
A = 16'h0070; B = 16'h0016; #100;
A = 16'h0070; B = 16'h0017; #100;
A = 16'h0070; B = 16'h0018; #100;
A = 16'h0070; B = 16'h0019; #100;
A = 16'h0070; B = 16'h001A; #100;
A = 16'h0070; B = 16'h001B; #100;
A = 16'h0070; B = 16'h001C; #100;
A = 16'h0070; B = 16'h001D; #100;
A = 16'h0070; B = 16'h001E; #100;
A = 16'h0070; B = 16'h001F; #100;
A = 16'h0070; B = 16'h0020; #100;
A = 16'h0070; B = 16'h0021; #100;
A = 16'h0070; B = 16'h0022; #100;
A = 16'h0070; B = 16'h0023; #100;
A = 16'h0070; B = 16'h0024; #100;
A = 16'h0070; B = 16'h0025; #100;
A = 16'h0070; B = 16'h0026; #100;
A = 16'h0070; B = 16'h0027; #100;
A = 16'h0070; B = 16'h0028; #100;
A = 16'h0070; B = 16'h0029; #100;
A = 16'h0070; B = 16'h002A; #100;
A = 16'h0070; B = 16'h002B; #100;
A = 16'h0070; B = 16'h002C; #100;
A = 16'h0070; B = 16'h002D; #100;
A = 16'h0070; B = 16'h002E; #100;
A = 16'h0070; B = 16'h002F; #100;
A = 16'h0070; B = 16'h0030; #100;
A = 16'h0070; B = 16'h0031; #100;
A = 16'h0070; B = 16'h0032; #100;
A = 16'h0070; B = 16'h0033; #100;
A = 16'h0070; B = 16'h0034; #100;
A = 16'h0070; B = 16'h0035; #100;
A = 16'h0070; B = 16'h0036; #100;
A = 16'h0070; B = 16'h0037; #100;
A = 16'h0070; B = 16'h0038; #100;
A = 16'h0070; B = 16'h0039; #100;
A = 16'h0070; B = 16'h003A; #100;
A = 16'h0070; B = 16'h003B; #100;
A = 16'h0070; B = 16'h003C; #100;
A = 16'h0070; B = 16'h003D; #100;
A = 16'h0070; B = 16'h003E; #100;
A = 16'h0070; B = 16'h003F; #100;
A = 16'h0070; B = 16'h0040; #100;
A = 16'h0070; B = 16'h0041; #100;
A = 16'h0070; B = 16'h0042; #100;
A = 16'h0070; B = 16'h0043; #100;
A = 16'h0070; B = 16'h0044; #100;
A = 16'h0070; B = 16'h0045; #100;
A = 16'h0070; B = 16'h0046; #100;
A = 16'h0070; B = 16'h0047; #100;
A = 16'h0070; B = 16'h0048; #100;
A = 16'h0070; B = 16'h0049; #100;
A = 16'h0070; B = 16'h004A; #100;
A = 16'h0070; B = 16'h004B; #100;
A = 16'h0070; B = 16'h004C; #100;
A = 16'h0070; B = 16'h004D; #100;
A = 16'h0070; B = 16'h004E; #100;
A = 16'h0070; B = 16'h004F; #100;
A = 16'h0070; B = 16'h0050; #100;
A = 16'h0070; B = 16'h0051; #100;
A = 16'h0070; B = 16'h0052; #100;
A = 16'h0070; B = 16'h0053; #100;
A = 16'h0070; B = 16'h0054; #100;
A = 16'h0070; B = 16'h0055; #100;
A = 16'h0070; B = 16'h0056; #100;
A = 16'h0070; B = 16'h0057; #100;
A = 16'h0070; B = 16'h0058; #100;
A = 16'h0070; B = 16'h0059; #100;
A = 16'h0070; B = 16'h005A; #100;
A = 16'h0070; B = 16'h005B; #100;
A = 16'h0070; B = 16'h005C; #100;
A = 16'h0070; B = 16'h005D; #100;
A = 16'h0070; B = 16'h005E; #100;
A = 16'h0070; B = 16'h005F; #100;
A = 16'h0070; B = 16'h0060; #100;
A = 16'h0070; B = 16'h0061; #100;
A = 16'h0070; B = 16'h0062; #100;
A = 16'h0070; B = 16'h0063; #100;
A = 16'h0070; B = 16'h0064; #100;
A = 16'h0070; B = 16'h0065; #100;
A = 16'h0070; B = 16'h0066; #100;
A = 16'h0070; B = 16'h0067; #100;
A = 16'h0070; B = 16'h0068; #100;
A = 16'h0070; B = 16'h0069; #100;
A = 16'h0070; B = 16'h006A; #100;
A = 16'h0070; B = 16'h006B; #100;
A = 16'h0070; B = 16'h006C; #100;
A = 16'h0070; B = 16'h006D; #100;
A = 16'h0070; B = 16'h006E; #100;
A = 16'h0070; B = 16'h006F; #100;
A = 16'h0070; B = 16'h0070; #100;
A = 16'h0070; B = 16'h0071; #100;
A = 16'h0070; B = 16'h0072; #100;
A = 16'h0070; B = 16'h0073; #100;
A = 16'h0070; B = 16'h0074; #100;
A = 16'h0070; B = 16'h0075; #100;
A = 16'h0070; B = 16'h0076; #100;
A = 16'h0070; B = 16'h0077; #100;
A = 16'h0070; B = 16'h0078; #100;
A = 16'h0070; B = 16'h0079; #100;
A = 16'h0070; B = 16'h007A; #100;
A = 16'h0070; B = 16'h007B; #100;
A = 16'h0070; B = 16'h007C; #100;
A = 16'h0070; B = 16'h007D; #100;
A = 16'h0070; B = 16'h007E; #100;
A = 16'h0070; B = 16'h007F; #100;
A = 16'h0070; B = 16'h0080; #100;
A = 16'h0070; B = 16'h0081; #100;
A = 16'h0070; B = 16'h0082; #100;
A = 16'h0070; B = 16'h0083; #100;
A = 16'h0070; B = 16'h0084; #100;
A = 16'h0070; B = 16'h0085; #100;
A = 16'h0070; B = 16'h0086; #100;
A = 16'h0070; B = 16'h0087; #100;
A = 16'h0070; B = 16'h0088; #100;
A = 16'h0070; B = 16'h0089; #100;
A = 16'h0070; B = 16'h008A; #100;
A = 16'h0070; B = 16'h008B; #100;
A = 16'h0070; B = 16'h008C; #100;
A = 16'h0070; B = 16'h008D; #100;
A = 16'h0070; B = 16'h008E; #100;
A = 16'h0070; B = 16'h008F; #100;
A = 16'h0070; B = 16'h0090; #100;
A = 16'h0070; B = 16'h0091; #100;
A = 16'h0070; B = 16'h0092; #100;
A = 16'h0070; B = 16'h0093; #100;
A = 16'h0070; B = 16'h0094; #100;
A = 16'h0070; B = 16'h0095; #100;
A = 16'h0070; B = 16'h0096; #100;
A = 16'h0070; B = 16'h0097; #100;
A = 16'h0070; B = 16'h0098; #100;
A = 16'h0070; B = 16'h0099; #100;
A = 16'h0070; B = 16'h009A; #100;
A = 16'h0070; B = 16'h009B; #100;
A = 16'h0070; B = 16'h009C; #100;
A = 16'h0070; B = 16'h009D; #100;
A = 16'h0070; B = 16'h009E; #100;
A = 16'h0070; B = 16'h009F; #100;
A = 16'h0070; B = 16'h00A0; #100;
A = 16'h0070; B = 16'h00A1; #100;
A = 16'h0070; B = 16'h00A2; #100;
A = 16'h0070; B = 16'h00A3; #100;
A = 16'h0070; B = 16'h00A4; #100;
A = 16'h0070; B = 16'h00A5; #100;
A = 16'h0070; B = 16'h00A6; #100;
A = 16'h0070; B = 16'h00A7; #100;
A = 16'h0070; B = 16'h00A8; #100;
A = 16'h0070; B = 16'h00A9; #100;
A = 16'h0070; B = 16'h00AA; #100;
A = 16'h0070; B = 16'h00AB; #100;
A = 16'h0070; B = 16'h00AC; #100;
A = 16'h0070; B = 16'h00AD; #100;
A = 16'h0070; B = 16'h00AE; #100;
A = 16'h0070; B = 16'h00AF; #100;
A = 16'h0070; B = 16'h00B0; #100;
A = 16'h0070; B = 16'h00B1; #100;
A = 16'h0070; B = 16'h00B2; #100;
A = 16'h0070; B = 16'h00B3; #100;
A = 16'h0070; B = 16'h00B4; #100;
A = 16'h0070; B = 16'h00B5; #100;
A = 16'h0070; B = 16'h00B6; #100;
A = 16'h0070; B = 16'h00B7; #100;
A = 16'h0070; B = 16'h00B8; #100;
A = 16'h0070; B = 16'h00B9; #100;
A = 16'h0070; B = 16'h00BA; #100;
A = 16'h0070; B = 16'h00BB; #100;
A = 16'h0070; B = 16'h00BC; #100;
A = 16'h0070; B = 16'h00BD; #100;
A = 16'h0070; B = 16'h00BE; #100;
A = 16'h0070; B = 16'h00BF; #100;
A = 16'h0070; B = 16'h00C0; #100;
A = 16'h0070; B = 16'h00C1; #100;
A = 16'h0070; B = 16'h00C2; #100;
A = 16'h0070; B = 16'h00C3; #100;
A = 16'h0070; B = 16'h00C4; #100;
A = 16'h0070; B = 16'h00C5; #100;
A = 16'h0070; B = 16'h00C6; #100;
A = 16'h0070; B = 16'h00C7; #100;
A = 16'h0070; B = 16'h00C8; #100;
A = 16'h0070; B = 16'h00C9; #100;
A = 16'h0070; B = 16'h00CA; #100;
A = 16'h0070; B = 16'h00CB; #100;
A = 16'h0070; B = 16'h00CC; #100;
A = 16'h0070; B = 16'h00CD; #100;
A = 16'h0070; B = 16'h00CE; #100;
A = 16'h0070; B = 16'h00CF; #100;
A = 16'h0070; B = 16'h00D0; #100;
A = 16'h0070; B = 16'h00D1; #100;
A = 16'h0070; B = 16'h00D2; #100;
A = 16'h0070; B = 16'h00D3; #100;
A = 16'h0070; B = 16'h00D4; #100;
A = 16'h0070; B = 16'h00D5; #100;
A = 16'h0070; B = 16'h00D6; #100;
A = 16'h0070; B = 16'h00D7; #100;
A = 16'h0070; B = 16'h00D8; #100;
A = 16'h0070; B = 16'h00D9; #100;
A = 16'h0070; B = 16'h00DA; #100;
A = 16'h0070; B = 16'h00DB; #100;
A = 16'h0070; B = 16'h00DC; #100;
A = 16'h0070; B = 16'h00DD; #100;
A = 16'h0070; B = 16'h00DE; #100;
A = 16'h0070; B = 16'h00DF; #100;
A = 16'h0070; B = 16'h00E0; #100;
A = 16'h0070; B = 16'h00E1; #100;
A = 16'h0070; B = 16'h00E2; #100;
A = 16'h0070; B = 16'h00E3; #100;
A = 16'h0070; B = 16'h00E4; #100;
A = 16'h0070; B = 16'h00E5; #100;
A = 16'h0070; B = 16'h00E6; #100;
A = 16'h0070; B = 16'h00E7; #100;
A = 16'h0070; B = 16'h00E8; #100;
A = 16'h0070; B = 16'h00E9; #100;
A = 16'h0070; B = 16'h00EA; #100;
A = 16'h0070; B = 16'h00EB; #100;
A = 16'h0070; B = 16'h00EC; #100;
A = 16'h0070; B = 16'h00ED; #100;
A = 16'h0070; B = 16'h00EE; #100;
A = 16'h0070; B = 16'h00EF; #100;
A = 16'h0070; B = 16'h00F0; #100;
A = 16'h0070; B = 16'h00F1; #100;
A = 16'h0070; B = 16'h00F2; #100;
A = 16'h0070; B = 16'h00F3; #100;
A = 16'h0070; B = 16'h00F4; #100;
A = 16'h0070; B = 16'h00F5; #100;
A = 16'h0070; B = 16'h00F6; #100;
A = 16'h0070; B = 16'h00F7; #100;
A = 16'h0070; B = 16'h00F8; #100;
A = 16'h0070; B = 16'h00F9; #100;
A = 16'h0070; B = 16'h00FA; #100;
A = 16'h0070; B = 16'h00FB; #100;
A = 16'h0070; B = 16'h00FC; #100;
A = 16'h0070; B = 16'h00FD; #100;
A = 16'h0070; B = 16'h00FE; #100;
A = 16'h0070; B = 16'h00FF; #100;
A = 16'h0071; B = 16'h000; #100;
A = 16'h0071; B = 16'h001; #100;
A = 16'h0071; B = 16'h002; #100;
A = 16'h0071; B = 16'h003; #100;
A = 16'h0071; B = 16'h004; #100;
A = 16'h0071; B = 16'h005; #100;
A = 16'h0071; B = 16'h006; #100;
A = 16'h0071; B = 16'h007; #100;
A = 16'h0071; B = 16'h008; #100;
A = 16'h0071; B = 16'h009; #100;
A = 16'h0071; B = 16'h00A; #100;
A = 16'h0071; B = 16'h00B; #100;
A = 16'h0071; B = 16'h00C; #100;
A = 16'h0071; B = 16'h00D; #100;
A = 16'h0071; B = 16'h00E; #100;
A = 16'h0071; B = 16'h00F; #100;
A = 16'h0071; B = 16'h0010; #100;
A = 16'h0071; B = 16'h0011; #100;
A = 16'h0071; B = 16'h0012; #100;
A = 16'h0071; B = 16'h0013; #100;
A = 16'h0071; B = 16'h0014; #100;
A = 16'h0071; B = 16'h0015; #100;
A = 16'h0071; B = 16'h0016; #100;
A = 16'h0071; B = 16'h0017; #100;
A = 16'h0071; B = 16'h0018; #100;
A = 16'h0071; B = 16'h0019; #100;
A = 16'h0071; B = 16'h001A; #100;
A = 16'h0071; B = 16'h001B; #100;
A = 16'h0071; B = 16'h001C; #100;
A = 16'h0071; B = 16'h001D; #100;
A = 16'h0071; B = 16'h001E; #100;
A = 16'h0071; B = 16'h001F; #100;
A = 16'h0071; B = 16'h0020; #100;
A = 16'h0071; B = 16'h0021; #100;
A = 16'h0071; B = 16'h0022; #100;
A = 16'h0071; B = 16'h0023; #100;
A = 16'h0071; B = 16'h0024; #100;
A = 16'h0071; B = 16'h0025; #100;
A = 16'h0071; B = 16'h0026; #100;
A = 16'h0071; B = 16'h0027; #100;
A = 16'h0071; B = 16'h0028; #100;
A = 16'h0071; B = 16'h0029; #100;
A = 16'h0071; B = 16'h002A; #100;
A = 16'h0071; B = 16'h002B; #100;
A = 16'h0071; B = 16'h002C; #100;
A = 16'h0071; B = 16'h002D; #100;
A = 16'h0071; B = 16'h002E; #100;
A = 16'h0071; B = 16'h002F; #100;
A = 16'h0071; B = 16'h0030; #100;
A = 16'h0071; B = 16'h0031; #100;
A = 16'h0071; B = 16'h0032; #100;
A = 16'h0071; B = 16'h0033; #100;
A = 16'h0071; B = 16'h0034; #100;
A = 16'h0071; B = 16'h0035; #100;
A = 16'h0071; B = 16'h0036; #100;
A = 16'h0071; B = 16'h0037; #100;
A = 16'h0071; B = 16'h0038; #100;
A = 16'h0071; B = 16'h0039; #100;
A = 16'h0071; B = 16'h003A; #100;
A = 16'h0071; B = 16'h003B; #100;
A = 16'h0071; B = 16'h003C; #100;
A = 16'h0071; B = 16'h003D; #100;
A = 16'h0071; B = 16'h003E; #100;
A = 16'h0071; B = 16'h003F; #100;
A = 16'h0071; B = 16'h0040; #100;
A = 16'h0071; B = 16'h0041; #100;
A = 16'h0071; B = 16'h0042; #100;
A = 16'h0071; B = 16'h0043; #100;
A = 16'h0071; B = 16'h0044; #100;
A = 16'h0071; B = 16'h0045; #100;
A = 16'h0071; B = 16'h0046; #100;
A = 16'h0071; B = 16'h0047; #100;
A = 16'h0071; B = 16'h0048; #100;
A = 16'h0071; B = 16'h0049; #100;
A = 16'h0071; B = 16'h004A; #100;
A = 16'h0071; B = 16'h004B; #100;
A = 16'h0071; B = 16'h004C; #100;
A = 16'h0071; B = 16'h004D; #100;
A = 16'h0071; B = 16'h004E; #100;
A = 16'h0071; B = 16'h004F; #100;
A = 16'h0071; B = 16'h0050; #100;
A = 16'h0071; B = 16'h0051; #100;
A = 16'h0071; B = 16'h0052; #100;
A = 16'h0071; B = 16'h0053; #100;
A = 16'h0071; B = 16'h0054; #100;
A = 16'h0071; B = 16'h0055; #100;
A = 16'h0071; B = 16'h0056; #100;
A = 16'h0071; B = 16'h0057; #100;
A = 16'h0071; B = 16'h0058; #100;
A = 16'h0071; B = 16'h0059; #100;
A = 16'h0071; B = 16'h005A; #100;
A = 16'h0071; B = 16'h005B; #100;
A = 16'h0071; B = 16'h005C; #100;
A = 16'h0071; B = 16'h005D; #100;
A = 16'h0071; B = 16'h005E; #100;
A = 16'h0071; B = 16'h005F; #100;
A = 16'h0071; B = 16'h0060; #100;
A = 16'h0071; B = 16'h0061; #100;
A = 16'h0071; B = 16'h0062; #100;
A = 16'h0071; B = 16'h0063; #100;
A = 16'h0071; B = 16'h0064; #100;
A = 16'h0071; B = 16'h0065; #100;
A = 16'h0071; B = 16'h0066; #100;
A = 16'h0071; B = 16'h0067; #100;
A = 16'h0071; B = 16'h0068; #100;
A = 16'h0071; B = 16'h0069; #100;
A = 16'h0071; B = 16'h006A; #100;
A = 16'h0071; B = 16'h006B; #100;
A = 16'h0071; B = 16'h006C; #100;
A = 16'h0071; B = 16'h006D; #100;
A = 16'h0071; B = 16'h006E; #100;
A = 16'h0071; B = 16'h006F; #100;
A = 16'h0071; B = 16'h0070; #100;
A = 16'h0071; B = 16'h0071; #100;
A = 16'h0071; B = 16'h0072; #100;
A = 16'h0071; B = 16'h0073; #100;
A = 16'h0071; B = 16'h0074; #100;
A = 16'h0071; B = 16'h0075; #100;
A = 16'h0071; B = 16'h0076; #100;
A = 16'h0071; B = 16'h0077; #100;
A = 16'h0071; B = 16'h0078; #100;
A = 16'h0071; B = 16'h0079; #100;
A = 16'h0071; B = 16'h007A; #100;
A = 16'h0071; B = 16'h007B; #100;
A = 16'h0071; B = 16'h007C; #100;
A = 16'h0071; B = 16'h007D; #100;
A = 16'h0071; B = 16'h007E; #100;
A = 16'h0071; B = 16'h007F; #100;
A = 16'h0071; B = 16'h0080; #100;
A = 16'h0071; B = 16'h0081; #100;
A = 16'h0071; B = 16'h0082; #100;
A = 16'h0071; B = 16'h0083; #100;
A = 16'h0071; B = 16'h0084; #100;
A = 16'h0071; B = 16'h0085; #100;
A = 16'h0071; B = 16'h0086; #100;
A = 16'h0071; B = 16'h0087; #100;
A = 16'h0071; B = 16'h0088; #100;
A = 16'h0071; B = 16'h0089; #100;
A = 16'h0071; B = 16'h008A; #100;
A = 16'h0071; B = 16'h008B; #100;
A = 16'h0071; B = 16'h008C; #100;
A = 16'h0071; B = 16'h008D; #100;
A = 16'h0071; B = 16'h008E; #100;
A = 16'h0071; B = 16'h008F; #100;
A = 16'h0071; B = 16'h0090; #100;
A = 16'h0071; B = 16'h0091; #100;
A = 16'h0071; B = 16'h0092; #100;
A = 16'h0071; B = 16'h0093; #100;
A = 16'h0071; B = 16'h0094; #100;
A = 16'h0071; B = 16'h0095; #100;
A = 16'h0071; B = 16'h0096; #100;
A = 16'h0071; B = 16'h0097; #100;
A = 16'h0071; B = 16'h0098; #100;
A = 16'h0071; B = 16'h0099; #100;
A = 16'h0071; B = 16'h009A; #100;
A = 16'h0071; B = 16'h009B; #100;
A = 16'h0071; B = 16'h009C; #100;
A = 16'h0071; B = 16'h009D; #100;
A = 16'h0071; B = 16'h009E; #100;
A = 16'h0071; B = 16'h009F; #100;
A = 16'h0071; B = 16'h00A0; #100;
A = 16'h0071; B = 16'h00A1; #100;
A = 16'h0071; B = 16'h00A2; #100;
A = 16'h0071; B = 16'h00A3; #100;
A = 16'h0071; B = 16'h00A4; #100;
A = 16'h0071; B = 16'h00A5; #100;
A = 16'h0071; B = 16'h00A6; #100;
A = 16'h0071; B = 16'h00A7; #100;
A = 16'h0071; B = 16'h00A8; #100;
A = 16'h0071; B = 16'h00A9; #100;
A = 16'h0071; B = 16'h00AA; #100;
A = 16'h0071; B = 16'h00AB; #100;
A = 16'h0071; B = 16'h00AC; #100;
A = 16'h0071; B = 16'h00AD; #100;
A = 16'h0071; B = 16'h00AE; #100;
A = 16'h0071; B = 16'h00AF; #100;
A = 16'h0071; B = 16'h00B0; #100;
A = 16'h0071; B = 16'h00B1; #100;
A = 16'h0071; B = 16'h00B2; #100;
A = 16'h0071; B = 16'h00B3; #100;
A = 16'h0071; B = 16'h00B4; #100;
A = 16'h0071; B = 16'h00B5; #100;
A = 16'h0071; B = 16'h00B6; #100;
A = 16'h0071; B = 16'h00B7; #100;
A = 16'h0071; B = 16'h00B8; #100;
A = 16'h0071; B = 16'h00B9; #100;
A = 16'h0071; B = 16'h00BA; #100;
A = 16'h0071; B = 16'h00BB; #100;
A = 16'h0071; B = 16'h00BC; #100;
A = 16'h0071; B = 16'h00BD; #100;
A = 16'h0071; B = 16'h00BE; #100;
A = 16'h0071; B = 16'h00BF; #100;
A = 16'h0071; B = 16'h00C0; #100;
A = 16'h0071; B = 16'h00C1; #100;
A = 16'h0071; B = 16'h00C2; #100;
A = 16'h0071; B = 16'h00C3; #100;
A = 16'h0071; B = 16'h00C4; #100;
A = 16'h0071; B = 16'h00C5; #100;
A = 16'h0071; B = 16'h00C6; #100;
A = 16'h0071; B = 16'h00C7; #100;
A = 16'h0071; B = 16'h00C8; #100;
A = 16'h0071; B = 16'h00C9; #100;
A = 16'h0071; B = 16'h00CA; #100;
A = 16'h0071; B = 16'h00CB; #100;
A = 16'h0071; B = 16'h00CC; #100;
A = 16'h0071; B = 16'h00CD; #100;
A = 16'h0071; B = 16'h00CE; #100;
A = 16'h0071; B = 16'h00CF; #100;
A = 16'h0071; B = 16'h00D0; #100;
A = 16'h0071; B = 16'h00D1; #100;
A = 16'h0071; B = 16'h00D2; #100;
A = 16'h0071; B = 16'h00D3; #100;
A = 16'h0071; B = 16'h00D4; #100;
A = 16'h0071; B = 16'h00D5; #100;
A = 16'h0071; B = 16'h00D6; #100;
A = 16'h0071; B = 16'h00D7; #100;
A = 16'h0071; B = 16'h00D8; #100;
A = 16'h0071; B = 16'h00D9; #100;
A = 16'h0071; B = 16'h00DA; #100;
A = 16'h0071; B = 16'h00DB; #100;
A = 16'h0071; B = 16'h00DC; #100;
A = 16'h0071; B = 16'h00DD; #100;
A = 16'h0071; B = 16'h00DE; #100;
A = 16'h0071; B = 16'h00DF; #100;
A = 16'h0071; B = 16'h00E0; #100;
A = 16'h0071; B = 16'h00E1; #100;
A = 16'h0071; B = 16'h00E2; #100;
A = 16'h0071; B = 16'h00E3; #100;
A = 16'h0071; B = 16'h00E4; #100;
A = 16'h0071; B = 16'h00E5; #100;
A = 16'h0071; B = 16'h00E6; #100;
A = 16'h0071; B = 16'h00E7; #100;
A = 16'h0071; B = 16'h00E8; #100;
A = 16'h0071; B = 16'h00E9; #100;
A = 16'h0071; B = 16'h00EA; #100;
A = 16'h0071; B = 16'h00EB; #100;
A = 16'h0071; B = 16'h00EC; #100;
A = 16'h0071; B = 16'h00ED; #100;
A = 16'h0071; B = 16'h00EE; #100;
A = 16'h0071; B = 16'h00EF; #100;
A = 16'h0071; B = 16'h00F0; #100;
A = 16'h0071; B = 16'h00F1; #100;
A = 16'h0071; B = 16'h00F2; #100;
A = 16'h0071; B = 16'h00F3; #100;
A = 16'h0071; B = 16'h00F4; #100;
A = 16'h0071; B = 16'h00F5; #100;
A = 16'h0071; B = 16'h00F6; #100;
A = 16'h0071; B = 16'h00F7; #100;
A = 16'h0071; B = 16'h00F8; #100;
A = 16'h0071; B = 16'h00F9; #100;
A = 16'h0071; B = 16'h00FA; #100;
A = 16'h0071; B = 16'h00FB; #100;
A = 16'h0071; B = 16'h00FC; #100;
A = 16'h0071; B = 16'h00FD; #100;
A = 16'h0071; B = 16'h00FE; #100;
A = 16'h0071; B = 16'h00FF; #100;
A = 16'h0072; B = 16'h000; #100;
A = 16'h0072; B = 16'h001; #100;
A = 16'h0072; B = 16'h002; #100;
A = 16'h0072; B = 16'h003; #100;
A = 16'h0072; B = 16'h004; #100;
A = 16'h0072; B = 16'h005; #100;
A = 16'h0072; B = 16'h006; #100;
A = 16'h0072; B = 16'h007; #100;
A = 16'h0072; B = 16'h008; #100;
A = 16'h0072; B = 16'h009; #100;
A = 16'h0072; B = 16'h00A; #100;
A = 16'h0072; B = 16'h00B; #100;
A = 16'h0072; B = 16'h00C; #100;
A = 16'h0072; B = 16'h00D; #100;
A = 16'h0072; B = 16'h00E; #100;
A = 16'h0072; B = 16'h00F; #100;
A = 16'h0072; B = 16'h0010; #100;
A = 16'h0072; B = 16'h0011; #100;
A = 16'h0072; B = 16'h0012; #100;
A = 16'h0072; B = 16'h0013; #100;
A = 16'h0072; B = 16'h0014; #100;
A = 16'h0072; B = 16'h0015; #100;
A = 16'h0072; B = 16'h0016; #100;
A = 16'h0072; B = 16'h0017; #100;
A = 16'h0072; B = 16'h0018; #100;
A = 16'h0072; B = 16'h0019; #100;
A = 16'h0072; B = 16'h001A; #100;
A = 16'h0072; B = 16'h001B; #100;
A = 16'h0072; B = 16'h001C; #100;
A = 16'h0072; B = 16'h001D; #100;
A = 16'h0072; B = 16'h001E; #100;
A = 16'h0072; B = 16'h001F; #100;
A = 16'h0072; B = 16'h0020; #100;
A = 16'h0072; B = 16'h0021; #100;
A = 16'h0072; B = 16'h0022; #100;
A = 16'h0072; B = 16'h0023; #100;
A = 16'h0072; B = 16'h0024; #100;
A = 16'h0072; B = 16'h0025; #100;
A = 16'h0072; B = 16'h0026; #100;
A = 16'h0072; B = 16'h0027; #100;
A = 16'h0072; B = 16'h0028; #100;
A = 16'h0072; B = 16'h0029; #100;
A = 16'h0072; B = 16'h002A; #100;
A = 16'h0072; B = 16'h002B; #100;
A = 16'h0072; B = 16'h002C; #100;
A = 16'h0072; B = 16'h002D; #100;
A = 16'h0072; B = 16'h002E; #100;
A = 16'h0072; B = 16'h002F; #100;
A = 16'h0072; B = 16'h0030; #100;
A = 16'h0072; B = 16'h0031; #100;
A = 16'h0072; B = 16'h0032; #100;
A = 16'h0072; B = 16'h0033; #100;
A = 16'h0072; B = 16'h0034; #100;
A = 16'h0072; B = 16'h0035; #100;
A = 16'h0072; B = 16'h0036; #100;
A = 16'h0072; B = 16'h0037; #100;
A = 16'h0072; B = 16'h0038; #100;
A = 16'h0072; B = 16'h0039; #100;
A = 16'h0072; B = 16'h003A; #100;
A = 16'h0072; B = 16'h003B; #100;
A = 16'h0072; B = 16'h003C; #100;
A = 16'h0072; B = 16'h003D; #100;
A = 16'h0072; B = 16'h003E; #100;
A = 16'h0072; B = 16'h003F; #100;
A = 16'h0072; B = 16'h0040; #100;
A = 16'h0072; B = 16'h0041; #100;
A = 16'h0072; B = 16'h0042; #100;
A = 16'h0072; B = 16'h0043; #100;
A = 16'h0072; B = 16'h0044; #100;
A = 16'h0072; B = 16'h0045; #100;
A = 16'h0072; B = 16'h0046; #100;
A = 16'h0072; B = 16'h0047; #100;
A = 16'h0072; B = 16'h0048; #100;
A = 16'h0072; B = 16'h0049; #100;
A = 16'h0072; B = 16'h004A; #100;
A = 16'h0072; B = 16'h004B; #100;
A = 16'h0072; B = 16'h004C; #100;
A = 16'h0072; B = 16'h004D; #100;
A = 16'h0072; B = 16'h004E; #100;
A = 16'h0072; B = 16'h004F; #100;
A = 16'h0072; B = 16'h0050; #100;
A = 16'h0072; B = 16'h0051; #100;
A = 16'h0072; B = 16'h0052; #100;
A = 16'h0072; B = 16'h0053; #100;
A = 16'h0072; B = 16'h0054; #100;
A = 16'h0072; B = 16'h0055; #100;
A = 16'h0072; B = 16'h0056; #100;
A = 16'h0072; B = 16'h0057; #100;
A = 16'h0072; B = 16'h0058; #100;
A = 16'h0072; B = 16'h0059; #100;
A = 16'h0072; B = 16'h005A; #100;
A = 16'h0072; B = 16'h005B; #100;
A = 16'h0072; B = 16'h005C; #100;
A = 16'h0072; B = 16'h005D; #100;
A = 16'h0072; B = 16'h005E; #100;
A = 16'h0072; B = 16'h005F; #100;
A = 16'h0072; B = 16'h0060; #100;
A = 16'h0072; B = 16'h0061; #100;
A = 16'h0072; B = 16'h0062; #100;
A = 16'h0072; B = 16'h0063; #100;
A = 16'h0072; B = 16'h0064; #100;
A = 16'h0072; B = 16'h0065; #100;
A = 16'h0072; B = 16'h0066; #100;
A = 16'h0072; B = 16'h0067; #100;
A = 16'h0072; B = 16'h0068; #100;
A = 16'h0072; B = 16'h0069; #100;
A = 16'h0072; B = 16'h006A; #100;
A = 16'h0072; B = 16'h006B; #100;
A = 16'h0072; B = 16'h006C; #100;
A = 16'h0072; B = 16'h006D; #100;
A = 16'h0072; B = 16'h006E; #100;
A = 16'h0072; B = 16'h006F; #100;
A = 16'h0072; B = 16'h0070; #100;
A = 16'h0072; B = 16'h0071; #100;
A = 16'h0072; B = 16'h0072; #100;
A = 16'h0072; B = 16'h0073; #100;
A = 16'h0072; B = 16'h0074; #100;
A = 16'h0072; B = 16'h0075; #100;
A = 16'h0072; B = 16'h0076; #100;
A = 16'h0072; B = 16'h0077; #100;
A = 16'h0072; B = 16'h0078; #100;
A = 16'h0072; B = 16'h0079; #100;
A = 16'h0072; B = 16'h007A; #100;
A = 16'h0072; B = 16'h007B; #100;
A = 16'h0072; B = 16'h007C; #100;
A = 16'h0072; B = 16'h007D; #100;
A = 16'h0072; B = 16'h007E; #100;
A = 16'h0072; B = 16'h007F; #100;
A = 16'h0072; B = 16'h0080; #100;
A = 16'h0072; B = 16'h0081; #100;
A = 16'h0072; B = 16'h0082; #100;
A = 16'h0072; B = 16'h0083; #100;
A = 16'h0072; B = 16'h0084; #100;
A = 16'h0072; B = 16'h0085; #100;
A = 16'h0072; B = 16'h0086; #100;
A = 16'h0072; B = 16'h0087; #100;
A = 16'h0072; B = 16'h0088; #100;
A = 16'h0072; B = 16'h0089; #100;
A = 16'h0072; B = 16'h008A; #100;
A = 16'h0072; B = 16'h008B; #100;
A = 16'h0072; B = 16'h008C; #100;
A = 16'h0072; B = 16'h008D; #100;
A = 16'h0072; B = 16'h008E; #100;
A = 16'h0072; B = 16'h008F; #100;
A = 16'h0072; B = 16'h0090; #100;
A = 16'h0072; B = 16'h0091; #100;
A = 16'h0072; B = 16'h0092; #100;
A = 16'h0072; B = 16'h0093; #100;
A = 16'h0072; B = 16'h0094; #100;
A = 16'h0072; B = 16'h0095; #100;
A = 16'h0072; B = 16'h0096; #100;
A = 16'h0072; B = 16'h0097; #100;
A = 16'h0072; B = 16'h0098; #100;
A = 16'h0072; B = 16'h0099; #100;
A = 16'h0072; B = 16'h009A; #100;
A = 16'h0072; B = 16'h009B; #100;
A = 16'h0072; B = 16'h009C; #100;
A = 16'h0072; B = 16'h009D; #100;
A = 16'h0072; B = 16'h009E; #100;
A = 16'h0072; B = 16'h009F; #100;
A = 16'h0072; B = 16'h00A0; #100;
A = 16'h0072; B = 16'h00A1; #100;
A = 16'h0072; B = 16'h00A2; #100;
A = 16'h0072; B = 16'h00A3; #100;
A = 16'h0072; B = 16'h00A4; #100;
A = 16'h0072; B = 16'h00A5; #100;
A = 16'h0072; B = 16'h00A6; #100;
A = 16'h0072; B = 16'h00A7; #100;
A = 16'h0072; B = 16'h00A8; #100;
A = 16'h0072; B = 16'h00A9; #100;
A = 16'h0072; B = 16'h00AA; #100;
A = 16'h0072; B = 16'h00AB; #100;
A = 16'h0072; B = 16'h00AC; #100;
A = 16'h0072; B = 16'h00AD; #100;
A = 16'h0072; B = 16'h00AE; #100;
A = 16'h0072; B = 16'h00AF; #100;
A = 16'h0072; B = 16'h00B0; #100;
A = 16'h0072; B = 16'h00B1; #100;
A = 16'h0072; B = 16'h00B2; #100;
A = 16'h0072; B = 16'h00B3; #100;
A = 16'h0072; B = 16'h00B4; #100;
A = 16'h0072; B = 16'h00B5; #100;
A = 16'h0072; B = 16'h00B6; #100;
A = 16'h0072; B = 16'h00B7; #100;
A = 16'h0072; B = 16'h00B8; #100;
A = 16'h0072; B = 16'h00B9; #100;
A = 16'h0072; B = 16'h00BA; #100;
A = 16'h0072; B = 16'h00BB; #100;
A = 16'h0072; B = 16'h00BC; #100;
A = 16'h0072; B = 16'h00BD; #100;
A = 16'h0072; B = 16'h00BE; #100;
A = 16'h0072; B = 16'h00BF; #100;
A = 16'h0072; B = 16'h00C0; #100;
A = 16'h0072; B = 16'h00C1; #100;
A = 16'h0072; B = 16'h00C2; #100;
A = 16'h0072; B = 16'h00C3; #100;
A = 16'h0072; B = 16'h00C4; #100;
A = 16'h0072; B = 16'h00C5; #100;
A = 16'h0072; B = 16'h00C6; #100;
A = 16'h0072; B = 16'h00C7; #100;
A = 16'h0072; B = 16'h00C8; #100;
A = 16'h0072; B = 16'h00C9; #100;
A = 16'h0072; B = 16'h00CA; #100;
A = 16'h0072; B = 16'h00CB; #100;
A = 16'h0072; B = 16'h00CC; #100;
A = 16'h0072; B = 16'h00CD; #100;
A = 16'h0072; B = 16'h00CE; #100;
A = 16'h0072; B = 16'h00CF; #100;
A = 16'h0072; B = 16'h00D0; #100;
A = 16'h0072; B = 16'h00D1; #100;
A = 16'h0072; B = 16'h00D2; #100;
A = 16'h0072; B = 16'h00D3; #100;
A = 16'h0072; B = 16'h00D4; #100;
A = 16'h0072; B = 16'h00D5; #100;
A = 16'h0072; B = 16'h00D6; #100;
A = 16'h0072; B = 16'h00D7; #100;
A = 16'h0072; B = 16'h00D8; #100;
A = 16'h0072; B = 16'h00D9; #100;
A = 16'h0072; B = 16'h00DA; #100;
A = 16'h0072; B = 16'h00DB; #100;
A = 16'h0072; B = 16'h00DC; #100;
A = 16'h0072; B = 16'h00DD; #100;
A = 16'h0072; B = 16'h00DE; #100;
A = 16'h0072; B = 16'h00DF; #100;
A = 16'h0072; B = 16'h00E0; #100;
A = 16'h0072; B = 16'h00E1; #100;
A = 16'h0072; B = 16'h00E2; #100;
A = 16'h0072; B = 16'h00E3; #100;
A = 16'h0072; B = 16'h00E4; #100;
A = 16'h0072; B = 16'h00E5; #100;
A = 16'h0072; B = 16'h00E6; #100;
A = 16'h0072; B = 16'h00E7; #100;
A = 16'h0072; B = 16'h00E8; #100;
A = 16'h0072; B = 16'h00E9; #100;
A = 16'h0072; B = 16'h00EA; #100;
A = 16'h0072; B = 16'h00EB; #100;
A = 16'h0072; B = 16'h00EC; #100;
A = 16'h0072; B = 16'h00ED; #100;
A = 16'h0072; B = 16'h00EE; #100;
A = 16'h0072; B = 16'h00EF; #100;
A = 16'h0072; B = 16'h00F0; #100;
A = 16'h0072; B = 16'h00F1; #100;
A = 16'h0072; B = 16'h00F2; #100;
A = 16'h0072; B = 16'h00F3; #100;
A = 16'h0072; B = 16'h00F4; #100;
A = 16'h0072; B = 16'h00F5; #100;
A = 16'h0072; B = 16'h00F6; #100;
A = 16'h0072; B = 16'h00F7; #100;
A = 16'h0072; B = 16'h00F8; #100;
A = 16'h0072; B = 16'h00F9; #100;
A = 16'h0072; B = 16'h00FA; #100;
A = 16'h0072; B = 16'h00FB; #100;
A = 16'h0072; B = 16'h00FC; #100;
A = 16'h0072; B = 16'h00FD; #100;
A = 16'h0072; B = 16'h00FE; #100;
A = 16'h0072; B = 16'h00FF; #100;
A = 16'h0073; B = 16'h000; #100;
A = 16'h0073; B = 16'h001; #100;
A = 16'h0073; B = 16'h002; #100;
A = 16'h0073; B = 16'h003; #100;
A = 16'h0073; B = 16'h004; #100;
A = 16'h0073; B = 16'h005; #100;
A = 16'h0073; B = 16'h006; #100;
A = 16'h0073; B = 16'h007; #100;
A = 16'h0073; B = 16'h008; #100;
A = 16'h0073; B = 16'h009; #100;
A = 16'h0073; B = 16'h00A; #100;
A = 16'h0073; B = 16'h00B; #100;
A = 16'h0073; B = 16'h00C; #100;
A = 16'h0073; B = 16'h00D; #100;
A = 16'h0073; B = 16'h00E; #100;
A = 16'h0073; B = 16'h00F; #100;
A = 16'h0073; B = 16'h0010; #100;
A = 16'h0073; B = 16'h0011; #100;
A = 16'h0073; B = 16'h0012; #100;
A = 16'h0073; B = 16'h0013; #100;
A = 16'h0073; B = 16'h0014; #100;
A = 16'h0073; B = 16'h0015; #100;
A = 16'h0073; B = 16'h0016; #100;
A = 16'h0073; B = 16'h0017; #100;
A = 16'h0073; B = 16'h0018; #100;
A = 16'h0073; B = 16'h0019; #100;
A = 16'h0073; B = 16'h001A; #100;
A = 16'h0073; B = 16'h001B; #100;
A = 16'h0073; B = 16'h001C; #100;
A = 16'h0073; B = 16'h001D; #100;
A = 16'h0073; B = 16'h001E; #100;
A = 16'h0073; B = 16'h001F; #100;
A = 16'h0073; B = 16'h0020; #100;
A = 16'h0073; B = 16'h0021; #100;
A = 16'h0073; B = 16'h0022; #100;
A = 16'h0073; B = 16'h0023; #100;
A = 16'h0073; B = 16'h0024; #100;
A = 16'h0073; B = 16'h0025; #100;
A = 16'h0073; B = 16'h0026; #100;
A = 16'h0073; B = 16'h0027; #100;
A = 16'h0073; B = 16'h0028; #100;
A = 16'h0073; B = 16'h0029; #100;
A = 16'h0073; B = 16'h002A; #100;
A = 16'h0073; B = 16'h002B; #100;
A = 16'h0073; B = 16'h002C; #100;
A = 16'h0073; B = 16'h002D; #100;
A = 16'h0073; B = 16'h002E; #100;
A = 16'h0073; B = 16'h002F; #100;
A = 16'h0073; B = 16'h0030; #100;
A = 16'h0073; B = 16'h0031; #100;
A = 16'h0073; B = 16'h0032; #100;
A = 16'h0073; B = 16'h0033; #100;
A = 16'h0073; B = 16'h0034; #100;
A = 16'h0073; B = 16'h0035; #100;
A = 16'h0073; B = 16'h0036; #100;
A = 16'h0073; B = 16'h0037; #100;
A = 16'h0073; B = 16'h0038; #100;
A = 16'h0073; B = 16'h0039; #100;
A = 16'h0073; B = 16'h003A; #100;
A = 16'h0073; B = 16'h003B; #100;
A = 16'h0073; B = 16'h003C; #100;
A = 16'h0073; B = 16'h003D; #100;
A = 16'h0073; B = 16'h003E; #100;
A = 16'h0073; B = 16'h003F; #100;
A = 16'h0073; B = 16'h0040; #100;
A = 16'h0073; B = 16'h0041; #100;
A = 16'h0073; B = 16'h0042; #100;
A = 16'h0073; B = 16'h0043; #100;
A = 16'h0073; B = 16'h0044; #100;
A = 16'h0073; B = 16'h0045; #100;
A = 16'h0073; B = 16'h0046; #100;
A = 16'h0073; B = 16'h0047; #100;
A = 16'h0073; B = 16'h0048; #100;
A = 16'h0073; B = 16'h0049; #100;
A = 16'h0073; B = 16'h004A; #100;
A = 16'h0073; B = 16'h004B; #100;
A = 16'h0073; B = 16'h004C; #100;
A = 16'h0073; B = 16'h004D; #100;
A = 16'h0073; B = 16'h004E; #100;
A = 16'h0073; B = 16'h004F; #100;
A = 16'h0073; B = 16'h0050; #100;
A = 16'h0073; B = 16'h0051; #100;
A = 16'h0073; B = 16'h0052; #100;
A = 16'h0073; B = 16'h0053; #100;
A = 16'h0073; B = 16'h0054; #100;
A = 16'h0073; B = 16'h0055; #100;
A = 16'h0073; B = 16'h0056; #100;
A = 16'h0073; B = 16'h0057; #100;
A = 16'h0073; B = 16'h0058; #100;
A = 16'h0073; B = 16'h0059; #100;
A = 16'h0073; B = 16'h005A; #100;
A = 16'h0073; B = 16'h005B; #100;
A = 16'h0073; B = 16'h005C; #100;
A = 16'h0073; B = 16'h005D; #100;
A = 16'h0073; B = 16'h005E; #100;
A = 16'h0073; B = 16'h005F; #100;
A = 16'h0073; B = 16'h0060; #100;
A = 16'h0073; B = 16'h0061; #100;
A = 16'h0073; B = 16'h0062; #100;
A = 16'h0073; B = 16'h0063; #100;
A = 16'h0073; B = 16'h0064; #100;
A = 16'h0073; B = 16'h0065; #100;
A = 16'h0073; B = 16'h0066; #100;
A = 16'h0073; B = 16'h0067; #100;
A = 16'h0073; B = 16'h0068; #100;
A = 16'h0073; B = 16'h0069; #100;
A = 16'h0073; B = 16'h006A; #100;
A = 16'h0073; B = 16'h006B; #100;
A = 16'h0073; B = 16'h006C; #100;
A = 16'h0073; B = 16'h006D; #100;
A = 16'h0073; B = 16'h006E; #100;
A = 16'h0073; B = 16'h006F; #100;
A = 16'h0073; B = 16'h0070; #100;
A = 16'h0073; B = 16'h0071; #100;
A = 16'h0073; B = 16'h0072; #100;
A = 16'h0073; B = 16'h0073; #100;
A = 16'h0073; B = 16'h0074; #100;
A = 16'h0073; B = 16'h0075; #100;
A = 16'h0073; B = 16'h0076; #100;
A = 16'h0073; B = 16'h0077; #100;
A = 16'h0073; B = 16'h0078; #100;
A = 16'h0073; B = 16'h0079; #100;
A = 16'h0073; B = 16'h007A; #100;
A = 16'h0073; B = 16'h007B; #100;
A = 16'h0073; B = 16'h007C; #100;
A = 16'h0073; B = 16'h007D; #100;
A = 16'h0073; B = 16'h007E; #100;
A = 16'h0073; B = 16'h007F; #100;
A = 16'h0073; B = 16'h0080; #100;
A = 16'h0073; B = 16'h0081; #100;
A = 16'h0073; B = 16'h0082; #100;
A = 16'h0073; B = 16'h0083; #100;
A = 16'h0073; B = 16'h0084; #100;
A = 16'h0073; B = 16'h0085; #100;
A = 16'h0073; B = 16'h0086; #100;
A = 16'h0073; B = 16'h0087; #100;
A = 16'h0073; B = 16'h0088; #100;
A = 16'h0073; B = 16'h0089; #100;
A = 16'h0073; B = 16'h008A; #100;
A = 16'h0073; B = 16'h008B; #100;
A = 16'h0073; B = 16'h008C; #100;
A = 16'h0073; B = 16'h008D; #100;
A = 16'h0073; B = 16'h008E; #100;
A = 16'h0073; B = 16'h008F; #100;
A = 16'h0073; B = 16'h0090; #100;
A = 16'h0073; B = 16'h0091; #100;
A = 16'h0073; B = 16'h0092; #100;
A = 16'h0073; B = 16'h0093; #100;
A = 16'h0073; B = 16'h0094; #100;
A = 16'h0073; B = 16'h0095; #100;
A = 16'h0073; B = 16'h0096; #100;
A = 16'h0073; B = 16'h0097; #100;
A = 16'h0073; B = 16'h0098; #100;
A = 16'h0073; B = 16'h0099; #100;
A = 16'h0073; B = 16'h009A; #100;
A = 16'h0073; B = 16'h009B; #100;
A = 16'h0073; B = 16'h009C; #100;
A = 16'h0073; B = 16'h009D; #100;
A = 16'h0073; B = 16'h009E; #100;
A = 16'h0073; B = 16'h009F; #100;
A = 16'h0073; B = 16'h00A0; #100;
A = 16'h0073; B = 16'h00A1; #100;
A = 16'h0073; B = 16'h00A2; #100;
A = 16'h0073; B = 16'h00A3; #100;
A = 16'h0073; B = 16'h00A4; #100;
A = 16'h0073; B = 16'h00A5; #100;
A = 16'h0073; B = 16'h00A6; #100;
A = 16'h0073; B = 16'h00A7; #100;
A = 16'h0073; B = 16'h00A8; #100;
A = 16'h0073; B = 16'h00A9; #100;
A = 16'h0073; B = 16'h00AA; #100;
A = 16'h0073; B = 16'h00AB; #100;
A = 16'h0073; B = 16'h00AC; #100;
A = 16'h0073; B = 16'h00AD; #100;
A = 16'h0073; B = 16'h00AE; #100;
A = 16'h0073; B = 16'h00AF; #100;
A = 16'h0073; B = 16'h00B0; #100;
A = 16'h0073; B = 16'h00B1; #100;
A = 16'h0073; B = 16'h00B2; #100;
A = 16'h0073; B = 16'h00B3; #100;
A = 16'h0073; B = 16'h00B4; #100;
A = 16'h0073; B = 16'h00B5; #100;
A = 16'h0073; B = 16'h00B6; #100;
A = 16'h0073; B = 16'h00B7; #100;
A = 16'h0073; B = 16'h00B8; #100;
A = 16'h0073; B = 16'h00B9; #100;
A = 16'h0073; B = 16'h00BA; #100;
A = 16'h0073; B = 16'h00BB; #100;
A = 16'h0073; B = 16'h00BC; #100;
A = 16'h0073; B = 16'h00BD; #100;
A = 16'h0073; B = 16'h00BE; #100;
A = 16'h0073; B = 16'h00BF; #100;
A = 16'h0073; B = 16'h00C0; #100;
A = 16'h0073; B = 16'h00C1; #100;
A = 16'h0073; B = 16'h00C2; #100;
A = 16'h0073; B = 16'h00C3; #100;
A = 16'h0073; B = 16'h00C4; #100;
A = 16'h0073; B = 16'h00C5; #100;
A = 16'h0073; B = 16'h00C6; #100;
A = 16'h0073; B = 16'h00C7; #100;
A = 16'h0073; B = 16'h00C8; #100;
A = 16'h0073; B = 16'h00C9; #100;
A = 16'h0073; B = 16'h00CA; #100;
A = 16'h0073; B = 16'h00CB; #100;
A = 16'h0073; B = 16'h00CC; #100;
A = 16'h0073; B = 16'h00CD; #100;
A = 16'h0073; B = 16'h00CE; #100;
A = 16'h0073; B = 16'h00CF; #100;
A = 16'h0073; B = 16'h00D0; #100;
A = 16'h0073; B = 16'h00D1; #100;
A = 16'h0073; B = 16'h00D2; #100;
A = 16'h0073; B = 16'h00D3; #100;
A = 16'h0073; B = 16'h00D4; #100;
A = 16'h0073; B = 16'h00D5; #100;
A = 16'h0073; B = 16'h00D6; #100;
A = 16'h0073; B = 16'h00D7; #100;
A = 16'h0073; B = 16'h00D8; #100;
A = 16'h0073; B = 16'h00D9; #100;
A = 16'h0073; B = 16'h00DA; #100;
A = 16'h0073; B = 16'h00DB; #100;
A = 16'h0073; B = 16'h00DC; #100;
A = 16'h0073; B = 16'h00DD; #100;
A = 16'h0073; B = 16'h00DE; #100;
A = 16'h0073; B = 16'h00DF; #100;
A = 16'h0073; B = 16'h00E0; #100;
A = 16'h0073; B = 16'h00E1; #100;
A = 16'h0073; B = 16'h00E2; #100;
A = 16'h0073; B = 16'h00E3; #100;
A = 16'h0073; B = 16'h00E4; #100;
A = 16'h0073; B = 16'h00E5; #100;
A = 16'h0073; B = 16'h00E6; #100;
A = 16'h0073; B = 16'h00E7; #100;
A = 16'h0073; B = 16'h00E8; #100;
A = 16'h0073; B = 16'h00E9; #100;
A = 16'h0073; B = 16'h00EA; #100;
A = 16'h0073; B = 16'h00EB; #100;
A = 16'h0073; B = 16'h00EC; #100;
A = 16'h0073; B = 16'h00ED; #100;
A = 16'h0073; B = 16'h00EE; #100;
A = 16'h0073; B = 16'h00EF; #100;
A = 16'h0073; B = 16'h00F0; #100;
A = 16'h0073; B = 16'h00F1; #100;
A = 16'h0073; B = 16'h00F2; #100;
A = 16'h0073; B = 16'h00F3; #100;
A = 16'h0073; B = 16'h00F4; #100;
A = 16'h0073; B = 16'h00F5; #100;
A = 16'h0073; B = 16'h00F6; #100;
A = 16'h0073; B = 16'h00F7; #100;
A = 16'h0073; B = 16'h00F8; #100;
A = 16'h0073; B = 16'h00F9; #100;
A = 16'h0073; B = 16'h00FA; #100;
A = 16'h0073; B = 16'h00FB; #100;
A = 16'h0073; B = 16'h00FC; #100;
A = 16'h0073; B = 16'h00FD; #100;
A = 16'h0073; B = 16'h00FE; #100;
A = 16'h0073; B = 16'h00FF; #100;
A = 16'h0074; B = 16'h000; #100;
A = 16'h0074; B = 16'h001; #100;
A = 16'h0074; B = 16'h002; #100;
A = 16'h0074; B = 16'h003; #100;
A = 16'h0074; B = 16'h004; #100;
A = 16'h0074; B = 16'h005; #100;
A = 16'h0074; B = 16'h006; #100;
A = 16'h0074; B = 16'h007; #100;
A = 16'h0074; B = 16'h008; #100;
A = 16'h0074; B = 16'h009; #100;
A = 16'h0074; B = 16'h00A; #100;
A = 16'h0074; B = 16'h00B; #100;
A = 16'h0074; B = 16'h00C; #100;
A = 16'h0074; B = 16'h00D; #100;
A = 16'h0074; B = 16'h00E; #100;
A = 16'h0074; B = 16'h00F; #100;
A = 16'h0074; B = 16'h0010; #100;
A = 16'h0074; B = 16'h0011; #100;
A = 16'h0074; B = 16'h0012; #100;
A = 16'h0074; B = 16'h0013; #100;
A = 16'h0074; B = 16'h0014; #100;
A = 16'h0074; B = 16'h0015; #100;
A = 16'h0074; B = 16'h0016; #100;
A = 16'h0074; B = 16'h0017; #100;
A = 16'h0074; B = 16'h0018; #100;
A = 16'h0074; B = 16'h0019; #100;
A = 16'h0074; B = 16'h001A; #100;
A = 16'h0074; B = 16'h001B; #100;
A = 16'h0074; B = 16'h001C; #100;
A = 16'h0074; B = 16'h001D; #100;
A = 16'h0074; B = 16'h001E; #100;
A = 16'h0074; B = 16'h001F; #100;
A = 16'h0074; B = 16'h0020; #100;
A = 16'h0074; B = 16'h0021; #100;
A = 16'h0074; B = 16'h0022; #100;
A = 16'h0074; B = 16'h0023; #100;
A = 16'h0074; B = 16'h0024; #100;
A = 16'h0074; B = 16'h0025; #100;
A = 16'h0074; B = 16'h0026; #100;
A = 16'h0074; B = 16'h0027; #100;
A = 16'h0074; B = 16'h0028; #100;
A = 16'h0074; B = 16'h0029; #100;
A = 16'h0074; B = 16'h002A; #100;
A = 16'h0074; B = 16'h002B; #100;
A = 16'h0074; B = 16'h002C; #100;
A = 16'h0074; B = 16'h002D; #100;
A = 16'h0074; B = 16'h002E; #100;
A = 16'h0074; B = 16'h002F; #100;
A = 16'h0074; B = 16'h0030; #100;
A = 16'h0074; B = 16'h0031; #100;
A = 16'h0074; B = 16'h0032; #100;
A = 16'h0074; B = 16'h0033; #100;
A = 16'h0074; B = 16'h0034; #100;
A = 16'h0074; B = 16'h0035; #100;
A = 16'h0074; B = 16'h0036; #100;
A = 16'h0074; B = 16'h0037; #100;
A = 16'h0074; B = 16'h0038; #100;
A = 16'h0074; B = 16'h0039; #100;
A = 16'h0074; B = 16'h003A; #100;
A = 16'h0074; B = 16'h003B; #100;
A = 16'h0074; B = 16'h003C; #100;
A = 16'h0074; B = 16'h003D; #100;
A = 16'h0074; B = 16'h003E; #100;
A = 16'h0074; B = 16'h003F; #100;
A = 16'h0074; B = 16'h0040; #100;
A = 16'h0074; B = 16'h0041; #100;
A = 16'h0074; B = 16'h0042; #100;
A = 16'h0074; B = 16'h0043; #100;
A = 16'h0074; B = 16'h0044; #100;
A = 16'h0074; B = 16'h0045; #100;
A = 16'h0074; B = 16'h0046; #100;
A = 16'h0074; B = 16'h0047; #100;
A = 16'h0074; B = 16'h0048; #100;
A = 16'h0074; B = 16'h0049; #100;
A = 16'h0074; B = 16'h004A; #100;
A = 16'h0074; B = 16'h004B; #100;
A = 16'h0074; B = 16'h004C; #100;
A = 16'h0074; B = 16'h004D; #100;
A = 16'h0074; B = 16'h004E; #100;
A = 16'h0074; B = 16'h004F; #100;
A = 16'h0074; B = 16'h0050; #100;
A = 16'h0074; B = 16'h0051; #100;
A = 16'h0074; B = 16'h0052; #100;
A = 16'h0074; B = 16'h0053; #100;
A = 16'h0074; B = 16'h0054; #100;
A = 16'h0074; B = 16'h0055; #100;
A = 16'h0074; B = 16'h0056; #100;
A = 16'h0074; B = 16'h0057; #100;
A = 16'h0074; B = 16'h0058; #100;
A = 16'h0074; B = 16'h0059; #100;
A = 16'h0074; B = 16'h005A; #100;
A = 16'h0074; B = 16'h005B; #100;
A = 16'h0074; B = 16'h005C; #100;
A = 16'h0074; B = 16'h005D; #100;
A = 16'h0074; B = 16'h005E; #100;
A = 16'h0074; B = 16'h005F; #100;
A = 16'h0074; B = 16'h0060; #100;
A = 16'h0074; B = 16'h0061; #100;
A = 16'h0074; B = 16'h0062; #100;
A = 16'h0074; B = 16'h0063; #100;
A = 16'h0074; B = 16'h0064; #100;
A = 16'h0074; B = 16'h0065; #100;
A = 16'h0074; B = 16'h0066; #100;
A = 16'h0074; B = 16'h0067; #100;
A = 16'h0074; B = 16'h0068; #100;
A = 16'h0074; B = 16'h0069; #100;
A = 16'h0074; B = 16'h006A; #100;
A = 16'h0074; B = 16'h006B; #100;
A = 16'h0074; B = 16'h006C; #100;
A = 16'h0074; B = 16'h006D; #100;
A = 16'h0074; B = 16'h006E; #100;
A = 16'h0074; B = 16'h006F; #100;
A = 16'h0074; B = 16'h0070; #100;
A = 16'h0074; B = 16'h0071; #100;
A = 16'h0074; B = 16'h0072; #100;
A = 16'h0074; B = 16'h0073; #100;
A = 16'h0074; B = 16'h0074; #100;
A = 16'h0074; B = 16'h0075; #100;
A = 16'h0074; B = 16'h0076; #100;
A = 16'h0074; B = 16'h0077; #100;
A = 16'h0074; B = 16'h0078; #100;
A = 16'h0074; B = 16'h0079; #100;
A = 16'h0074; B = 16'h007A; #100;
A = 16'h0074; B = 16'h007B; #100;
A = 16'h0074; B = 16'h007C; #100;
A = 16'h0074; B = 16'h007D; #100;
A = 16'h0074; B = 16'h007E; #100;
A = 16'h0074; B = 16'h007F; #100;
A = 16'h0074; B = 16'h0080; #100;
A = 16'h0074; B = 16'h0081; #100;
A = 16'h0074; B = 16'h0082; #100;
A = 16'h0074; B = 16'h0083; #100;
A = 16'h0074; B = 16'h0084; #100;
A = 16'h0074; B = 16'h0085; #100;
A = 16'h0074; B = 16'h0086; #100;
A = 16'h0074; B = 16'h0087; #100;
A = 16'h0074; B = 16'h0088; #100;
A = 16'h0074; B = 16'h0089; #100;
A = 16'h0074; B = 16'h008A; #100;
A = 16'h0074; B = 16'h008B; #100;
A = 16'h0074; B = 16'h008C; #100;
A = 16'h0074; B = 16'h008D; #100;
A = 16'h0074; B = 16'h008E; #100;
A = 16'h0074; B = 16'h008F; #100;
A = 16'h0074; B = 16'h0090; #100;
A = 16'h0074; B = 16'h0091; #100;
A = 16'h0074; B = 16'h0092; #100;
A = 16'h0074; B = 16'h0093; #100;
A = 16'h0074; B = 16'h0094; #100;
A = 16'h0074; B = 16'h0095; #100;
A = 16'h0074; B = 16'h0096; #100;
A = 16'h0074; B = 16'h0097; #100;
A = 16'h0074; B = 16'h0098; #100;
A = 16'h0074; B = 16'h0099; #100;
A = 16'h0074; B = 16'h009A; #100;
A = 16'h0074; B = 16'h009B; #100;
A = 16'h0074; B = 16'h009C; #100;
A = 16'h0074; B = 16'h009D; #100;
A = 16'h0074; B = 16'h009E; #100;
A = 16'h0074; B = 16'h009F; #100;
A = 16'h0074; B = 16'h00A0; #100;
A = 16'h0074; B = 16'h00A1; #100;
A = 16'h0074; B = 16'h00A2; #100;
A = 16'h0074; B = 16'h00A3; #100;
A = 16'h0074; B = 16'h00A4; #100;
A = 16'h0074; B = 16'h00A5; #100;
A = 16'h0074; B = 16'h00A6; #100;
A = 16'h0074; B = 16'h00A7; #100;
A = 16'h0074; B = 16'h00A8; #100;
A = 16'h0074; B = 16'h00A9; #100;
A = 16'h0074; B = 16'h00AA; #100;
A = 16'h0074; B = 16'h00AB; #100;
A = 16'h0074; B = 16'h00AC; #100;
A = 16'h0074; B = 16'h00AD; #100;
A = 16'h0074; B = 16'h00AE; #100;
A = 16'h0074; B = 16'h00AF; #100;
A = 16'h0074; B = 16'h00B0; #100;
A = 16'h0074; B = 16'h00B1; #100;
A = 16'h0074; B = 16'h00B2; #100;
A = 16'h0074; B = 16'h00B3; #100;
A = 16'h0074; B = 16'h00B4; #100;
A = 16'h0074; B = 16'h00B5; #100;
A = 16'h0074; B = 16'h00B6; #100;
A = 16'h0074; B = 16'h00B7; #100;
A = 16'h0074; B = 16'h00B8; #100;
A = 16'h0074; B = 16'h00B9; #100;
A = 16'h0074; B = 16'h00BA; #100;
A = 16'h0074; B = 16'h00BB; #100;
A = 16'h0074; B = 16'h00BC; #100;
A = 16'h0074; B = 16'h00BD; #100;
A = 16'h0074; B = 16'h00BE; #100;
A = 16'h0074; B = 16'h00BF; #100;
A = 16'h0074; B = 16'h00C0; #100;
A = 16'h0074; B = 16'h00C1; #100;
A = 16'h0074; B = 16'h00C2; #100;
A = 16'h0074; B = 16'h00C3; #100;
A = 16'h0074; B = 16'h00C4; #100;
A = 16'h0074; B = 16'h00C5; #100;
A = 16'h0074; B = 16'h00C6; #100;
A = 16'h0074; B = 16'h00C7; #100;
A = 16'h0074; B = 16'h00C8; #100;
A = 16'h0074; B = 16'h00C9; #100;
A = 16'h0074; B = 16'h00CA; #100;
A = 16'h0074; B = 16'h00CB; #100;
A = 16'h0074; B = 16'h00CC; #100;
A = 16'h0074; B = 16'h00CD; #100;
A = 16'h0074; B = 16'h00CE; #100;
A = 16'h0074; B = 16'h00CF; #100;
A = 16'h0074; B = 16'h00D0; #100;
A = 16'h0074; B = 16'h00D1; #100;
A = 16'h0074; B = 16'h00D2; #100;
A = 16'h0074; B = 16'h00D3; #100;
A = 16'h0074; B = 16'h00D4; #100;
A = 16'h0074; B = 16'h00D5; #100;
A = 16'h0074; B = 16'h00D6; #100;
A = 16'h0074; B = 16'h00D7; #100;
A = 16'h0074; B = 16'h00D8; #100;
A = 16'h0074; B = 16'h00D9; #100;
A = 16'h0074; B = 16'h00DA; #100;
A = 16'h0074; B = 16'h00DB; #100;
A = 16'h0074; B = 16'h00DC; #100;
A = 16'h0074; B = 16'h00DD; #100;
A = 16'h0074; B = 16'h00DE; #100;
A = 16'h0074; B = 16'h00DF; #100;
A = 16'h0074; B = 16'h00E0; #100;
A = 16'h0074; B = 16'h00E1; #100;
A = 16'h0074; B = 16'h00E2; #100;
A = 16'h0074; B = 16'h00E3; #100;
A = 16'h0074; B = 16'h00E4; #100;
A = 16'h0074; B = 16'h00E5; #100;
A = 16'h0074; B = 16'h00E6; #100;
A = 16'h0074; B = 16'h00E7; #100;
A = 16'h0074; B = 16'h00E8; #100;
A = 16'h0074; B = 16'h00E9; #100;
A = 16'h0074; B = 16'h00EA; #100;
A = 16'h0074; B = 16'h00EB; #100;
A = 16'h0074; B = 16'h00EC; #100;
A = 16'h0074; B = 16'h00ED; #100;
A = 16'h0074; B = 16'h00EE; #100;
A = 16'h0074; B = 16'h00EF; #100;
A = 16'h0074; B = 16'h00F0; #100;
A = 16'h0074; B = 16'h00F1; #100;
A = 16'h0074; B = 16'h00F2; #100;
A = 16'h0074; B = 16'h00F3; #100;
A = 16'h0074; B = 16'h00F4; #100;
A = 16'h0074; B = 16'h00F5; #100;
A = 16'h0074; B = 16'h00F6; #100;
A = 16'h0074; B = 16'h00F7; #100;
A = 16'h0074; B = 16'h00F8; #100;
A = 16'h0074; B = 16'h00F9; #100;
A = 16'h0074; B = 16'h00FA; #100;
A = 16'h0074; B = 16'h00FB; #100;
A = 16'h0074; B = 16'h00FC; #100;
A = 16'h0074; B = 16'h00FD; #100;
A = 16'h0074; B = 16'h00FE; #100;
A = 16'h0074; B = 16'h00FF; #100;
A = 16'h0075; B = 16'h000; #100;
A = 16'h0075; B = 16'h001; #100;
A = 16'h0075; B = 16'h002; #100;
A = 16'h0075; B = 16'h003; #100;
A = 16'h0075; B = 16'h004; #100;
A = 16'h0075; B = 16'h005; #100;
A = 16'h0075; B = 16'h006; #100;
A = 16'h0075; B = 16'h007; #100;
A = 16'h0075; B = 16'h008; #100;
A = 16'h0075; B = 16'h009; #100;
A = 16'h0075; B = 16'h00A; #100;
A = 16'h0075; B = 16'h00B; #100;
A = 16'h0075; B = 16'h00C; #100;
A = 16'h0075; B = 16'h00D; #100;
A = 16'h0075; B = 16'h00E; #100;
A = 16'h0075; B = 16'h00F; #100;
A = 16'h0075; B = 16'h0010; #100;
A = 16'h0075; B = 16'h0011; #100;
A = 16'h0075; B = 16'h0012; #100;
A = 16'h0075; B = 16'h0013; #100;
A = 16'h0075; B = 16'h0014; #100;
A = 16'h0075; B = 16'h0015; #100;
A = 16'h0075; B = 16'h0016; #100;
A = 16'h0075; B = 16'h0017; #100;
A = 16'h0075; B = 16'h0018; #100;
A = 16'h0075; B = 16'h0019; #100;
A = 16'h0075; B = 16'h001A; #100;
A = 16'h0075; B = 16'h001B; #100;
A = 16'h0075; B = 16'h001C; #100;
A = 16'h0075; B = 16'h001D; #100;
A = 16'h0075; B = 16'h001E; #100;
A = 16'h0075; B = 16'h001F; #100;
A = 16'h0075; B = 16'h0020; #100;
A = 16'h0075; B = 16'h0021; #100;
A = 16'h0075; B = 16'h0022; #100;
A = 16'h0075; B = 16'h0023; #100;
A = 16'h0075; B = 16'h0024; #100;
A = 16'h0075; B = 16'h0025; #100;
A = 16'h0075; B = 16'h0026; #100;
A = 16'h0075; B = 16'h0027; #100;
A = 16'h0075; B = 16'h0028; #100;
A = 16'h0075; B = 16'h0029; #100;
A = 16'h0075; B = 16'h002A; #100;
A = 16'h0075; B = 16'h002B; #100;
A = 16'h0075; B = 16'h002C; #100;
A = 16'h0075; B = 16'h002D; #100;
A = 16'h0075; B = 16'h002E; #100;
A = 16'h0075; B = 16'h002F; #100;
A = 16'h0075; B = 16'h0030; #100;
A = 16'h0075; B = 16'h0031; #100;
A = 16'h0075; B = 16'h0032; #100;
A = 16'h0075; B = 16'h0033; #100;
A = 16'h0075; B = 16'h0034; #100;
A = 16'h0075; B = 16'h0035; #100;
A = 16'h0075; B = 16'h0036; #100;
A = 16'h0075; B = 16'h0037; #100;
A = 16'h0075; B = 16'h0038; #100;
A = 16'h0075; B = 16'h0039; #100;
A = 16'h0075; B = 16'h003A; #100;
A = 16'h0075; B = 16'h003B; #100;
A = 16'h0075; B = 16'h003C; #100;
A = 16'h0075; B = 16'h003D; #100;
A = 16'h0075; B = 16'h003E; #100;
A = 16'h0075; B = 16'h003F; #100;
A = 16'h0075; B = 16'h0040; #100;
A = 16'h0075; B = 16'h0041; #100;
A = 16'h0075; B = 16'h0042; #100;
A = 16'h0075; B = 16'h0043; #100;
A = 16'h0075; B = 16'h0044; #100;
A = 16'h0075; B = 16'h0045; #100;
A = 16'h0075; B = 16'h0046; #100;
A = 16'h0075; B = 16'h0047; #100;
A = 16'h0075; B = 16'h0048; #100;
A = 16'h0075; B = 16'h0049; #100;
A = 16'h0075; B = 16'h004A; #100;
A = 16'h0075; B = 16'h004B; #100;
A = 16'h0075; B = 16'h004C; #100;
A = 16'h0075; B = 16'h004D; #100;
A = 16'h0075; B = 16'h004E; #100;
A = 16'h0075; B = 16'h004F; #100;
A = 16'h0075; B = 16'h0050; #100;
A = 16'h0075; B = 16'h0051; #100;
A = 16'h0075; B = 16'h0052; #100;
A = 16'h0075; B = 16'h0053; #100;
A = 16'h0075; B = 16'h0054; #100;
A = 16'h0075; B = 16'h0055; #100;
A = 16'h0075; B = 16'h0056; #100;
A = 16'h0075; B = 16'h0057; #100;
A = 16'h0075; B = 16'h0058; #100;
A = 16'h0075; B = 16'h0059; #100;
A = 16'h0075; B = 16'h005A; #100;
A = 16'h0075; B = 16'h005B; #100;
A = 16'h0075; B = 16'h005C; #100;
A = 16'h0075; B = 16'h005D; #100;
A = 16'h0075; B = 16'h005E; #100;
A = 16'h0075; B = 16'h005F; #100;
A = 16'h0075; B = 16'h0060; #100;
A = 16'h0075; B = 16'h0061; #100;
A = 16'h0075; B = 16'h0062; #100;
A = 16'h0075; B = 16'h0063; #100;
A = 16'h0075; B = 16'h0064; #100;
A = 16'h0075; B = 16'h0065; #100;
A = 16'h0075; B = 16'h0066; #100;
A = 16'h0075; B = 16'h0067; #100;
A = 16'h0075; B = 16'h0068; #100;
A = 16'h0075; B = 16'h0069; #100;
A = 16'h0075; B = 16'h006A; #100;
A = 16'h0075; B = 16'h006B; #100;
A = 16'h0075; B = 16'h006C; #100;
A = 16'h0075; B = 16'h006D; #100;
A = 16'h0075; B = 16'h006E; #100;
A = 16'h0075; B = 16'h006F; #100;
A = 16'h0075; B = 16'h0070; #100;
A = 16'h0075; B = 16'h0071; #100;
A = 16'h0075; B = 16'h0072; #100;
A = 16'h0075; B = 16'h0073; #100;
A = 16'h0075; B = 16'h0074; #100;
A = 16'h0075; B = 16'h0075; #100;
A = 16'h0075; B = 16'h0076; #100;
A = 16'h0075; B = 16'h0077; #100;
A = 16'h0075; B = 16'h0078; #100;
A = 16'h0075; B = 16'h0079; #100;
A = 16'h0075; B = 16'h007A; #100;
A = 16'h0075; B = 16'h007B; #100;
A = 16'h0075; B = 16'h007C; #100;
A = 16'h0075; B = 16'h007D; #100;
A = 16'h0075; B = 16'h007E; #100;
A = 16'h0075; B = 16'h007F; #100;
A = 16'h0075; B = 16'h0080; #100;
A = 16'h0075; B = 16'h0081; #100;
A = 16'h0075; B = 16'h0082; #100;
A = 16'h0075; B = 16'h0083; #100;
A = 16'h0075; B = 16'h0084; #100;
A = 16'h0075; B = 16'h0085; #100;
A = 16'h0075; B = 16'h0086; #100;
A = 16'h0075; B = 16'h0087; #100;
A = 16'h0075; B = 16'h0088; #100;
A = 16'h0075; B = 16'h0089; #100;
A = 16'h0075; B = 16'h008A; #100;
A = 16'h0075; B = 16'h008B; #100;
A = 16'h0075; B = 16'h008C; #100;
A = 16'h0075; B = 16'h008D; #100;
A = 16'h0075; B = 16'h008E; #100;
A = 16'h0075; B = 16'h008F; #100;
A = 16'h0075; B = 16'h0090; #100;
A = 16'h0075; B = 16'h0091; #100;
A = 16'h0075; B = 16'h0092; #100;
A = 16'h0075; B = 16'h0093; #100;
A = 16'h0075; B = 16'h0094; #100;
A = 16'h0075; B = 16'h0095; #100;
A = 16'h0075; B = 16'h0096; #100;
A = 16'h0075; B = 16'h0097; #100;
A = 16'h0075; B = 16'h0098; #100;
A = 16'h0075; B = 16'h0099; #100;
A = 16'h0075; B = 16'h009A; #100;
A = 16'h0075; B = 16'h009B; #100;
A = 16'h0075; B = 16'h009C; #100;
A = 16'h0075; B = 16'h009D; #100;
A = 16'h0075; B = 16'h009E; #100;
A = 16'h0075; B = 16'h009F; #100;
A = 16'h0075; B = 16'h00A0; #100;
A = 16'h0075; B = 16'h00A1; #100;
A = 16'h0075; B = 16'h00A2; #100;
A = 16'h0075; B = 16'h00A3; #100;
A = 16'h0075; B = 16'h00A4; #100;
A = 16'h0075; B = 16'h00A5; #100;
A = 16'h0075; B = 16'h00A6; #100;
A = 16'h0075; B = 16'h00A7; #100;
A = 16'h0075; B = 16'h00A8; #100;
A = 16'h0075; B = 16'h00A9; #100;
A = 16'h0075; B = 16'h00AA; #100;
A = 16'h0075; B = 16'h00AB; #100;
A = 16'h0075; B = 16'h00AC; #100;
A = 16'h0075; B = 16'h00AD; #100;
A = 16'h0075; B = 16'h00AE; #100;
A = 16'h0075; B = 16'h00AF; #100;
A = 16'h0075; B = 16'h00B0; #100;
A = 16'h0075; B = 16'h00B1; #100;
A = 16'h0075; B = 16'h00B2; #100;
A = 16'h0075; B = 16'h00B3; #100;
A = 16'h0075; B = 16'h00B4; #100;
A = 16'h0075; B = 16'h00B5; #100;
A = 16'h0075; B = 16'h00B6; #100;
A = 16'h0075; B = 16'h00B7; #100;
A = 16'h0075; B = 16'h00B8; #100;
A = 16'h0075; B = 16'h00B9; #100;
A = 16'h0075; B = 16'h00BA; #100;
A = 16'h0075; B = 16'h00BB; #100;
A = 16'h0075; B = 16'h00BC; #100;
A = 16'h0075; B = 16'h00BD; #100;
A = 16'h0075; B = 16'h00BE; #100;
A = 16'h0075; B = 16'h00BF; #100;
A = 16'h0075; B = 16'h00C0; #100;
A = 16'h0075; B = 16'h00C1; #100;
A = 16'h0075; B = 16'h00C2; #100;
A = 16'h0075; B = 16'h00C3; #100;
A = 16'h0075; B = 16'h00C4; #100;
A = 16'h0075; B = 16'h00C5; #100;
A = 16'h0075; B = 16'h00C6; #100;
A = 16'h0075; B = 16'h00C7; #100;
A = 16'h0075; B = 16'h00C8; #100;
A = 16'h0075; B = 16'h00C9; #100;
A = 16'h0075; B = 16'h00CA; #100;
A = 16'h0075; B = 16'h00CB; #100;
A = 16'h0075; B = 16'h00CC; #100;
A = 16'h0075; B = 16'h00CD; #100;
A = 16'h0075; B = 16'h00CE; #100;
A = 16'h0075; B = 16'h00CF; #100;
A = 16'h0075; B = 16'h00D0; #100;
A = 16'h0075; B = 16'h00D1; #100;
A = 16'h0075; B = 16'h00D2; #100;
A = 16'h0075; B = 16'h00D3; #100;
A = 16'h0075; B = 16'h00D4; #100;
A = 16'h0075; B = 16'h00D5; #100;
A = 16'h0075; B = 16'h00D6; #100;
A = 16'h0075; B = 16'h00D7; #100;
A = 16'h0075; B = 16'h00D8; #100;
A = 16'h0075; B = 16'h00D9; #100;
A = 16'h0075; B = 16'h00DA; #100;
A = 16'h0075; B = 16'h00DB; #100;
A = 16'h0075; B = 16'h00DC; #100;
A = 16'h0075; B = 16'h00DD; #100;
A = 16'h0075; B = 16'h00DE; #100;
A = 16'h0075; B = 16'h00DF; #100;
A = 16'h0075; B = 16'h00E0; #100;
A = 16'h0075; B = 16'h00E1; #100;
A = 16'h0075; B = 16'h00E2; #100;
A = 16'h0075; B = 16'h00E3; #100;
A = 16'h0075; B = 16'h00E4; #100;
A = 16'h0075; B = 16'h00E5; #100;
A = 16'h0075; B = 16'h00E6; #100;
A = 16'h0075; B = 16'h00E7; #100;
A = 16'h0075; B = 16'h00E8; #100;
A = 16'h0075; B = 16'h00E9; #100;
A = 16'h0075; B = 16'h00EA; #100;
A = 16'h0075; B = 16'h00EB; #100;
A = 16'h0075; B = 16'h00EC; #100;
A = 16'h0075; B = 16'h00ED; #100;
A = 16'h0075; B = 16'h00EE; #100;
A = 16'h0075; B = 16'h00EF; #100;
A = 16'h0075; B = 16'h00F0; #100;
A = 16'h0075; B = 16'h00F1; #100;
A = 16'h0075; B = 16'h00F2; #100;
A = 16'h0075; B = 16'h00F3; #100;
A = 16'h0075; B = 16'h00F4; #100;
A = 16'h0075; B = 16'h00F5; #100;
A = 16'h0075; B = 16'h00F6; #100;
A = 16'h0075; B = 16'h00F7; #100;
A = 16'h0075; B = 16'h00F8; #100;
A = 16'h0075; B = 16'h00F9; #100;
A = 16'h0075; B = 16'h00FA; #100;
A = 16'h0075; B = 16'h00FB; #100;
A = 16'h0075; B = 16'h00FC; #100;
A = 16'h0075; B = 16'h00FD; #100;
A = 16'h0075; B = 16'h00FE; #100;
A = 16'h0075; B = 16'h00FF; #100;
A = 16'h0076; B = 16'h000; #100;
A = 16'h0076; B = 16'h001; #100;
A = 16'h0076; B = 16'h002; #100;
A = 16'h0076; B = 16'h003; #100;
A = 16'h0076; B = 16'h004; #100;
A = 16'h0076; B = 16'h005; #100;
A = 16'h0076; B = 16'h006; #100;
A = 16'h0076; B = 16'h007; #100;
A = 16'h0076; B = 16'h008; #100;
A = 16'h0076; B = 16'h009; #100;
A = 16'h0076; B = 16'h00A; #100;
A = 16'h0076; B = 16'h00B; #100;
A = 16'h0076; B = 16'h00C; #100;
A = 16'h0076; B = 16'h00D; #100;
A = 16'h0076; B = 16'h00E; #100;
A = 16'h0076; B = 16'h00F; #100;
A = 16'h0076; B = 16'h0010; #100;
A = 16'h0076; B = 16'h0011; #100;
A = 16'h0076; B = 16'h0012; #100;
A = 16'h0076; B = 16'h0013; #100;
A = 16'h0076; B = 16'h0014; #100;
A = 16'h0076; B = 16'h0015; #100;
A = 16'h0076; B = 16'h0016; #100;
A = 16'h0076; B = 16'h0017; #100;
A = 16'h0076; B = 16'h0018; #100;
A = 16'h0076; B = 16'h0019; #100;
A = 16'h0076; B = 16'h001A; #100;
A = 16'h0076; B = 16'h001B; #100;
A = 16'h0076; B = 16'h001C; #100;
A = 16'h0076; B = 16'h001D; #100;
A = 16'h0076; B = 16'h001E; #100;
A = 16'h0076; B = 16'h001F; #100;
A = 16'h0076; B = 16'h0020; #100;
A = 16'h0076; B = 16'h0021; #100;
A = 16'h0076; B = 16'h0022; #100;
A = 16'h0076; B = 16'h0023; #100;
A = 16'h0076; B = 16'h0024; #100;
A = 16'h0076; B = 16'h0025; #100;
A = 16'h0076; B = 16'h0026; #100;
A = 16'h0076; B = 16'h0027; #100;
A = 16'h0076; B = 16'h0028; #100;
A = 16'h0076; B = 16'h0029; #100;
A = 16'h0076; B = 16'h002A; #100;
A = 16'h0076; B = 16'h002B; #100;
A = 16'h0076; B = 16'h002C; #100;
A = 16'h0076; B = 16'h002D; #100;
A = 16'h0076; B = 16'h002E; #100;
A = 16'h0076; B = 16'h002F; #100;
A = 16'h0076; B = 16'h0030; #100;
A = 16'h0076; B = 16'h0031; #100;
A = 16'h0076; B = 16'h0032; #100;
A = 16'h0076; B = 16'h0033; #100;
A = 16'h0076; B = 16'h0034; #100;
A = 16'h0076; B = 16'h0035; #100;
A = 16'h0076; B = 16'h0036; #100;
A = 16'h0076; B = 16'h0037; #100;
A = 16'h0076; B = 16'h0038; #100;
A = 16'h0076; B = 16'h0039; #100;
A = 16'h0076; B = 16'h003A; #100;
A = 16'h0076; B = 16'h003B; #100;
A = 16'h0076; B = 16'h003C; #100;
A = 16'h0076; B = 16'h003D; #100;
A = 16'h0076; B = 16'h003E; #100;
A = 16'h0076; B = 16'h003F; #100;
A = 16'h0076; B = 16'h0040; #100;
A = 16'h0076; B = 16'h0041; #100;
A = 16'h0076; B = 16'h0042; #100;
A = 16'h0076; B = 16'h0043; #100;
A = 16'h0076; B = 16'h0044; #100;
A = 16'h0076; B = 16'h0045; #100;
A = 16'h0076; B = 16'h0046; #100;
A = 16'h0076; B = 16'h0047; #100;
A = 16'h0076; B = 16'h0048; #100;
A = 16'h0076; B = 16'h0049; #100;
A = 16'h0076; B = 16'h004A; #100;
A = 16'h0076; B = 16'h004B; #100;
A = 16'h0076; B = 16'h004C; #100;
A = 16'h0076; B = 16'h004D; #100;
A = 16'h0076; B = 16'h004E; #100;
A = 16'h0076; B = 16'h004F; #100;
A = 16'h0076; B = 16'h0050; #100;
A = 16'h0076; B = 16'h0051; #100;
A = 16'h0076; B = 16'h0052; #100;
A = 16'h0076; B = 16'h0053; #100;
A = 16'h0076; B = 16'h0054; #100;
A = 16'h0076; B = 16'h0055; #100;
A = 16'h0076; B = 16'h0056; #100;
A = 16'h0076; B = 16'h0057; #100;
A = 16'h0076; B = 16'h0058; #100;
A = 16'h0076; B = 16'h0059; #100;
A = 16'h0076; B = 16'h005A; #100;
A = 16'h0076; B = 16'h005B; #100;
A = 16'h0076; B = 16'h005C; #100;
A = 16'h0076; B = 16'h005D; #100;
A = 16'h0076; B = 16'h005E; #100;
A = 16'h0076; B = 16'h005F; #100;
A = 16'h0076; B = 16'h0060; #100;
A = 16'h0076; B = 16'h0061; #100;
A = 16'h0076; B = 16'h0062; #100;
A = 16'h0076; B = 16'h0063; #100;
A = 16'h0076; B = 16'h0064; #100;
A = 16'h0076; B = 16'h0065; #100;
A = 16'h0076; B = 16'h0066; #100;
A = 16'h0076; B = 16'h0067; #100;
A = 16'h0076; B = 16'h0068; #100;
A = 16'h0076; B = 16'h0069; #100;
A = 16'h0076; B = 16'h006A; #100;
A = 16'h0076; B = 16'h006B; #100;
A = 16'h0076; B = 16'h006C; #100;
A = 16'h0076; B = 16'h006D; #100;
A = 16'h0076; B = 16'h006E; #100;
A = 16'h0076; B = 16'h006F; #100;
A = 16'h0076; B = 16'h0070; #100;
A = 16'h0076; B = 16'h0071; #100;
A = 16'h0076; B = 16'h0072; #100;
A = 16'h0076; B = 16'h0073; #100;
A = 16'h0076; B = 16'h0074; #100;
A = 16'h0076; B = 16'h0075; #100;
A = 16'h0076; B = 16'h0076; #100;
A = 16'h0076; B = 16'h0077; #100;
A = 16'h0076; B = 16'h0078; #100;
A = 16'h0076; B = 16'h0079; #100;
A = 16'h0076; B = 16'h007A; #100;
A = 16'h0076; B = 16'h007B; #100;
A = 16'h0076; B = 16'h007C; #100;
A = 16'h0076; B = 16'h007D; #100;
A = 16'h0076; B = 16'h007E; #100;
A = 16'h0076; B = 16'h007F; #100;
A = 16'h0076; B = 16'h0080; #100;
A = 16'h0076; B = 16'h0081; #100;
A = 16'h0076; B = 16'h0082; #100;
A = 16'h0076; B = 16'h0083; #100;
A = 16'h0076; B = 16'h0084; #100;
A = 16'h0076; B = 16'h0085; #100;
A = 16'h0076; B = 16'h0086; #100;
A = 16'h0076; B = 16'h0087; #100;
A = 16'h0076; B = 16'h0088; #100;
A = 16'h0076; B = 16'h0089; #100;
A = 16'h0076; B = 16'h008A; #100;
A = 16'h0076; B = 16'h008B; #100;
A = 16'h0076; B = 16'h008C; #100;
A = 16'h0076; B = 16'h008D; #100;
A = 16'h0076; B = 16'h008E; #100;
A = 16'h0076; B = 16'h008F; #100;
A = 16'h0076; B = 16'h0090; #100;
A = 16'h0076; B = 16'h0091; #100;
A = 16'h0076; B = 16'h0092; #100;
A = 16'h0076; B = 16'h0093; #100;
A = 16'h0076; B = 16'h0094; #100;
A = 16'h0076; B = 16'h0095; #100;
A = 16'h0076; B = 16'h0096; #100;
A = 16'h0076; B = 16'h0097; #100;
A = 16'h0076; B = 16'h0098; #100;
A = 16'h0076; B = 16'h0099; #100;
A = 16'h0076; B = 16'h009A; #100;
A = 16'h0076; B = 16'h009B; #100;
A = 16'h0076; B = 16'h009C; #100;
A = 16'h0076; B = 16'h009D; #100;
A = 16'h0076; B = 16'h009E; #100;
A = 16'h0076; B = 16'h009F; #100;
A = 16'h0076; B = 16'h00A0; #100;
A = 16'h0076; B = 16'h00A1; #100;
A = 16'h0076; B = 16'h00A2; #100;
A = 16'h0076; B = 16'h00A3; #100;
A = 16'h0076; B = 16'h00A4; #100;
A = 16'h0076; B = 16'h00A5; #100;
A = 16'h0076; B = 16'h00A6; #100;
A = 16'h0076; B = 16'h00A7; #100;
A = 16'h0076; B = 16'h00A8; #100;
A = 16'h0076; B = 16'h00A9; #100;
A = 16'h0076; B = 16'h00AA; #100;
A = 16'h0076; B = 16'h00AB; #100;
A = 16'h0076; B = 16'h00AC; #100;
A = 16'h0076; B = 16'h00AD; #100;
A = 16'h0076; B = 16'h00AE; #100;
A = 16'h0076; B = 16'h00AF; #100;
A = 16'h0076; B = 16'h00B0; #100;
A = 16'h0076; B = 16'h00B1; #100;
A = 16'h0076; B = 16'h00B2; #100;
A = 16'h0076; B = 16'h00B3; #100;
A = 16'h0076; B = 16'h00B4; #100;
A = 16'h0076; B = 16'h00B5; #100;
A = 16'h0076; B = 16'h00B6; #100;
A = 16'h0076; B = 16'h00B7; #100;
A = 16'h0076; B = 16'h00B8; #100;
A = 16'h0076; B = 16'h00B9; #100;
A = 16'h0076; B = 16'h00BA; #100;
A = 16'h0076; B = 16'h00BB; #100;
A = 16'h0076; B = 16'h00BC; #100;
A = 16'h0076; B = 16'h00BD; #100;
A = 16'h0076; B = 16'h00BE; #100;
A = 16'h0076; B = 16'h00BF; #100;
A = 16'h0076; B = 16'h00C0; #100;
A = 16'h0076; B = 16'h00C1; #100;
A = 16'h0076; B = 16'h00C2; #100;
A = 16'h0076; B = 16'h00C3; #100;
A = 16'h0076; B = 16'h00C4; #100;
A = 16'h0076; B = 16'h00C5; #100;
A = 16'h0076; B = 16'h00C6; #100;
A = 16'h0076; B = 16'h00C7; #100;
A = 16'h0076; B = 16'h00C8; #100;
A = 16'h0076; B = 16'h00C9; #100;
A = 16'h0076; B = 16'h00CA; #100;
A = 16'h0076; B = 16'h00CB; #100;
A = 16'h0076; B = 16'h00CC; #100;
A = 16'h0076; B = 16'h00CD; #100;
A = 16'h0076; B = 16'h00CE; #100;
A = 16'h0076; B = 16'h00CF; #100;
A = 16'h0076; B = 16'h00D0; #100;
A = 16'h0076; B = 16'h00D1; #100;
A = 16'h0076; B = 16'h00D2; #100;
A = 16'h0076; B = 16'h00D3; #100;
A = 16'h0076; B = 16'h00D4; #100;
A = 16'h0076; B = 16'h00D5; #100;
A = 16'h0076; B = 16'h00D6; #100;
A = 16'h0076; B = 16'h00D7; #100;
A = 16'h0076; B = 16'h00D8; #100;
A = 16'h0076; B = 16'h00D9; #100;
A = 16'h0076; B = 16'h00DA; #100;
A = 16'h0076; B = 16'h00DB; #100;
A = 16'h0076; B = 16'h00DC; #100;
A = 16'h0076; B = 16'h00DD; #100;
A = 16'h0076; B = 16'h00DE; #100;
A = 16'h0076; B = 16'h00DF; #100;
A = 16'h0076; B = 16'h00E0; #100;
A = 16'h0076; B = 16'h00E1; #100;
A = 16'h0076; B = 16'h00E2; #100;
A = 16'h0076; B = 16'h00E3; #100;
A = 16'h0076; B = 16'h00E4; #100;
A = 16'h0076; B = 16'h00E5; #100;
A = 16'h0076; B = 16'h00E6; #100;
A = 16'h0076; B = 16'h00E7; #100;
A = 16'h0076; B = 16'h00E8; #100;
A = 16'h0076; B = 16'h00E9; #100;
A = 16'h0076; B = 16'h00EA; #100;
A = 16'h0076; B = 16'h00EB; #100;
A = 16'h0076; B = 16'h00EC; #100;
A = 16'h0076; B = 16'h00ED; #100;
A = 16'h0076; B = 16'h00EE; #100;
A = 16'h0076; B = 16'h00EF; #100;
A = 16'h0076; B = 16'h00F0; #100;
A = 16'h0076; B = 16'h00F1; #100;
A = 16'h0076; B = 16'h00F2; #100;
A = 16'h0076; B = 16'h00F3; #100;
A = 16'h0076; B = 16'h00F4; #100;
A = 16'h0076; B = 16'h00F5; #100;
A = 16'h0076; B = 16'h00F6; #100;
A = 16'h0076; B = 16'h00F7; #100;
A = 16'h0076; B = 16'h00F8; #100;
A = 16'h0076; B = 16'h00F9; #100;
A = 16'h0076; B = 16'h00FA; #100;
A = 16'h0076; B = 16'h00FB; #100;
A = 16'h0076; B = 16'h00FC; #100;
A = 16'h0076; B = 16'h00FD; #100;
A = 16'h0076; B = 16'h00FE; #100;
A = 16'h0076; B = 16'h00FF; #100;
A = 16'h0077; B = 16'h000; #100;
A = 16'h0077; B = 16'h001; #100;
A = 16'h0077; B = 16'h002; #100;
A = 16'h0077; B = 16'h003; #100;
A = 16'h0077; B = 16'h004; #100;
A = 16'h0077; B = 16'h005; #100;
A = 16'h0077; B = 16'h006; #100;
A = 16'h0077; B = 16'h007; #100;
A = 16'h0077; B = 16'h008; #100;
A = 16'h0077; B = 16'h009; #100;
A = 16'h0077; B = 16'h00A; #100;
A = 16'h0077; B = 16'h00B; #100;
A = 16'h0077; B = 16'h00C; #100;
A = 16'h0077; B = 16'h00D; #100;
A = 16'h0077; B = 16'h00E; #100;
A = 16'h0077; B = 16'h00F; #100;
A = 16'h0077; B = 16'h0010; #100;
A = 16'h0077; B = 16'h0011; #100;
A = 16'h0077; B = 16'h0012; #100;
A = 16'h0077; B = 16'h0013; #100;
A = 16'h0077; B = 16'h0014; #100;
A = 16'h0077; B = 16'h0015; #100;
A = 16'h0077; B = 16'h0016; #100;
A = 16'h0077; B = 16'h0017; #100;
A = 16'h0077; B = 16'h0018; #100;
A = 16'h0077; B = 16'h0019; #100;
A = 16'h0077; B = 16'h001A; #100;
A = 16'h0077; B = 16'h001B; #100;
A = 16'h0077; B = 16'h001C; #100;
A = 16'h0077; B = 16'h001D; #100;
A = 16'h0077; B = 16'h001E; #100;
A = 16'h0077; B = 16'h001F; #100;
A = 16'h0077; B = 16'h0020; #100;
A = 16'h0077; B = 16'h0021; #100;
A = 16'h0077; B = 16'h0022; #100;
A = 16'h0077; B = 16'h0023; #100;
A = 16'h0077; B = 16'h0024; #100;
A = 16'h0077; B = 16'h0025; #100;
A = 16'h0077; B = 16'h0026; #100;
A = 16'h0077; B = 16'h0027; #100;
A = 16'h0077; B = 16'h0028; #100;
A = 16'h0077; B = 16'h0029; #100;
A = 16'h0077; B = 16'h002A; #100;
A = 16'h0077; B = 16'h002B; #100;
A = 16'h0077; B = 16'h002C; #100;
A = 16'h0077; B = 16'h002D; #100;
A = 16'h0077; B = 16'h002E; #100;
A = 16'h0077; B = 16'h002F; #100;
A = 16'h0077; B = 16'h0030; #100;
A = 16'h0077; B = 16'h0031; #100;
A = 16'h0077; B = 16'h0032; #100;
A = 16'h0077; B = 16'h0033; #100;
A = 16'h0077; B = 16'h0034; #100;
A = 16'h0077; B = 16'h0035; #100;
A = 16'h0077; B = 16'h0036; #100;
A = 16'h0077; B = 16'h0037; #100;
A = 16'h0077; B = 16'h0038; #100;
A = 16'h0077; B = 16'h0039; #100;
A = 16'h0077; B = 16'h003A; #100;
A = 16'h0077; B = 16'h003B; #100;
A = 16'h0077; B = 16'h003C; #100;
A = 16'h0077; B = 16'h003D; #100;
A = 16'h0077; B = 16'h003E; #100;
A = 16'h0077; B = 16'h003F; #100;
A = 16'h0077; B = 16'h0040; #100;
A = 16'h0077; B = 16'h0041; #100;
A = 16'h0077; B = 16'h0042; #100;
A = 16'h0077; B = 16'h0043; #100;
A = 16'h0077; B = 16'h0044; #100;
A = 16'h0077; B = 16'h0045; #100;
A = 16'h0077; B = 16'h0046; #100;
A = 16'h0077; B = 16'h0047; #100;
A = 16'h0077; B = 16'h0048; #100;
A = 16'h0077; B = 16'h0049; #100;
A = 16'h0077; B = 16'h004A; #100;
A = 16'h0077; B = 16'h004B; #100;
A = 16'h0077; B = 16'h004C; #100;
A = 16'h0077; B = 16'h004D; #100;
A = 16'h0077; B = 16'h004E; #100;
A = 16'h0077; B = 16'h004F; #100;
A = 16'h0077; B = 16'h0050; #100;
A = 16'h0077; B = 16'h0051; #100;
A = 16'h0077; B = 16'h0052; #100;
A = 16'h0077; B = 16'h0053; #100;
A = 16'h0077; B = 16'h0054; #100;
A = 16'h0077; B = 16'h0055; #100;
A = 16'h0077; B = 16'h0056; #100;
A = 16'h0077; B = 16'h0057; #100;
A = 16'h0077; B = 16'h0058; #100;
A = 16'h0077; B = 16'h0059; #100;
A = 16'h0077; B = 16'h005A; #100;
A = 16'h0077; B = 16'h005B; #100;
A = 16'h0077; B = 16'h005C; #100;
A = 16'h0077; B = 16'h005D; #100;
A = 16'h0077; B = 16'h005E; #100;
A = 16'h0077; B = 16'h005F; #100;
A = 16'h0077; B = 16'h0060; #100;
A = 16'h0077; B = 16'h0061; #100;
A = 16'h0077; B = 16'h0062; #100;
A = 16'h0077; B = 16'h0063; #100;
A = 16'h0077; B = 16'h0064; #100;
A = 16'h0077; B = 16'h0065; #100;
A = 16'h0077; B = 16'h0066; #100;
A = 16'h0077; B = 16'h0067; #100;
A = 16'h0077; B = 16'h0068; #100;
A = 16'h0077; B = 16'h0069; #100;
A = 16'h0077; B = 16'h006A; #100;
A = 16'h0077; B = 16'h006B; #100;
A = 16'h0077; B = 16'h006C; #100;
A = 16'h0077; B = 16'h006D; #100;
A = 16'h0077; B = 16'h006E; #100;
A = 16'h0077; B = 16'h006F; #100;
A = 16'h0077; B = 16'h0070; #100;
A = 16'h0077; B = 16'h0071; #100;
A = 16'h0077; B = 16'h0072; #100;
A = 16'h0077; B = 16'h0073; #100;
A = 16'h0077; B = 16'h0074; #100;
A = 16'h0077; B = 16'h0075; #100;
A = 16'h0077; B = 16'h0076; #100;
A = 16'h0077; B = 16'h0077; #100;
A = 16'h0077; B = 16'h0078; #100;
A = 16'h0077; B = 16'h0079; #100;
A = 16'h0077; B = 16'h007A; #100;
A = 16'h0077; B = 16'h007B; #100;
A = 16'h0077; B = 16'h007C; #100;
A = 16'h0077; B = 16'h007D; #100;
A = 16'h0077; B = 16'h007E; #100;
A = 16'h0077; B = 16'h007F; #100;
A = 16'h0077; B = 16'h0080; #100;
A = 16'h0077; B = 16'h0081; #100;
A = 16'h0077; B = 16'h0082; #100;
A = 16'h0077; B = 16'h0083; #100;
A = 16'h0077; B = 16'h0084; #100;
A = 16'h0077; B = 16'h0085; #100;
A = 16'h0077; B = 16'h0086; #100;
A = 16'h0077; B = 16'h0087; #100;
A = 16'h0077; B = 16'h0088; #100;
A = 16'h0077; B = 16'h0089; #100;
A = 16'h0077; B = 16'h008A; #100;
A = 16'h0077; B = 16'h008B; #100;
A = 16'h0077; B = 16'h008C; #100;
A = 16'h0077; B = 16'h008D; #100;
A = 16'h0077; B = 16'h008E; #100;
A = 16'h0077; B = 16'h008F; #100;
A = 16'h0077; B = 16'h0090; #100;
A = 16'h0077; B = 16'h0091; #100;
A = 16'h0077; B = 16'h0092; #100;
A = 16'h0077; B = 16'h0093; #100;
A = 16'h0077; B = 16'h0094; #100;
A = 16'h0077; B = 16'h0095; #100;
A = 16'h0077; B = 16'h0096; #100;
A = 16'h0077; B = 16'h0097; #100;
A = 16'h0077; B = 16'h0098; #100;
A = 16'h0077; B = 16'h0099; #100;
A = 16'h0077; B = 16'h009A; #100;
A = 16'h0077; B = 16'h009B; #100;
A = 16'h0077; B = 16'h009C; #100;
A = 16'h0077; B = 16'h009D; #100;
A = 16'h0077; B = 16'h009E; #100;
A = 16'h0077; B = 16'h009F; #100;
A = 16'h0077; B = 16'h00A0; #100;
A = 16'h0077; B = 16'h00A1; #100;
A = 16'h0077; B = 16'h00A2; #100;
A = 16'h0077; B = 16'h00A3; #100;
A = 16'h0077; B = 16'h00A4; #100;
A = 16'h0077; B = 16'h00A5; #100;
A = 16'h0077; B = 16'h00A6; #100;
A = 16'h0077; B = 16'h00A7; #100;
A = 16'h0077; B = 16'h00A8; #100;
A = 16'h0077; B = 16'h00A9; #100;
A = 16'h0077; B = 16'h00AA; #100;
A = 16'h0077; B = 16'h00AB; #100;
A = 16'h0077; B = 16'h00AC; #100;
A = 16'h0077; B = 16'h00AD; #100;
A = 16'h0077; B = 16'h00AE; #100;
A = 16'h0077; B = 16'h00AF; #100;
A = 16'h0077; B = 16'h00B0; #100;
A = 16'h0077; B = 16'h00B1; #100;
A = 16'h0077; B = 16'h00B2; #100;
A = 16'h0077; B = 16'h00B3; #100;
A = 16'h0077; B = 16'h00B4; #100;
A = 16'h0077; B = 16'h00B5; #100;
A = 16'h0077; B = 16'h00B6; #100;
A = 16'h0077; B = 16'h00B7; #100;
A = 16'h0077; B = 16'h00B8; #100;
A = 16'h0077; B = 16'h00B9; #100;
A = 16'h0077; B = 16'h00BA; #100;
A = 16'h0077; B = 16'h00BB; #100;
A = 16'h0077; B = 16'h00BC; #100;
A = 16'h0077; B = 16'h00BD; #100;
A = 16'h0077; B = 16'h00BE; #100;
A = 16'h0077; B = 16'h00BF; #100;
A = 16'h0077; B = 16'h00C0; #100;
A = 16'h0077; B = 16'h00C1; #100;
A = 16'h0077; B = 16'h00C2; #100;
A = 16'h0077; B = 16'h00C3; #100;
A = 16'h0077; B = 16'h00C4; #100;
A = 16'h0077; B = 16'h00C5; #100;
A = 16'h0077; B = 16'h00C6; #100;
A = 16'h0077; B = 16'h00C7; #100;
A = 16'h0077; B = 16'h00C8; #100;
A = 16'h0077; B = 16'h00C9; #100;
A = 16'h0077; B = 16'h00CA; #100;
A = 16'h0077; B = 16'h00CB; #100;
A = 16'h0077; B = 16'h00CC; #100;
A = 16'h0077; B = 16'h00CD; #100;
A = 16'h0077; B = 16'h00CE; #100;
A = 16'h0077; B = 16'h00CF; #100;
A = 16'h0077; B = 16'h00D0; #100;
A = 16'h0077; B = 16'h00D1; #100;
A = 16'h0077; B = 16'h00D2; #100;
A = 16'h0077; B = 16'h00D3; #100;
A = 16'h0077; B = 16'h00D4; #100;
A = 16'h0077; B = 16'h00D5; #100;
A = 16'h0077; B = 16'h00D6; #100;
A = 16'h0077; B = 16'h00D7; #100;
A = 16'h0077; B = 16'h00D8; #100;
A = 16'h0077; B = 16'h00D9; #100;
A = 16'h0077; B = 16'h00DA; #100;
A = 16'h0077; B = 16'h00DB; #100;
A = 16'h0077; B = 16'h00DC; #100;
A = 16'h0077; B = 16'h00DD; #100;
A = 16'h0077; B = 16'h00DE; #100;
A = 16'h0077; B = 16'h00DF; #100;
A = 16'h0077; B = 16'h00E0; #100;
A = 16'h0077; B = 16'h00E1; #100;
A = 16'h0077; B = 16'h00E2; #100;
A = 16'h0077; B = 16'h00E3; #100;
A = 16'h0077; B = 16'h00E4; #100;
A = 16'h0077; B = 16'h00E5; #100;
A = 16'h0077; B = 16'h00E6; #100;
A = 16'h0077; B = 16'h00E7; #100;
A = 16'h0077; B = 16'h00E8; #100;
A = 16'h0077; B = 16'h00E9; #100;
A = 16'h0077; B = 16'h00EA; #100;
A = 16'h0077; B = 16'h00EB; #100;
A = 16'h0077; B = 16'h00EC; #100;
A = 16'h0077; B = 16'h00ED; #100;
A = 16'h0077; B = 16'h00EE; #100;
A = 16'h0077; B = 16'h00EF; #100;
A = 16'h0077; B = 16'h00F0; #100;
A = 16'h0077; B = 16'h00F1; #100;
A = 16'h0077; B = 16'h00F2; #100;
A = 16'h0077; B = 16'h00F3; #100;
A = 16'h0077; B = 16'h00F4; #100;
A = 16'h0077; B = 16'h00F5; #100;
A = 16'h0077; B = 16'h00F6; #100;
A = 16'h0077; B = 16'h00F7; #100;
A = 16'h0077; B = 16'h00F8; #100;
A = 16'h0077; B = 16'h00F9; #100;
A = 16'h0077; B = 16'h00FA; #100;
A = 16'h0077; B = 16'h00FB; #100;
A = 16'h0077; B = 16'h00FC; #100;
A = 16'h0077; B = 16'h00FD; #100;
A = 16'h0077; B = 16'h00FE; #100;
A = 16'h0077; B = 16'h00FF; #100;
A = 16'h0078; B = 16'h000; #100;
A = 16'h0078; B = 16'h001; #100;
A = 16'h0078; B = 16'h002; #100;
A = 16'h0078; B = 16'h003; #100;
A = 16'h0078; B = 16'h004; #100;
A = 16'h0078; B = 16'h005; #100;
A = 16'h0078; B = 16'h006; #100;
A = 16'h0078; B = 16'h007; #100;
A = 16'h0078; B = 16'h008; #100;
A = 16'h0078; B = 16'h009; #100;
A = 16'h0078; B = 16'h00A; #100;
A = 16'h0078; B = 16'h00B; #100;
A = 16'h0078; B = 16'h00C; #100;
A = 16'h0078; B = 16'h00D; #100;
A = 16'h0078; B = 16'h00E; #100;
A = 16'h0078; B = 16'h00F; #100;
A = 16'h0078; B = 16'h0010; #100;
A = 16'h0078; B = 16'h0011; #100;
A = 16'h0078; B = 16'h0012; #100;
A = 16'h0078; B = 16'h0013; #100;
A = 16'h0078; B = 16'h0014; #100;
A = 16'h0078; B = 16'h0015; #100;
A = 16'h0078; B = 16'h0016; #100;
A = 16'h0078; B = 16'h0017; #100;
A = 16'h0078; B = 16'h0018; #100;
A = 16'h0078; B = 16'h0019; #100;
A = 16'h0078; B = 16'h001A; #100;
A = 16'h0078; B = 16'h001B; #100;
A = 16'h0078; B = 16'h001C; #100;
A = 16'h0078; B = 16'h001D; #100;
A = 16'h0078; B = 16'h001E; #100;
A = 16'h0078; B = 16'h001F; #100;
A = 16'h0078; B = 16'h0020; #100;
A = 16'h0078; B = 16'h0021; #100;
A = 16'h0078; B = 16'h0022; #100;
A = 16'h0078; B = 16'h0023; #100;
A = 16'h0078; B = 16'h0024; #100;
A = 16'h0078; B = 16'h0025; #100;
A = 16'h0078; B = 16'h0026; #100;
A = 16'h0078; B = 16'h0027; #100;
A = 16'h0078; B = 16'h0028; #100;
A = 16'h0078; B = 16'h0029; #100;
A = 16'h0078; B = 16'h002A; #100;
A = 16'h0078; B = 16'h002B; #100;
A = 16'h0078; B = 16'h002C; #100;
A = 16'h0078; B = 16'h002D; #100;
A = 16'h0078; B = 16'h002E; #100;
A = 16'h0078; B = 16'h002F; #100;
A = 16'h0078; B = 16'h0030; #100;
A = 16'h0078; B = 16'h0031; #100;
A = 16'h0078; B = 16'h0032; #100;
A = 16'h0078; B = 16'h0033; #100;
A = 16'h0078; B = 16'h0034; #100;
A = 16'h0078; B = 16'h0035; #100;
A = 16'h0078; B = 16'h0036; #100;
A = 16'h0078; B = 16'h0037; #100;
A = 16'h0078; B = 16'h0038; #100;
A = 16'h0078; B = 16'h0039; #100;
A = 16'h0078; B = 16'h003A; #100;
A = 16'h0078; B = 16'h003B; #100;
A = 16'h0078; B = 16'h003C; #100;
A = 16'h0078; B = 16'h003D; #100;
A = 16'h0078; B = 16'h003E; #100;
A = 16'h0078; B = 16'h003F; #100;
A = 16'h0078; B = 16'h0040; #100;
A = 16'h0078; B = 16'h0041; #100;
A = 16'h0078; B = 16'h0042; #100;
A = 16'h0078; B = 16'h0043; #100;
A = 16'h0078; B = 16'h0044; #100;
A = 16'h0078; B = 16'h0045; #100;
A = 16'h0078; B = 16'h0046; #100;
A = 16'h0078; B = 16'h0047; #100;
A = 16'h0078; B = 16'h0048; #100;
A = 16'h0078; B = 16'h0049; #100;
A = 16'h0078; B = 16'h004A; #100;
A = 16'h0078; B = 16'h004B; #100;
A = 16'h0078; B = 16'h004C; #100;
A = 16'h0078; B = 16'h004D; #100;
A = 16'h0078; B = 16'h004E; #100;
A = 16'h0078; B = 16'h004F; #100;
A = 16'h0078; B = 16'h0050; #100;
A = 16'h0078; B = 16'h0051; #100;
A = 16'h0078; B = 16'h0052; #100;
A = 16'h0078; B = 16'h0053; #100;
A = 16'h0078; B = 16'h0054; #100;
A = 16'h0078; B = 16'h0055; #100;
A = 16'h0078; B = 16'h0056; #100;
A = 16'h0078; B = 16'h0057; #100;
A = 16'h0078; B = 16'h0058; #100;
A = 16'h0078; B = 16'h0059; #100;
A = 16'h0078; B = 16'h005A; #100;
A = 16'h0078; B = 16'h005B; #100;
A = 16'h0078; B = 16'h005C; #100;
A = 16'h0078; B = 16'h005D; #100;
A = 16'h0078; B = 16'h005E; #100;
A = 16'h0078; B = 16'h005F; #100;
A = 16'h0078; B = 16'h0060; #100;
A = 16'h0078; B = 16'h0061; #100;
A = 16'h0078; B = 16'h0062; #100;
A = 16'h0078; B = 16'h0063; #100;
A = 16'h0078; B = 16'h0064; #100;
A = 16'h0078; B = 16'h0065; #100;
A = 16'h0078; B = 16'h0066; #100;
A = 16'h0078; B = 16'h0067; #100;
A = 16'h0078; B = 16'h0068; #100;
A = 16'h0078; B = 16'h0069; #100;
A = 16'h0078; B = 16'h006A; #100;
A = 16'h0078; B = 16'h006B; #100;
A = 16'h0078; B = 16'h006C; #100;
A = 16'h0078; B = 16'h006D; #100;
A = 16'h0078; B = 16'h006E; #100;
A = 16'h0078; B = 16'h006F; #100;
A = 16'h0078; B = 16'h0070; #100;
A = 16'h0078; B = 16'h0071; #100;
A = 16'h0078; B = 16'h0072; #100;
A = 16'h0078; B = 16'h0073; #100;
A = 16'h0078; B = 16'h0074; #100;
A = 16'h0078; B = 16'h0075; #100;
A = 16'h0078; B = 16'h0076; #100;
A = 16'h0078; B = 16'h0077; #100;
A = 16'h0078; B = 16'h0078; #100;
A = 16'h0078; B = 16'h0079; #100;
A = 16'h0078; B = 16'h007A; #100;
A = 16'h0078; B = 16'h007B; #100;
A = 16'h0078; B = 16'h007C; #100;
A = 16'h0078; B = 16'h007D; #100;
A = 16'h0078; B = 16'h007E; #100;
A = 16'h0078; B = 16'h007F; #100;
A = 16'h0078; B = 16'h0080; #100;
A = 16'h0078; B = 16'h0081; #100;
A = 16'h0078; B = 16'h0082; #100;
A = 16'h0078; B = 16'h0083; #100;
A = 16'h0078; B = 16'h0084; #100;
A = 16'h0078; B = 16'h0085; #100;
A = 16'h0078; B = 16'h0086; #100;
A = 16'h0078; B = 16'h0087; #100;
A = 16'h0078; B = 16'h0088; #100;
A = 16'h0078; B = 16'h0089; #100;
A = 16'h0078; B = 16'h008A; #100;
A = 16'h0078; B = 16'h008B; #100;
A = 16'h0078; B = 16'h008C; #100;
A = 16'h0078; B = 16'h008D; #100;
A = 16'h0078; B = 16'h008E; #100;
A = 16'h0078; B = 16'h008F; #100;
A = 16'h0078; B = 16'h0090; #100;
A = 16'h0078; B = 16'h0091; #100;
A = 16'h0078; B = 16'h0092; #100;
A = 16'h0078; B = 16'h0093; #100;
A = 16'h0078; B = 16'h0094; #100;
A = 16'h0078; B = 16'h0095; #100;
A = 16'h0078; B = 16'h0096; #100;
A = 16'h0078; B = 16'h0097; #100;
A = 16'h0078; B = 16'h0098; #100;
A = 16'h0078; B = 16'h0099; #100;
A = 16'h0078; B = 16'h009A; #100;
A = 16'h0078; B = 16'h009B; #100;
A = 16'h0078; B = 16'h009C; #100;
A = 16'h0078; B = 16'h009D; #100;
A = 16'h0078; B = 16'h009E; #100;
A = 16'h0078; B = 16'h009F; #100;
A = 16'h0078; B = 16'h00A0; #100;
A = 16'h0078; B = 16'h00A1; #100;
A = 16'h0078; B = 16'h00A2; #100;
A = 16'h0078; B = 16'h00A3; #100;
A = 16'h0078; B = 16'h00A4; #100;
A = 16'h0078; B = 16'h00A5; #100;
A = 16'h0078; B = 16'h00A6; #100;
A = 16'h0078; B = 16'h00A7; #100;
A = 16'h0078; B = 16'h00A8; #100;
A = 16'h0078; B = 16'h00A9; #100;
A = 16'h0078; B = 16'h00AA; #100;
A = 16'h0078; B = 16'h00AB; #100;
A = 16'h0078; B = 16'h00AC; #100;
A = 16'h0078; B = 16'h00AD; #100;
A = 16'h0078; B = 16'h00AE; #100;
A = 16'h0078; B = 16'h00AF; #100;
A = 16'h0078; B = 16'h00B0; #100;
A = 16'h0078; B = 16'h00B1; #100;
A = 16'h0078; B = 16'h00B2; #100;
A = 16'h0078; B = 16'h00B3; #100;
A = 16'h0078; B = 16'h00B4; #100;
A = 16'h0078; B = 16'h00B5; #100;
A = 16'h0078; B = 16'h00B6; #100;
A = 16'h0078; B = 16'h00B7; #100;
A = 16'h0078; B = 16'h00B8; #100;
A = 16'h0078; B = 16'h00B9; #100;
A = 16'h0078; B = 16'h00BA; #100;
A = 16'h0078; B = 16'h00BB; #100;
A = 16'h0078; B = 16'h00BC; #100;
A = 16'h0078; B = 16'h00BD; #100;
A = 16'h0078; B = 16'h00BE; #100;
A = 16'h0078; B = 16'h00BF; #100;
A = 16'h0078; B = 16'h00C0; #100;
A = 16'h0078; B = 16'h00C1; #100;
A = 16'h0078; B = 16'h00C2; #100;
A = 16'h0078; B = 16'h00C3; #100;
A = 16'h0078; B = 16'h00C4; #100;
A = 16'h0078; B = 16'h00C5; #100;
A = 16'h0078; B = 16'h00C6; #100;
A = 16'h0078; B = 16'h00C7; #100;
A = 16'h0078; B = 16'h00C8; #100;
A = 16'h0078; B = 16'h00C9; #100;
A = 16'h0078; B = 16'h00CA; #100;
A = 16'h0078; B = 16'h00CB; #100;
A = 16'h0078; B = 16'h00CC; #100;
A = 16'h0078; B = 16'h00CD; #100;
A = 16'h0078; B = 16'h00CE; #100;
A = 16'h0078; B = 16'h00CF; #100;
A = 16'h0078; B = 16'h00D0; #100;
A = 16'h0078; B = 16'h00D1; #100;
A = 16'h0078; B = 16'h00D2; #100;
A = 16'h0078; B = 16'h00D3; #100;
A = 16'h0078; B = 16'h00D4; #100;
A = 16'h0078; B = 16'h00D5; #100;
A = 16'h0078; B = 16'h00D6; #100;
A = 16'h0078; B = 16'h00D7; #100;
A = 16'h0078; B = 16'h00D8; #100;
A = 16'h0078; B = 16'h00D9; #100;
A = 16'h0078; B = 16'h00DA; #100;
A = 16'h0078; B = 16'h00DB; #100;
A = 16'h0078; B = 16'h00DC; #100;
A = 16'h0078; B = 16'h00DD; #100;
A = 16'h0078; B = 16'h00DE; #100;
A = 16'h0078; B = 16'h00DF; #100;
A = 16'h0078; B = 16'h00E0; #100;
A = 16'h0078; B = 16'h00E1; #100;
A = 16'h0078; B = 16'h00E2; #100;
A = 16'h0078; B = 16'h00E3; #100;
A = 16'h0078; B = 16'h00E4; #100;
A = 16'h0078; B = 16'h00E5; #100;
A = 16'h0078; B = 16'h00E6; #100;
A = 16'h0078; B = 16'h00E7; #100;
A = 16'h0078; B = 16'h00E8; #100;
A = 16'h0078; B = 16'h00E9; #100;
A = 16'h0078; B = 16'h00EA; #100;
A = 16'h0078; B = 16'h00EB; #100;
A = 16'h0078; B = 16'h00EC; #100;
A = 16'h0078; B = 16'h00ED; #100;
A = 16'h0078; B = 16'h00EE; #100;
A = 16'h0078; B = 16'h00EF; #100;
A = 16'h0078; B = 16'h00F0; #100;
A = 16'h0078; B = 16'h00F1; #100;
A = 16'h0078; B = 16'h00F2; #100;
A = 16'h0078; B = 16'h00F3; #100;
A = 16'h0078; B = 16'h00F4; #100;
A = 16'h0078; B = 16'h00F5; #100;
A = 16'h0078; B = 16'h00F6; #100;
A = 16'h0078; B = 16'h00F7; #100;
A = 16'h0078; B = 16'h00F8; #100;
A = 16'h0078; B = 16'h00F9; #100;
A = 16'h0078; B = 16'h00FA; #100;
A = 16'h0078; B = 16'h00FB; #100;
A = 16'h0078; B = 16'h00FC; #100;
A = 16'h0078; B = 16'h00FD; #100;
A = 16'h0078; B = 16'h00FE; #100;
A = 16'h0078; B = 16'h00FF; #100;
A = 16'h0079; B = 16'h000; #100;
A = 16'h0079; B = 16'h001; #100;
A = 16'h0079; B = 16'h002; #100;
A = 16'h0079; B = 16'h003; #100;
A = 16'h0079; B = 16'h004; #100;
A = 16'h0079; B = 16'h005; #100;
A = 16'h0079; B = 16'h006; #100;
A = 16'h0079; B = 16'h007; #100;
A = 16'h0079; B = 16'h008; #100;
A = 16'h0079; B = 16'h009; #100;
A = 16'h0079; B = 16'h00A; #100;
A = 16'h0079; B = 16'h00B; #100;
A = 16'h0079; B = 16'h00C; #100;
A = 16'h0079; B = 16'h00D; #100;
A = 16'h0079; B = 16'h00E; #100;
A = 16'h0079; B = 16'h00F; #100;
A = 16'h0079; B = 16'h0010; #100;
A = 16'h0079; B = 16'h0011; #100;
A = 16'h0079; B = 16'h0012; #100;
A = 16'h0079; B = 16'h0013; #100;
A = 16'h0079; B = 16'h0014; #100;
A = 16'h0079; B = 16'h0015; #100;
A = 16'h0079; B = 16'h0016; #100;
A = 16'h0079; B = 16'h0017; #100;
A = 16'h0079; B = 16'h0018; #100;
A = 16'h0079; B = 16'h0019; #100;
A = 16'h0079; B = 16'h001A; #100;
A = 16'h0079; B = 16'h001B; #100;
A = 16'h0079; B = 16'h001C; #100;
A = 16'h0079; B = 16'h001D; #100;
A = 16'h0079; B = 16'h001E; #100;
A = 16'h0079; B = 16'h001F; #100;
A = 16'h0079; B = 16'h0020; #100;
A = 16'h0079; B = 16'h0021; #100;
A = 16'h0079; B = 16'h0022; #100;
A = 16'h0079; B = 16'h0023; #100;
A = 16'h0079; B = 16'h0024; #100;
A = 16'h0079; B = 16'h0025; #100;
A = 16'h0079; B = 16'h0026; #100;
A = 16'h0079; B = 16'h0027; #100;
A = 16'h0079; B = 16'h0028; #100;
A = 16'h0079; B = 16'h0029; #100;
A = 16'h0079; B = 16'h002A; #100;
A = 16'h0079; B = 16'h002B; #100;
A = 16'h0079; B = 16'h002C; #100;
A = 16'h0079; B = 16'h002D; #100;
A = 16'h0079; B = 16'h002E; #100;
A = 16'h0079; B = 16'h002F; #100;
A = 16'h0079; B = 16'h0030; #100;
A = 16'h0079; B = 16'h0031; #100;
A = 16'h0079; B = 16'h0032; #100;
A = 16'h0079; B = 16'h0033; #100;
A = 16'h0079; B = 16'h0034; #100;
A = 16'h0079; B = 16'h0035; #100;
A = 16'h0079; B = 16'h0036; #100;
A = 16'h0079; B = 16'h0037; #100;
A = 16'h0079; B = 16'h0038; #100;
A = 16'h0079; B = 16'h0039; #100;
A = 16'h0079; B = 16'h003A; #100;
A = 16'h0079; B = 16'h003B; #100;
A = 16'h0079; B = 16'h003C; #100;
A = 16'h0079; B = 16'h003D; #100;
A = 16'h0079; B = 16'h003E; #100;
A = 16'h0079; B = 16'h003F; #100;
A = 16'h0079; B = 16'h0040; #100;
A = 16'h0079; B = 16'h0041; #100;
A = 16'h0079; B = 16'h0042; #100;
A = 16'h0079; B = 16'h0043; #100;
A = 16'h0079; B = 16'h0044; #100;
A = 16'h0079; B = 16'h0045; #100;
A = 16'h0079; B = 16'h0046; #100;
A = 16'h0079; B = 16'h0047; #100;
A = 16'h0079; B = 16'h0048; #100;
A = 16'h0079; B = 16'h0049; #100;
A = 16'h0079; B = 16'h004A; #100;
A = 16'h0079; B = 16'h004B; #100;
A = 16'h0079; B = 16'h004C; #100;
A = 16'h0079; B = 16'h004D; #100;
A = 16'h0079; B = 16'h004E; #100;
A = 16'h0079; B = 16'h004F; #100;
A = 16'h0079; B = 16'h0050; #100;
A = 16'h0079; B = 16'h0051; #100;
A = 16'h0079; B = 16'h0052; #100;
A = 16'h0079; B = 16'h0053; #100;
A = 16'h0079; B = 16'h0054; #100;
A = 16'h0079; B = 16'h0055; #100;
A = 16'h0079; B = 16'h0056; #100;
A = 16'h0079; B = 16'h0057; #100;
A = 16'h0079; B = 16'h0058; #100;
A = 16'h0079; B = 16'h0059; #100;
A = 16'h0079; B = 16'h005A; #100;
A = 16'h0079; B = 16'h005B; #100;
A = 16'h0079; B = 16'h005C; #100;
A = 16'h0079; B = 16'h005D; #100;
A = 16'h0079; B = 16'h005E; #100;
A = 16'h0079; B = 16'h005F; #100;
A = 16'h0079; B = 16'h0060; #100;
A = 16'h0079; B = 16'h0061; #100;
A = 16'h0079; B = 16'h0062; #100;
A = 16'h0079; B = 16'h0063; #100;
A = 16'h0079; B = 16'h0064; #100;
A = 16'h0079; B = 16'h0065; #100;
A = 16'h0079; B = 16'h0066; #100;
A = 16'h0079; B = 16'h0067; #100;
A = 16'h0079; B = 16'h0068; #100;
A = 16'h0079; B = 16'h0069; #100;
A = 16'h0079; B = 16'h006A; #100;
A = 16'h0079; B = 16'h006B; #100;
A = 16'h0079; B = 16'h006C; #100;
A = 16'h0079; B = 16'h006D; #100;
A = 16'h0079; B = 16'h006E; #100;
A = 16'h0079; B = 16'h006F; #100;
A = 16'h0079; B = 16'h0070; #100;
A = 16'h0079; B = 16'h0071; #100;
A = 16'h0079; B = 16'h0072; #100;
A = 16'h0079; B = 16'h0073; #100;
A = 16'h0079; B = 16'h0074; #100;
A = 16'h0079; B = 16'h0075; #100;
A = 16'h0079; B = 16'h0076; #100;
A = 16'h0079; B = 16'h0077; #100;
A = 16'h0079; B = 16'h0078; #100;
A = 16'h0079; B = 16'h0079; #100;
A = 16'h0079; B = 16'h007A; #100;
A = 16'h0079; B = 16'h007B; #100;
A = 16'h0079; B = 16'h007C; #100;
A = 16'h0079; B = 16'h007D; #100;
A = 16'h0079; B = 16'h007E; #100;
A = 16'h0079; B = 16'h007F; #100;
A = 16'h0079; B = 16'h0080; #100;
A = 16'h0079; B = 16'h0081; #100;
A = 16'h0079; B = 16'h0082; #100;
A = 16'h0079; B = 16'h0083; #100;
A = 16'h0079; B = 16'h0084; #100;
A = 16'h0079; B = 16'h0085; #100;
A = 16'h0079; B = 16'h0086; #100;
A = 16'h0079; B = 16'h0087; #100;
A = 16'h0079; B = 16'h0088; #100;
A = 16'h0079; B = 16'h0089; #100;
A = 16'h0079; B = 16'h008A; #100;
A = 16'h0079; B = 16'h008B; #100;
A = 16'h0079; B = 16'h008C; #100;
A = 16'h0079; B = 16'h008D; #100;
A = 16'h0079; B = 16'h008E; #100;
A = 16'h0079; B = 16'h008F; #100;
A = 16'h0079; B = 16'h0090; #100;
A = 16'h0079; B = 16'h0091; #100;
A = 16'h0079; B = 16'h0092; #100;
A = 16'h0079; B = 16'h0093; #100;
A = 16'h0079; B = 16'h0094; #100;
A = 16'h0079; B = 16'h0095; #100;
A = 16'h0079; B = 16'h0096; #100;
A = 16'h0079; B = 16'h0097; #100;
A = 16'h0079; B = 16'h0098; #100;
A = 16'h0079; B = 16'h0099; #100;
A = 16'h0079; B = 16'h009A; #100;
A = 16'h0079; B = 16'h009B; #100;
A = 16'h0079; B = 16'h009C; #100;
A = 16'h0079; B = 16'h009D; #100;
A = 16'h0079; B = 16'h009E; #100;
A = 16'h0079; B = 16'h009F; #100;
A = 16'h0079; B = 16'h00A0; #100;
A = 16'h0079; B = 16'h00A1; #100;
A = 16'h0079; B = 16'h00A2; #100;
A = 16'h0079; B = 16'h00A3; #100;
A = 16'h0079; B = 16'h00A4; #100;
A = 16'h0079; B = 16'h00A5; #100;
A = 16'h0079; B = 16'h00A6; #100;
A = 16'h0079; B = 16'h00A7; #100;
A = 16'h0079; B = 16'h00A8; #100;
A = 16'h0079; B = 16'h00A9; #100;
A = 16'h0079; B = 16'h00AA; #100;
A = 16'h0079; B = 16'h00AB; #100;
A = 16'h0079; B = 16'h00AC; #100;
A = 16'h0079; B = 16'h00AD; #100;
A = 16'h0079; B = 16'h00AE; #100;
A = 16'h0079; B = 16'h00AF; #100;
A = 16'h0079; B = 16'h00B0; #100;
A = 16'h0079; B = 16'h00B1; #100;
A = 16'h0079; B = 16'h00B2; #100;
A = 16'h0079; B = 16'h00B3; #100;
A = 16'h0079; B = 16'h00B4; #100;
A = 16'h0079; B = 16'h00B5; #100;
A = 16'h0079; B = 16'h00B6; #100;
A = 16'h0079; B = 16'h00B7; #100;
A = 16'h0079; B = 16'h00B8; #100;
A = 16'h0079; B = 16'h00B9; #100;
A = 16'h0079; B = 16'h00BA; #100;
A = 16'h0079; B = 16'h00BB; #100;
A = 16'h0079; B = 16'h00BC; #100;
A = 16'h0079; B = 16'h00BD; #100;
A = 16'h0079; B = 16'h00BE; #100;
A = 16'h0079; B = 16'h00BF; #100;
A = 16'h0079; B = 16'h00C0; #100;
A = 16'h0079; B = 16'h00C1; #100;
A = 16'h0079; B = 16'h00C2; #100;
A = 16'h0079; B = 16'h00C3; #100;
A = 16'h0079; B = 16'h00C4; #100;
A = 16'h0079; B = 16'h00C5; #100;
A = 16'h0079; B = 16'h00C6; #100;
A = 16'h0079; B = 16'h00C7; #100;
A = 16'h0079; B = 16'h00C8; #100;
A = 16'h0079; B = 16'h00C9; #100;
A = 16'h0079; B = 16'h00CA; #100;
A = 16'h0079; B = 16'h00CB; #100;
A = 16'h0079; B = 16'h00CC; #100;
A = 16'h0079; B = 16'h00CD; #100;
A = 16'h0079; B = 16'h00CE; #100;
A = 16'h0079; B = 16'h00CF; #100;
A = 16'h0079; B = 16'h00D0; #100;
A = 16'h0079; B = 16'h00D1; #100;
A = 16'h0079; B = 16'h00D2; #100;
A = 16'h0079; B = 16'h00D3; #100;
A = 16'h0079; B = 16'h00D4; #100;
A = 16'h0079; B = 16'h00D5; #100;
A = 16'h0079; B = 16'h00D6; #100;
A = 16'h0079; B = 16'h00D7; #100;
A = 16'h0079; B = 16'h00D8; #100;
A = 16'h0079; B = 16'h00D9; #100;
A = 16'h0079; B = 16'h00DA; #100;
A = 16'h0079; B = 16'h00DB; #100;
A = 16'h0079; B = 16'h00DC; #100;
A = 16'h0079; B = 16'h00DD; #100;
A = 16'h0079; B = 16'h00DE; #100;
A = 16'h0079; B = 16'h00DF; #100;
A = 16'h0079; B = 16'h00E0; #100;
A = 16'h0079; B = 16'h00E1; #100;
A = 16'h0079; B = 16'h00E2; #100;
A = 16'h0079; B = 16'h00E3; #100;
A = 16'h0079; B = 16'h00E4; #100;
A = 16'h0079; B = 16'h00E5; #100;
A = 16'h0079; B = 16'h00E6; #100;
A = 16'h0079; B = 16'h00E7; #100;
A = 16'h0079; B = 16'h00E8; #100;
A = 16'h0079; B = 16'h00E9; #100;
A = 16'h0079; B = 16'h00EA; #100;
A = 16'h0079; B = 16'h00EB; #100;
A = 16'h0079; B = 16'h00EC; #100;
A = 16'h0079; B = 16'h00ED; #100;
A = 16'h0079; B = 16'h00EE; #100;
A = 16'h0079; B = 16'h00EF; #100;
A = 16'h0079; B = 16'h00F0; #100;
A = 16'h0079; B = 16'h00F1; #100;
A = 16'h0079; B = 16'h00F2; #100;
A = 16'h0079; B = 16'h00F3; #100;
A = 16'h0079; B = 16'h00F4; #100;
A = 16'h0079; B = 16'h00F5; #100;
A = 16'h0079; B = 16'h00F6; #100;
A = 16'h0079; B = 16'h00F7; #100;
A = 16'h0079; B = 16'h00F8; #100;
A = 16'h0079; B = 16'h00F9; #100;
A = 16'h0079; B = 16'h00FA; #100;
A = 16'h0079; B = 16'h00FB; #100;
A = 16'h0079; B = 16'h00FC; #100;
A = 16'h0079; B = 16'h00FD; #100;
A = 16'h0079; B = 16'h00FE; #100;
A = 16'h0079; B = 16'h00FF; #100;
A = 16'h007A; B = 16'h000; #100;
A = 16'h007A; B = 16'h001; #100;
A = 16'h007A; B = 16'h002; #100;
A = 16'h007A; B = 16'h003; #100;
A = 16'h007A; B = 16'h004; #100;
A = 16'h007A; B = 16'h005; #100;
A = 16'h007A; B = 16'h006; #100;
A = 16'h007A; B = 16'h007; #100;
A = 16'h007A; B = 16'h008; #100;
A = 16'h007A; B = 16'h009; #100;
A = 16'h007A; B = 16'h00A; #100;
A = 16'h007A; B = 16'h00B; #100;
A = 16'h007A; B = 16'h00C; #100;
A = 16'h007A; B = 16'h00D; #100;
A = 16'h007A; B = 16'h00E; #100;
A = 16'h007A; B = 16'h00F; #100;
A = 16'h007A; B = 16'h0010; #100;
A = 16'h007A; B = 16'h0011; #100;
A = 16'h007A; B = 16'h0012; #100;
A = 16'h007A; B = 16'h0013; #100;
A = 16'h007A; B = 16'h0014; #100;
A = 16'h007A; B = 16'h0015; #100;
A = 16'h007A; B = 16'h0016; #100;
A = 16'h007A; B = 16'h0017; #100;
A = 16'h007A; B = 16'h0018; #100;
A = 16'h007A; B = 16'h0019; #100;
A = 16'h007A; B = 16'h001A; #100;
A = 16'h007A; B = 16'h001B; #100;
A = 16'h007A; B = 16'h001C; #100;
A = 16'h007A; B = 16'h001D; #100;
A = 16'h007A; B = 16'h001E; #100;
A = 16'h007A; B = 16'h001F; #100;
A = 16'h007A; B = 16'h0020; #100;
A = 16'h007A; B = 16'h0021; #100;
A = 16'h007A; B = 16'h0022; #100;
A = 16'h007A; B = 16'h0023; #100;
A = 16'h007A; B = 16'h0024; #100;
A = 16'h007A; B = 16'h0025; #100;
A = 16'h007A; B = 16'h0026; #100;
A = 16'h007A; B = 16'h0027; #100;
A = 16'h007A; B = 16'h0028; #100;
A = 16'h007A; B = 16'h0029; #100;
A = 16'h007A; B = 16'h002A; #100;
A = 16'h007A; B = 16'h002B; #100;
A = 16'h007A; B = 16'h002C; #100;
A = 16'h007A; B = 16'h002D; #100;
A = 16'h007A; B = 16'h002E; #100;
A = 16'h007A; B = 16'h002F; #100;
A = 16'h007A; B = 16'h0030; #100;
A = 16'h007A; B = 16'h0031; #100;
A = 16'h007A; B = 16'h0032; #100;
A = 16'h007A; B = 16'h0033; #100;
A = 16'h007A; B = 16'h0034; #100;
A = 16'h007A; B = 16'h0035; #100;
A = 16'h007A; B = 16'h0036; #100;
A = 16'h007A; B = 16'h0037; #100;
A = 16'h007A; B = 16'h0038; #100;
A = 16'h007A; B = 16'h0039; #100;
A = 16'h007A; B = 16'h003A; #100;
A = 16'h007A; B = 16'h003B; #100;
A = 16'h007A; B = 16'h003C; #100;
A = 16'h007A; B = 16'h003D; #100;
A = 16'h007A; B = 16'h003E; #100;
A = 16'h007A; B = 16'h003F; #100;
A = 16'h007A; B = 16'h0040; #100;
A = 16'h007A; B = 16'h0041; #100;
A = 16'h007A; B = 16'h0042; #100;
A = 16'h007A; B = 16'h0043; #100;
A = 16'h007A; B = 16'h0044; #100;
A = 16'h007A; B = 16'h0045; #100;
A = 16'h007A; B = 16'h0046; #100;
A = 16'h007A; B = 16'h0047; #100;
A = 16'h007A; B = 16'h0048; #100;
A = 16'h007A; B = 16'h0049; #100;
A = 16'h007A; B = 16'h004A; #100;
A = 16'h007A; B = 16'h004B; #100;
A = 16'h007A; B = 16'h004C; #100;
A = 16'h007A; B = 16'h004D; #100;
A = 16'h007A; B = 16'h004E; #100;
A = 16'h007A; B = 16'h004F; #100;
A = 16'h007A; B = 16'h0050; #100;
A = 16'h007A; B = 16'h0051; #100;
A = 16'h007A; B = 16'h0052; #100;
A = 16'h007A; B = 16'h0053; #100;
A = 16'h007A; B = 16'h0054; #100;
A = 16'h007A; B = 16'h0055; #100;
A = 16'h007A; B = 16'h0056; #100;
A = 16'h007A; B = 16'h0057; #100;
A = 16'h007A; B = 16'h0058; #100;
A = 16'h007A; B = 16'h0059; #100;
A = 16'h007A; B = 16'h005A; #100;
A = 16'h007A; B = 16'h005B; #100;
A = 16'h007A; B = 16'h005C; #100;
A = 16'h007A; B = 16'h005D; #100;
A = 16'h007A; B = 16'h005E; #100;
A = 16'h007A; B = 16'h005F; #100;
A = 16'h007A; B = 16'h0060; #100;
A = 16'h007A; B = 16'h0061; #100;
A = 16'h007A; B = 16'h0062; #100;
A = 16'h007A; B = 16'h0063; #100;
A = 16'h007A; B = 16'h0064; #100;
A = 16'h007A; B = 16'h0065; #100;
A = 16'h007A; B = 16'h0066; #100;
A = 16'h007A; B = 16'h0067; #100;
A = 16'h007A; B = 16'h0068; #100;
A = 16'h007A; B = 16'h0069; #100;
A = 16'h007A; B = 16'h006A; #100;
A = 16'h007A; B = 16'h006B; #100;
A = 16'h007A; B = 16'h006C; #100;
A = 16'h007A; B = 16'h006D; #100;
A = 16'h007A; B = 16'h006E; #100;
A = 16'h007A; B = 16'h006F; #100;
A = 16'h007A; B = 16'h0070; #100;
A = 16'h007A; B = 16'h0071; #100;
A = 16'h007A; B = 16'h0072; #100;
A = 16'h007A; B = 16'h0073; #100;
A = 16'h007A; B = 16'h0074; #100;
A = 16'h007A; B = 16'h0075; #100;
A = 16'h007A; B = 16'h0076; #100;
A = 16'h007A; B = 16'h0077; #100;
A = 16'h007A; B = 16'h0078; #100;
A = 16'h007A; B = 16'h0079; #100;
A = 16'h007A; B = 16'h007A; #100;
A = 16'h007A; B = 16'h007B; #100;
A = 16'h007A; B = 16'h007C; #100;
A = 16'h007A; B = 16'h007D; #100;
A = 16'h007A; B = 16'h007E; #100;
A = 16'h007A; B = 16'h007F; #100;
A = 16'h007A; B = 16'h0080; #100;
A = 16'h007A; B = 16'h0081; #100;
A = 16'h007A; B = 16'h0082; #100;
A = 16'h007A; B = 16'h0083; #100;
A = 16'h007A; B = 16'h0084; #100;
A = 16'h007A; B = 16'h0085; #100;
A = 16'h007A; B = 16'h0086; #100;
A = 16'h007A; B = 16'h0087; #100;
A = 16'h007A; B = 16'h0088; #100;
A = 16'h007A; B = 16'h0089; #100;
A = 16'h007A; B = 16'h008A; #100;
A = 16'h007A; B = 16'h008B; #100;
A = 16'h007A; B = 16'h008C; #100;
A = 16'h007A; B = 16'h008D; #100;
A = 16'h007A; B = 16'h008E; #100;
A = 16'h007A; B = 16'h008F; #100;
A = 16'h007A; B = 16'h0090; #100;
A = 16'h007A; B = 16'h0091; #100;
A = 16'h007A; B = 16'h0092; #100;
A = 16'h007A; B = 16'h0093; #100;
A = 16'h007A; B = 16'h0094; #100;
A = 16'h007A; B = 16'h0095; #100;
A = 16'h007A; B = 16'h0096; #100;
A = 16'h007A; B = 16'h0097; #100;
A = 16'h007A; B = 16'h0098; #100;
A = 16'h007A; B = 16'h0099; #100;
A = 16'h007A; B = 16'h009A; #100;
A = 16'h007A; B = 16'h009B; #100;
A = 16'h007A; B = 16'h009C; #100;
A = 16'h007A; B = 16'h009D; #100;
A = 16'h007A; B = 16'h009E; #100;
A = 16'h007A; B = 16'h009F; #100;
A = 16'h007A; B = 16'h00A0; #100;
A = 16'h007A; B = 16'h00A1; #100;
A = 16'h007A; B = 16'h00A2; #100;
A = 16'h007A; B = 16'h00A3; #100;
A = 16'h007A; B = 16'h00A4; #100;
A = 16'h007A; B = 16'h00A5; #100;
A = 16'h007A; B = 16'h00A6; #100;
A = 16'h007A; B = 16'h00A7; #100;
A = 16'h007A; B = 16'h00A8; #100;
A = 16'h007A; B = 16'h00A9; #100;
A = 16'h007A; B = 16'h00AA; #100;
A = 16'h007A; B = 16'h00AB; #100;
A = 16'h007A; B = 16'h00AC; #100;
A = 16'h007A; B = 16'h00AD; #100;
A = 16'h007A; B = 16'h00AE; #100;
A = 16'h007A; B = 16'h00AF; #100;
A = 16'h007A; B = 16'h00B0; #100;
A = 16'h007A; B = 16'h00B1; #100;
A = 16'h007A; B = 16'h00B2; #100;
A = 16'h007A; B = 16'h00B3; #100;
A = 16'h007A; B = 16'h00B4; #100;
A = 16'h007A; B = 16'h00B5; #100;
A = 16'h007A; B = 16'h00B6; #100;
A = 16'h007A; B = 16'h00B7; #100;
A = 16'h007A; B = 16'h00B8; #100;
A = 16'h007A; B = 16'h00B9; #100;
A = 16'h007A; B = 16'h00BA; #100;
A = 16'h007A; B = 16'h00BB; #100;
A = 16'h007A; B = 16'h00BC; #100;
A = 16'h007A; B = 16'h00BD; #100;
A = 16'h007A; B = 16'h00BE; #100;
A = 16'h007A; B = 16'h00BF; #100;
A = 16'h007A; B = 16'h00C0; #100;
A = 16'h007A; B = 16'h00C1; #100;
A = 16'h007A; B = 16'h00C2; #100;
A = 16'h007A; B = 16'h00C3; #100;
A = 16'h007A; B = 16'h00C4; #100;
A = 16'h007A; B = 16'h00C5; #100;
A = 16'h007A; B = 16'h00C6; #100;
A = 16'h007A; B = 16'h00C7; #100;
A = 16'h007A; B = 16'h00C8; #100;
A = 16'h007A; B = 16'h00C9; #100;
A = 16'h007A; B = 16'h00CA; #100;
A = 16'h007A; B = 16'h00CB; #100;
A = 16'h007A; B = 16'h00CC; #100;
A = 16'h007A; B = 16'h00CD; #100;
A = 16'h007A; B = 16'h00CE; #100;
A = 16'h007A; B = 16'h00CF; #100;
A = 16'h007A; B = 16'h00D0; #100;
A = 16'h007A; B = 16'h00D1; #100;
A = 16'h007A; B = 16'h00D2; #100;
A = 16'h007A; B = 16'h00D3; #100;
A = 16'h007A; B = 16'h00D4; #100;
A = 16'h007A; B = 16'h00D5; #100;
A = 16'h007A; B = 16'h00D6; #100;
A = 16'h007A; B = 16'h00D7; #100;
A = 16'h007A; B = 16'h00D8; #100;
A = 16'h007A; B = 16'h00D9; #100;
A = 16'h007A; B = 16'h00DA; #100;
A = 16'h007A; B = 16'h00DB; #100;
A = 16'h007A; B = 16'h00DC; #100;
A = 16'h007A; B = 16'h00DD; #100;
A = 16'h007A; B = 16'h00DE; #100;
A = 16'h007A; B = 16'h00DF; #100;
A = 16'h007A; B = 16'h00E0; #100;
A = 16'h007A; B = 16'h00E1; #100;
A = 16'h007A; B = 16'h00E2; #100;
A = 16'h007A; B = 16'h00E3; #100;
A = 16'h007A; B = 16'h00E4; #100;
A = 16'h007A; B = 16'h00E5; #100;
A = 16'h007A; B = 16'h00E6; #100;
A = 16'h007A; B = 16'h00E7; #100;
A = 16'h007A; B = 16'h00E8; #100;
A = 16'h007A; B = 16'h00E9; #100;
A = 16'h007A; B = 16'h00EA; #100;
A = 16'h007A; B = 16'h00EB; #100;
A = 16'h007A; B = 16'h00EC; #100;
A = 16'h007A; B = 16'h00ED; #100;
A = 16'h007A; B = 16'h00EE; #100;
A = 16'h007A; B = 16'h00EF; #100;
A = 16'h007A; B = 16'h00F0; #100;
A = 16'h007A; B = 16'h00F1; #100;
A = 16'h007A; B = 16'h00F2; #100;
A = 16'h007A; B = 16'h00F3; #100;
A = 16'h007A; B = 16'h00F4; #100;
A = 16'h007A; B = 16'h00F5; #100;
A = 16'h007A; B = 16'h00F6; #100;
A = 16'h007A; B = 16'h00F7; #100;
A = 16'h007A; B = 16'h00F8; #100;
A = 16'h007A; B = 16'h00F9; #100;
A = 16'h007A; B = 16'h00FA; #100;
A = 16'h007A; B = 16'h00FB; #100;
A = 16'h007A; B = 16'h00FC; #100;
A = 16'h007A; B = 16'h00FD; #100;
A = 16'h007A; B = 16'h00FE; #100;
A = 16'h007A; B = 16'h00FF; #100;
A = 16'h007B; B = 16'h000; #100;
A = 16'h007B; B = 16'h001; #100;
A = 16'h007B; B = 16'h002; #100;
A = 16'h007B; B = 16'h003; #100;
A = 16'h007B; B = 16'h004; #100;
A = 16'h007B; B = 16'h005; #100;
A = 16'h007B; B = 16'h006; #100;
A = 16'h007B; B = 16'h007; #100;
A = 16'h007B; B = 16'h008; #100;
A = 16'h007B; B = 16'h009; #100;
A = 16'h007B; B = 16'h00A; #100;
A = 16'h007B; B = 16'h00B; #100;
A = 16'h007B; B = 16'h00C; #100;
A = 16'h007B; B = 16'h00D; #100;
A = 16'h007B; B = 16'h00E; #100;
A = 16'h007B; B = 16'h00F; #100;
A = 16'h007B; B = 16'h0010; #100;
A = 16'h007B; B = 16'h0011; #100;
A = 16'h007B; B = 16'h0012; #100;
A = 16'h007B; B = 16'h0013; #100;
A = 16'h007B; B = 16'h0014; #100;
A = 16'h007B; B = 16'h0015; #100;
A = 16'h007B; B = 16'h0016; #100;
A = 16'h007B; B = 16'h0017; #100;
A = 16'h007B; B = 16'h0018; #100;
A = 16'h007B; B = 16'h0019; #100;
A = 16'h007B; B = 16'h001A; #100;
A = 16'h007B; B = 16'h001B; #100;
A = 16'h007B; B = 16'h001C; #100;
A = 16'h007B; B = 16'h001D; #100;
A = 16'h007B; B = 16'h001E; #100;
A = 16'h007B; B = 16'h001F; #100;
A = 16'h007B; B = 16'h0020; #100;
A = 16'h007B; B = 16'h0021; #100;
A = 16'h007B; B = 16'h0022; #100;
A = 16'h007B; B = 16'h0023; #100;
A = 16'h007B; B = 16'h0024; #100;
A = 16'h007B; B = 16'h0025; #100;
A = 16'h007B; B = 16'h0026; #100;
A = 16'h007B; B = 16'h0027; #100;
A = 16'h007B; B = 16'h0028; #100;
A = 16'h007B; B = 16'h0029; #100;
A = 16'h007B; B = 16'h002A; #100;
A = 16'h007B; B = 16'h002B; #100;
A = 16'h007B; B = 16'h002C; #100;
A = 16'h007B; B = 16'h002D; #100;
A = 16'h007B; B = 16'h002E; #100;
A = 16'h007B; B = 16'h002F; #100;
A = 16'h007B; B = 16'h0030; #100;
A = 16'h007B; B = 16'h0031; #100;
A = 16'h007B; B = 16'h0032; #100;
A = 16'h007B; B = 16'h0033; #100;
A = 16'h007B; B = 16'h0034; #100;
A = 16'h007B; B = 16'h0035; #100;
A = 16'h007B; B = 16'h0036; #100;
A = 16'h007B; B = 16'h0037; #100;
A = 16'h007B; B = 16'h0038; #100;
A = 16'h007B; B = 16'h0039; #100;
A = 16'h007B; B = 16'h003A; #100;
A = 16'h007B; B = 16'h003B; #100;
A = 16'h007B; B = 16'h003C; #100;
A = 16'h007B; B = 16'h003D; #100;
A = 16'h007B; B = 16'h003E; #100;
A = 16'h007B; B = 16'h003F; #100;
A = 16'h007B; B = 16'h0040; #100;
A = 16'h007B; B = 16'h0041; #100;
A = 16'h007B; B = 16'h0042; #100;
A = 16'h007B; B = 16'h0043; #100;
A = 16'h007B; B = 16'h0044; #100;
A = 16'h007B; B = 16'h0045; #100;
A = 16'h007B; B = 16'h0046; #100;
A = 16'h007B; B = 16'h0047; #100;
A = 16'h007B; B = 16'h0048; #100;
A = 16'h007B; B = 16'h0049; #100;
A = 16'h007B; B = 16'h004A; #100;
A = 16'h007B; B = 16'h004B; #100;
A = 16'h007B; B = 16'h004C; #100;
A = 16'h007B; B = 16'h004D; #100;
A = 16'h007B; B = 16'h004E; #100;
A = 16'h007B; B = 16'h004F; #100;
A = 16'h007B; B = 16'h0050; #100;
A = 16'h007B; B = 16'h0051; #100;
A = 16'h007B; B = 16'h0052; #100;
A = 16'h007B; B = 16'h0053; #100;
A = 16'h007B; B = 16'h0054; #100;
A = 16'h007B; B = 16'h0055; #100;
A = 16'h007B; B = 16'h0056; #100;
A = 16'h007B; B = 16'h0057; #100;
A = 16'h007B; B = 16'h0058; #100;
A = 16'h007B; B = 16'h0059; #100;
A = 16'h007B; B = 16'h005A; #100;
A = 16'h007B; B = 16'h005B; #100;
A = 16'h007B; B = 16'h005C; #100;
A = 16'h007B; B = 16'h005D; #100;
A = 16'h007B; B = 16'h005E; #100;
A = 16'h007B; B = 16'h005F; #100;
A = 16'h007B; B = 16'h0060; #100;
A = 16'h007B; B = 16'h0061; #100;
A = 16'h007B; B = 16'h0062; #100;
A = 16'h007B; B = 16'h0063; #100;
A = 16'h007B; B = 16'h0064; #100;
A = 16'h007B; B = 16'h0065; #100;
A = 16'h007B; B = 16'h0066; #100;
A = 16'h007B; B = 16'h0067; #100;
A = 16'h007B; B = 16'h0068; #100;
A = 16'h007B; B = 16'h0069; #100;
A = 16'h007B; B = 16'h006A; #100;
A = 16'h007B; B = 16'h006B; #100;
A = 16'h007B; B = 16'h006C; #100;
A = 16'h007B; B = 16'h006D; #100;
A = 16'h007B; B = 16'h006E; #100;
A = 16'h007B; B = 16'h006F; #100;
A = 16'h007B; B = 16'h0070; #100;
A = 16'h007B; B = 16'h0071; #100;
A = 16'h007B; B = 16'h0072; #100;
A = 16'h007B; B = 16'h0073; #100;
A = 16'h007B; B = 16'h0074; #100;
A = 16'h007B; B = 16'h0075; #100;
A = 16'h007B; B = 16'h0076; #100;
A = 16'h007B; B = 16'h0077; #100;
A = 16'h007B; B = 16'h0078; #100;
A = 16'h007B; B = 16'h0079; #100;
A = 16'h007B; B = 16'h007A; #100;
A = 16'h007B; B = 16'h007B; #100;
A = 16'h007B; B = 16'h007C; #100;
A = 16'h007B; B = 16'h007D; #100;
A = 16'h007B; B = 16'h007E; #100;
A = 16'h007B; B = 16'h007F; #100;
A = 16'h007B; B = 16'h0080; #100;
A = 16'h007B; B = 16'h0081; #100;
A = 16'h007B; B = 16'h0082; #100;
A = 16'h007B; B = 16'h0083; #100;
A = 16'h007B; B = 16'h0084; #100;
A = 16'h007B; B = 16'h0085; #100;
A = 16'h007B; B = 16'h0086; #100;
A = 16'h007B; B = 16'h0087; #100;
A = 16'h007B; B = 16'h0088; #100;
A = 16'h007B; B = 16'h0089; #100;
A = 16'h007B; B = 16'h008A; #100;
A = 16'h007B; B = 16'h008B; #100;
A = 16'h007B; B = 16'h008C; #100;
A = 16'h007B; B = 16'h008D; #100;
A = 16'h007B; B = 16'h008E; #100;
A = 16'h007B; B = 16'h008F; #100;
A = 16'h007B; B = 16'h0090; #100;
A = 16'h007B; B = 16'h0091; #100;
A = 16'h007B; B = 16'h0092; #100;
A = 16'h007B; B = 16'h0093; #100;
A = 16'h007B; B = 16'h0094; #100;
A = 16'h007B; B = 16'h0095; #100;
A = 16'h007B; B = 16'h0096; #100;
A = 16'h007B; B = 16'h0097; #100;
A = 16'h007B; B = 16'h0098; #100;
A = 16'h007B; B = 16'h0099; #100;
A = 16'h007B; B = 16'h009A; #100;
A = 16'h007B; B = 16'h009B; #100;
A = 16'h007B; B = 16'h009C; #100;
A = 16'h007B; B = 16'h009D; #100;
A = 16'h007B; B = 16'h009E; #100;
A = 16'h007B; B = 16'h009F; #100;
A = 16'h007B; B = 16'h00A0; #100;
A = 16'h007B; B = 16'h00A1; #100;
A = 16'h007B; B = 16'h00A2; #100;
A = 16'h007B; B = 16'h00A3; #100;
A = 16'h007B; B = 16'h00A4; #100;
A = 16'h007B; B = 16'h00A5; #100;
A = 16'h007B; B = 16'h00A6; #100;
A = 16'h007B; B = 16'h00A7; #100;
A = 16'h007B; B = 16'h00A8; #100;
A = 16'h007B; B = 16'h00A9; #100;
A = 16'h007B; B = 16'h00AA; #100;
A = 16'h007B; B = 16'h00AB; #100;
A = 16'h007B; B = 16'h00AC; #100;
A = 16'h007B; B = 16'h00AD; #100;
A = 16'h007B; B = 16'h00AE; #100;
A = 16'h007B; B = 16'h00AF; #100;
A = 16'h007B; B = 16'h00B0; #100;
A = 16'h007B; B = 16'h00B1; #100;
A = 16'h007B; B = 16'h00B2; #100;
A = 16'h007B; B = 16'h00B3; #100;
A = 16'h007B; B = 16'h00B4; #100;
A = 16'h007B; B = 16'h00B5; #100;
A = 16'h007B; B = 16'h00B6; #100;
A = 16'h007B; B = 16'h00B7; #100;
A = 16'h007B; B = 16'h00B8; #100;
A = 16'h007B; B = 16'h00B9; #100;
A = 16'h007B; B = 16'h00BA; #100;
A = 16'h007B; B = 16'h00BB; #100;
A = 16'h007B; B = 16'h00BC; #100;
A = 16'h007B; B = 16'h00BD; #100;
A = 16'h007B; B = 16'h00BE; #100;
A = 16'h007B; B = 16'h00BF; #100;
A = 16'h007B; B = 16'h00C0; #100;
A = 16'h007B; B = 16'h00C1; #100;
A = 16'h007B; B = 16'h00C2; #100;
A = 16'h007B; B = 16'h00C3; #100;
A = 16'h007B; B = 16'h00C4; #100;
A = 16'h007B; B = 16'h00C5; #100;
A = 16'h007B; B = 16'h00C6; #100;
A = 16'h007B; B = 16'h00C7; #100;
A = 16'h007B; B = 16'h00C8; #100;
A = 16'h007B; B = 16'h00C9; #100;
A = 16'h007B; B = 16'h00CA; #100;
A = 16'h007B; B = 16'h00CB; #100;
A = 16'h007B; B = 16'h00CC; #100;
A = 16'h007B; B = 16'h00CD; #100;
A = 16'h007B; B = 16'h00CE; #100;
A = 16'h007B; B = 16'h00CF; #100;
A = 16'h007B; B = 16'h00D0; #100;
A = 16'h007B; B = 16'h00D1; #100;
A = 16'h007B; B = 16'h00D2; #100;
A = 16'h007B; B = 16'h00D3; #100;
A = 16'h007B; B = 16'h00D4; #100;
A = 16'h007B; B = 16'h00D5; #100;
A = 16'h007B; B = 16'h00D6; #100;
A = 16'h007B; B = 16'h00D7; #100;
A = 16'h007B; B = 16'h00D8; #100;
A = 16'h007B; B = 16'h00D9; #100;
A = 16'h007B; B = 16'h00DA; #100;
A = 16'h007B; B = 16'h00DB; #100;
A = 16'h007B; B = 16'h00DC; #100;
A = 16'h007B; B = 16'h00DD; #100;
A = 16'h007B; B = 16'h00DE; #100;
A = 16'h007B; B = 16'h00DF; #100;
A = 16'h007B; B = 16'h00E0; #100;
A = 16'h007B; B = 16'h00E1; #100;
A = 16'h007B; B = 16'h00E2; #100;
A = 16'h007B; B = 16'h00E3; #100;
A = 16'h007B; B = 16'h00E4; #100;
A = 16'h007B; B = 16'h00E5; #100;
A = 16'h007B; B = 16'h00E6; #100;
A = 16'h007B; B = 16'h00E7; #100;
A = 16'h007B; B = 16'h00E8; #100;
A = 16'h007B; B = 16'h00E9; #100;
A = 16'h007B; B = 16'h00EA; #100;
A = 16'h007B; B = 16'h00EB; #100;
A = 16'h007B; B = 16'h00EC; #100;
A = 16'h007B; B = 16'h00ED; #100;
A = 16'h007B; B = 16'h00EE; #100;
A = 16'h007B; B = 16'h00EF; #100;
A = 16'h007B; B = 16'h00F0; #100;
A = 16'h007B; B = 16'h00F1; #100;
A = 16'h007B; B = 16'h00F2; #100;
A = 16'h007B; B = 16'h00F3; #100;
A = 16'h007B; B = 16'h00F4; #100;
A = 16'h007B; B = 16'h00F5; #100;
A = 16'h007B; B = 16'h00F6; #100;
A = 16'h007B; B = 16'h00F7; #100;
A = 16'h007B; B = 16'h00F8; #100;
A = 16'h007B; B = 16'h00F9; #100;
A = 16'h007B; B = 16'h00FA; #100;
A = 16'h007B; B = 16'h00FB; #100;
A = 16'h007B; B = 16'h00FC; #100;
A = 16'h007B; B = 16'h00FD; #100;
A = 16'h007B; B = 16'h00FE; #100;
A = 16'h007B; B = 16'h00FF; #100;
A = 16'h007C; B = 16'h000; #100;
A = 16'h007C; B = 16'h001; #100;
A = 16'h007C; B = 16'h002; #100;
A = 16'h007C; B = 16'h003; #100;
A = 16'h007C; B = 16'h004; #100;
A = 16'h007C; B = 16'h005; #100;
A = 16'h007C; B = 16'h006; #100;
A = 16'h007C; B = 16'h007; #100;
A = 16'h007C; B = 16'h008; #100;
A = 16'h007C; B = 16'h009; #100;
A = 16'h007C; B = 16'h00A; #100;
A = 16'h007C; B = 16'h00B; #100;
A = 16'h007C; B = 16'h00C; #100;
A = 16'h007C; B = 16'h00D; #100;
A = 16'h007C; B = 16'h00E; #100;
A = 16'h007C; B = 16'h00F; #100;
A = 16'h007C; B = 16'h0010; #100;
A = 16'h007C; B = 16'h0011; #100;
A = 16'h007C; B = 16'h0012; #100;
A = 16'h007C; B = 16'h0013; #100;
A = 16'h007C; B = 16'h0014; #100;
A = 16'h007C; B = 16'h0015; #100;
A = 16'h007C; B = 16'h0016; #100;
A = 16'h007C; B = 16'h0017; #100;
A = 16'h007C; B = 16'h0018; #100;
A = 16'h007C; B = 16'h0019; #100;
A = 16'h007C; B = 16'h001A; #100;
A = 16'h007C; B = 16'h001B; #100;
A = 16'h007C; B = 16'h001C; #100;
A = 16'h007C; B = 16'h001D; #100;
A = 16'h007C; B = 16'h001E; #100;
A = 16'h007C; B = 16'h001F; #100;
A = 16'h007C; B = 16'h0020; #100;
A = 16'h007C; B = 16'h0021; #100;
A = 16'h007C; B = 16'h0022; #100;
A = 16'h007C; B = 16'h0023; #100;
A = 16'h007C; B = 16'h0024; #100;
A = 16'h007C; B = 16'h0025; #100;
A = 16'h007C; B = 16'h0026; #100;
A = 16'h007C; B = 16'h0027; #100;
A = 16'h007C; B = 16'h0028; #100;
A = 16'h007C; B = 16'h0029; #100;
A = 16'h007C; B = 16'h002A; #100;
A = 16'h007C; B = 16'h002B; #100;
A = 16'h007C; B = 16'h002C; #100;
A = 16'h007C; B = 16'h002D; #100;
A = 16'h007C; B = 16'h002E; #100;
A = 16'h007C; B = 16'h002F; #100;
A = 16'h007C; B = 16'h0030; #100;
A = 16'h007C; B = 16'h0031; #100;
A = 16'h007C; B = 16'h0032; #100;
A = 16'h007C; B = 16'h0033; #100;
A = 16'h007C; B = 16'h0034; #100;
A = 16'h007C; B = 16'h0035; #100;
A = 16'h007C; B = 16'h0036; #100;
A = 16'h007C; B = 16'h0037; #100;
A = 16'h007C; B = 16'h0038; #100;
A = 16'h007C; B = 16'h0039; #100;
A = 16'h007C; B = 16'h003A; #100;
A = 16'h007C; B = 16'h003B; #100;
A = 16'h007C; B = 16'h003C; #100;
A = 16'h007C; B = 16'h003D; #100;
A = 16'h007C; B = 16'h003E; #100;
A = 16'h007C; B = 16'h003F; #100;
A = 16'h007C; B = 16'h0040; #100;
A = 16'h007C; B = 16'h0041; #100;
A = 16'h007C; B = 16'h0042; #100;
A = 16'h007C; B = 16'h0043; #100;
A = 16'h007C; B = 16'h0044; #100;
A = 16'h007C; B = 16'h0045; #100;
A = 16'h007C; B = 16'h0046; #100;
A = 16'h007C; B = 16'h0047; #100;
A = 16'h007C; B = 16'h0048; #100;
A = 16'h007C; B = 16'h0049; #100;
A = 16'h007C; B = 16'h004A; #100;
A = 16'h007C; B = 16'h004B; #100;
A = 16'h007C; B = 16'h004C; #100;
A = 16'h007C; B = 16'h004D; #100;
A = 16'h007C; B = 16'h004E; #100;
A = 16'h007C; B = 16'h004F; #100;
A = 16'h007C; B = 16'h0050; #100;
A = 16'h007C; B = 16'h0051; #100;
A = 16'h007C; B = 16'h0052; #100;
A = 16'h007C; B = 16'h0053; #100;
A = 16'h007C; B = 16'h0054; #100;
A = 16'h007C; B = 16'h0055; #100;
A = 16'h007C; B = 16'h0056; #100;
A = 16'h007C; B = 16'h0057; #100;
A = 16'h007C; B = 16'h0058; #100;
A = 16'h007C; B = 16'h0059; #100;
A = 16'h007C; B = 16'h005A; #100;
A = 16'h007C; B = 16'h005B; #100;
A = 16'h007C; B = 16'h005C; #100;
A = 16'h007C; B = 16'h005D; #100;
A = 16'h007C; B = 16'h005E; #100;
A = 16'h007C; B = 16'h005F; #100;
A = 16'h007C; B = 16'h0060; #100;
A = 16'h007C; B = 16'h0061; #100;
A = 16'h007C; B = 16'h0062; #100;
A = 16'h007C; B = 16'h0063; #100;
A = 16'h007C; B = 16'h0064; #100;
A = 16'h007C; B = 16'h0065; #100;
A = 16'h007C; B = 16'h0066; #100;
A = 16'h007C; B = 16'h0067; #100;
A = 16'h007C; B = 16'h0068; #100;
A = 16'h007C; B = 16'h0069; #100;
A = 16'h007C; B = 16'h006A; #100;
A = 16'h007C; B = 16'h006B; #100;
A = 16'h007C; B = 16'h006C; #100;
A = 16'h007C; B = 16'h006D; #100;
A = 16'h007C; B = 16'h006E; #100;
A = 16'h007C; B = 16'h006F; #100;
A = 16'h007C; B = 16'h0070; #100;
A = 16'h007C; B = 16'h0071; #100;
A = 16'h007C; B = 16'h0072; #100;
A = 16'h007C; B = 16'h0073; #100;
A = 16'h007C; B = 16'h0074; #100;
A = 16'h007C; B = 16'h0075; #100;
A = 16'h007C; B = 16'h0076; #100;
A = 16'h007C; B = 16'h0077; #100;
A = 16'h007C; B = 16'h0078; #100;
A = 16'h007C; B = 16'h0079; #100;
A = 16'h007C; B = 16'h007A; #100;
A = 16'h007C; B = 16'h007B; #100;
A = 16'h007C; B = 16'h007C; #100;
A = 16'h007C; B = 16'h007D; #100;
A = 16'h007C; B = 16'h007E; #100;
A = 16'h007C; B = 16'h007F; #100;
A = 16'h007C; B = 16'h0080; #100;
A = 16'h007C; B = 16'h0081; #100;
A = 16'h007C; B = 16'h0082; #100;
A = 16'h007C; B = 16'h0083; #100;
A = 16'h007C; B = 16'h0084; #100;
A = 16'h007C; B = 16'h0085; #100;
A = 16'h007C; B = 16'h0086; #100;
A = 16'h007C; B = 16'h0087; #100;
A = 16'h007C; B = 16'h0088; #100;
A = 16'h007C; B = 16'h0089; #100;
A = 16'h007C; B = 16'h008A; #100;
A = 16'h007C; B = 16'h008B; #100;
A = 16'h007C; B = 16'h008C; #100;
A = 16'h007C; B = 16'h008D; #100;
A = 16'h007C; B = 16'h008E; #100;
A = 16'h007C; B = 16'h008F; #100;
A = 16'h007C; B = 16'h0090; #100;
A = 16'h007C; B = 16'h0091; #100;
A = 16'h007C; B = 16'h0092; #100;
A = 16'h007C; B = 16'h0093; #100;
A = 16'h007C; B = 16'h0094; #100;
A = 16'h007C; B = 16'h0095; #100;
A = 16'h007C; B = 16'h0096; #100;
A = 16'h007C; B = 16'h0097; #100;
A = 16'h007C; B = 16'h0098; #100;
A = 16'h007C; B = 16'h0099; #100;
A = 16'h007C; B = 16'h009A; #100;
A = 16'h007C; B = 16'h009B; #100;
A = 16'h007C; B = 16'h009C; #100;
A = 16'h007C; B = 16'h009D; #100;
A = 16'h007C; B = 16'h009E; #100;
A = 16'h007C; B = 16'h009F; #100;
A = 16'h007C; B = 16'h00A0; #100;
A = 16'h007C; B = 16'h00A1; #100;
A = 16'h007C; B = 16'h00A2; #100;
A = 16'h007C; B = 16'h00A3; #100;
A = 16'h007C; B = 16'h00A4; #100;
A = 16'h007C; B = 16'h00A5; #100;
A = 16'h007C; B = 16'h00A6; #100;
A = 16'h007C; B = 16'h00A7; #100;
A = 16'h007C; B = 16'h00A8; #100;
A = 16'h007C; B = 16'h00A9; #100;
A = 16'h007C; B = 16'h00AA; #100;
A = 16'h007C; B = 16'h00AB; #100;
A = 16'h007C; B = 16'h00AC; #100;
A = 16'h007C; B = 16'h00AD; #100;
A = 16'h007C; B = 16'h00AE; #100;
A = 16'h007C; B = 16'h00AF; #100;
A = 16'h007C; B = 16'h00B0; #100;
A = 16'h007C; B = 16'h00B1; #100;
A = 16'h007C; B = 16'h00B2; #100;
A = 16'h007C; B = 16'h00B3; #100;
A = 16'h007C; B = 16'h00B4; #100;
A = 16'h007C; B = 16'h00B5; #100;
A = 16'h007C; B = 16'h00B6; #100;
A = 16'h007C; B = 16'h00B7; #100;
A = 16'h007C; B = 16'h00B8; #100;
A = 16'h007C; B = 16'h00B9; #100;
A = 16'h007C; B = 16'h00BA; #100;
A = 16'h007C; B = 16'h00BB; #100;
A = 16'h007C; B = 16'h00BC; #100;
A = 16'h007C; B = 16'h00BD; #100;
A = 16'h007C; B = 16'h00BE; #100;
A = 16'h007C; B = 16'h00BF; #100;
A = 16'h007C; B = 16'h00C0; #100;
A = 16'h007C; B = 16'h00C1; #100;
A = 16'h007C; B = 16'h00C2; #100;
A = 16'h007C; B = 16'h00C3; #100;
A = 16'h007C; B = 16'h00C4; #100;
A = 16'h007C; B = 16'h00C5; #100;
A = 16'h007C; B = 16'h00C6; #100;
A = 16'h007C; B = 16'h00C7; #100;
A = 16'h007C; B = 16'h00C8; #100;
A = 16'h007C; B = 16'h00C9; #100;
A = 16'h007C; B = 16'h00CA; #100;
A = 16'h007C; B = 16'h00CB; #100;
A = 16'h007C; B = 16'h00CC; #100;
A = 16'h007C; B = 16'h00CD; #100;
A = 16'h007C; B = 16'h00CE; #100;
A = 16'h007C; B = 16'h00CF; #100;
A = 16'h007C; B = 16'h00D0; #100;
A = 16'h007C; B = 16'h00D1; #100;
A = 16'h007C; B = 16'h00D2; #100;
A = 16'h007C; B = 16'h00D3; #100;
A = 16'h007C; B = 16'h00D4; #100;
A = 16'h007C; B = 16'h00D5; #100;
A = 16'h007C; B = 16'h00D6; #100;
A = 16'h007C; B = 16'h00D7; #100;
A = 16'h007C; B = 16'h00D8; #100;
A = 16'h007C; B = 16'h00D9; #100;
A = 16'h007C; B = 16'h00DA; #100;
A = 16'h007C; B = 16'h00DB; #100;
A = 16'h007C; B = 16'h00DC; #100;
A = 16'h007C; B = 16'h00DD; #100;
A = 16'h007C; B = 16'h00DE; #100;
A = 16'h007C; B = 16'h00DF; #100;
A = 16'h007C; B = 16'h00E0; #100;
A = 16'h007C; B = 16'h00E1; #100;
A = 16'h007C; B = 16'h00E2; #100;
A = 16'h007C; B = 16'h00E3; #100;
A = 16'h007C; B = 16'h00E4; #100;
A = 16'h007C; B = 16'h00E5; #100;
A = 16'h007C; B = 16'h00E6; #100;
A = 16'h007C; B = 16'h00E7; #100;
A = 16'h007C; B = 16'h00E8; #100;
A = 16'h007C; B = 16'h00E9; #100;
A = 16'h007C; B = 16'h00EA; #100;
A = 16'h007C; B = 16'h00EB; #100;
A = 16'h007C; B = 16'h00EC; #100;
A = 16'h007C; B = 16'h00ED; #100;
A = 16'h007C; B = 16'h00EE; #100;
A = 16'h007C; B = 16'h00EF; #100;
A = 16'h007C; B = 16'h00F0; #100;
A = 16'h007C; B = 16'h00F1; #100;
A = 16'h007C; B = 16'h00F2; #100;
A = 16'h007C; B = 16'h00F3; #100;
A = 16'h007C; B = 16'h00F4; #100;
A = 16'h007C; B = 16'h00F5; #100;
A = 16'h007C; B = 16'h00F6; #100;
A = 16'h007C; B = 16'h00F7; #100;
A = 16'h007C; B = 16'h00F8; #100;
A = 16'h007C; B = 16'h00F9; #100;
A = 16'h007C; B = 16'h00FA; #100;
A = 16'h007C; B = 16'h00FB; #100;
A = 16'h007C; B = 16'h00FC; #100;
A = 16'h007C; B = 16'h00FD; #100;
A = 16'h007C; B = 16'h00FE; #100;
A = 16'h007C; B = 16'h00FF; #100;
A = 16'h007D; B = 16'h000; #100;
A = 16'h007D; B = 16'h001; #100;
A = 16'h007D; B = 16'h002; #100;
A = 16'h007D; B = 16'h003; #100;
A = 16'h007D; B = 16'h004; #100;
A = 16'h007D; B = 16'h005; #100;
A = 16'h007D; B = 16'h006; #100;
A = 16'h007D; B = 16'h007; #100;
A = 16'h007D; B = 16'h008; #100;
A = 16'h007D; B = 16'h009; #100;
A = 16'h007D; B = 16'h00A; #100;
A = 16'h007D; B = 16'h00B; #100;
A = 16'h007D; B = 16'h00C; #100;
A = 16'h007D; B = 16'h00D; #100;
A = 16'h007D; B = 16'h00E; #100;
A = 16'h007D; B = 16'h00F; #100;
A = 16'h007D; B = 16'h0010; #100;
A = 16'h007D; B = 16'h0011; #100;
A = 16'h007D; B = 16'h0012; #100;
A = 16'h007D; B = 16'h0013; #100;
A = 16'h007D; B = 16'h0014; #100;
A = 16'h007D; B = 16'h0015; #100;
A = 16'h007D; B = 16'h0016; #100;
A = 16'h007D; B = 16'h0017; #100;
A = 16'h007D; B = 16'h0018; #100;
A = 16'h007D; B = 16'h0019; #100;
A = 16'h007D; B = 16'h001A; #100;
A = 16'h007D; B = 16'h001B; #100;
A = 16'h007D; B = 16'h001C; #100;
A = 16'h007D; B = 16'h001D; #100;
A = 16'h007D; B = 16'h001E; #100;
A = 16'h007D; B = 16'h001F; #100;
A = 16'h007D; B = 16'h0020; #100;
A = 16'h007D; B = 16'h0021; #100;
A = 16'h007D; B = 16'h0022; #100;
A = 16'h007D; B = 16'h0023; #100;
A = 16'h007D; B = 16'h0024; #100;
A = 16'h007D; B = 16'h0025; #100;
A = 16'h007D; B = 16'h0026; #100;
A = 16'h007D; B = 16'h0027; #100;
A = 16'h007D; B = 16'h0028; #100;
A = 16'h007D; B = 16'h0029; #100;
A = 16'h007D; B = 16'h002A; #100;
A = 16'h007D; B = 16'h002B; #100;
A = 16'h007D; B = 16'h002C; #100;
A = 16'h007D; B = 16'h002D; #100;
A = 16'h007D; B = 16'h002E; #100;
A = 16'h007D; B = 16'h002F; #100;
A = 16'h007D; B = 16'h0030; #100;
A = 16'h007D; B = 16'h0031; #100;
A = 16'h007D; B = 16'h0032; #100;
A = 16'h007D; B = 16'h0033; #100;
A = 16'h007D; B = 16'h0034; #100;
A = 16'h007D; B = 16'h0035; #100;
A = 16'h007D; B = 16'h0036; #100;
A = 16'h007D; B = 16'h0037; #100;
A = 16'h007D; B = 16'h0038; #100;
A = 16'h007D; B = 16'h0039; #100;
A = 16'h007D; B = 16'h003A; #100;
A = 16'h007D; B = 16'h003B; #100;
A = 16'h007D; B = 16'h003C; #100;
A = 16'h007D; B = 16'h003D; #100;
A = 16'h007D; B = 16'h003E; #100;
A = 16'h007D; B = 16'h003F; #100;
A = 16'h007D; B = 16'h0040; #100;
A = 16'h007D; B = 16'h0041; #100;
A = 16'h007D; B = 16'h0042; #100;
A = 16'h007D; B = 16'h0043; #100;
A = 16'h007D; B = 16'h0044; #100;
A = 16'h007D; B = 16'h0045; #100;
A = 16'h007D; B = 16'h0046; #100;
A = 16'h007D; B = 16'h0047; #100;
A = 16'h007D; B = 16'h0048; #100;
A = 16'h007D; B = 16'h0049; #100;
A = 16'h007D; B = 16'h004A; #100;
A = 16'h007D; B = 16'h004B; #100;
A = 16'h007D; B = 16'h004C; #100;
A = 16'h007D; B = 16'h004D; #100;
A = 16'h007D; B = 16'h004E; #100;
A = 16'h007D; B = 16'h004F; #100;
A = 16'h007D; B = 16'h0050; #100;
A = 16'h007D; B = 16'h0051; #100;
A = 16'h007D; B = 16'h0052; #100;
A = 16'h007D; B = 16'h0053; #100;
A = 16'h007D; B = 16'h0054; #100;
A = 16'h007D; B = 16'h0055; #100;
A = 16'h007D; B = 16'h0056; #100;
A = 16'h007D; B = 16'h0057; #100;
A = 16'h007D; B = 16'h0058; #100;
A = 16'h007D; B = 16'h0059; #100;
A = 16'h007D; B = 16'h005A; #100;
A = 16'h007D; B = 16'h005B; #100;
A = 16'h007D; B = 16'h005C; #100;
A = 16'h007D; B = 16'h005D; #100;
A = 16'h007D; B = 16'h005E; #100;
A = 16'h007D; B = 16'h005F; #100;
A = 16'h007D; B = 16'h0060; #100;
A = 16'h007D; B = 16'h0061; #100;
A = 16'h007D; B = 16'h0062; #100;
A = 16'h007D; B = 16'h0063; #100;
A = 16'h007D; B = 16'h0064; #100;
A = 16'h007D; B = 16'h0065; #100;
A = 16'h007D; B = 16'h0066; #100;
A = 16'h007D; B = 16'h0067; #100;
A = 16'h007D; B = 16'h0068; #100;
A = 16'h007D; B = 16'h0069; #100;
A = 16'h007D; B = 16'h006A; #100;
A = 16'h007D; B = 16'h006B; #100;
A = 16'h007D; B = 16'h006C; #100;
A = 16'h007D; B = 16'h006D; #100;
A = 16'h007D; B = 16'h006E; #100;
A = 16'h007D; B = 16'h006F; #100;
A = 16'h007D; B = 16'h0070; #100;
A = 16'h007D; B = 16'h0071; #100;
A = 16'h007D; B = 16'h0072; #100;
A = 16'h007D; B = 16'h0073; #100;
A = 16'h007D; B = 16'h0074; #100;
A = 16'h007D; B = 16'h0075; #100;
A = 16'h007D; B = 16'h0076; #100;
A = 16'h007D; B = 16'h0077; #100;
A = 16'h007D; B = 16'h0078; #100;
A = 16'h007D; B = 16'h0079; #100;
A = 16'h007D; B = 16'h007A; #100;
A = 16'h007D; B = 16'h007B; #100;
A = 16'h007D; B = 16'h007C; #100;
A = 16'h007D; B = 16'h007D; #100;
A = 16'h007D; B = 16'h007E; #100;
A = 16'h007D; B = 16'h007F; #100;
A = 16'h007D; B = 16'h0080; #100;
A = 16'h007D; B = 16'h0081; #100;
A = 16'h007D; B = 16'h0082; #100;
A = 16'h007D; B = 16'h0083; #100;
A = 16'h007D; B = 16'h0084; #100;
A = 16'h007D; B = 16'h0085; #100;
A = 16'h007D; B = 16'h0086; #100;
A = 16'h007D; B = 16'h0087; #100;
A = 16'h007D; B = 16'h0088; #100;
A = 16'h007D; B = 16'h0089; #100;
A = 16'h007D; B = 16'h008A; #100;
A = 16'h007D; B = 16'h008B; #100;
A = 16'h007D; B = 16'h008C; #100;
A = 16'h007D; B = 16'h008D; #100;
A = 16'h007D; B = 16'h008E; #100;
A = 16'h007D; B = 16'h008F; #100;
A = 16'h007D; B = 16'h0090; #100;
A = 16'h007D; B = 16'h0091; #100;
A = 16'h007D; B = 16'h0092; #100;
A = 16'h007D; B = 16'h0093; #100;
A = 16'h007D; B = 16'h0094; #100;
A = 16'h007D; B = 16'h0095; #100;
A = 16'h007D; B = 16'h0096; #100;
A = 16'h007D; B = 16'h0097; #100;
A = 16'h007D; B = 16'h0098; #100;
A = 16'h007D; B = 16'h0099; #100;
A = 16'h007D; B = 16'h009A; #100;
A = 16'h007D; B = 16'h009B; #100;
A = 16'h007D; B = 16'h009C; #100;
A = 16'h007D; B = 16'h009D; #100;
A = 16'h007D; B = 16'h009E; #100;
A = 16'h007D; B = 16'h009F; #100;
A = 16'h007D; B = 16'h00A0; #100;
A = 16'h007D; B = 16'h00A1; #100;
A = 16'h007D; B = 16'h00A2; #100;
A = 16'h007D; B = 16'h00A3; #100;
A = 16'h007D; B = 16'h00A4; #100;
A = 16'h007D; B = 16'h00A5; #100;
A = 16'h007D; B = 16'h00A6; #100;
A = 16'h007D; B = 16'h00A7; #100;
A = 16'h007D; B = 16'h00A8; #100;
A = 16'h007D; B = 16'h00A9; #100;
A = 16'h007D; B = 16'h00AA; #100;
A = 16'h007D; B = 16'h00AB; #100;
A = 16'h007D; B = 16'h00AC; #100;
A = 16'h007D; B = 16'h00AD; #100;
A = 16'h007D; B = 16'h00AE; #100;
A = 16'h007D; B = 16'h00AF; #100;
A = 16'h007D; B = 16'h00B0; #100;
A = 16'h007D; B = 16'h00B1; #100;
A = 16'h007D; B = 16'h00B2; #100;
A = 16'h007D; B = 16'h00B3; #100;
A = 16'h007D; B = 16'h00B4; #100;
A = 16'h007D; B = 16'h00B5; #100;
A = 16'h007D; B = 16'h00B6; #100;
A = 16'h007D; B = 16'h00B7; #100;
A = 16'h007D; B = 16'h00B8; #100;
A = 16'h007D; B = 16'h00B9; #100;
A = 16'h007D; B = 16'h00BA; #100;
A = 16'h007D; B = 16'h00BB; #100;
A = 16'h007D; B = 16'h00BC; #100;
A = 16'h007D; B = 16'h00BD; #100;
A = 16'h007D; B = 16'h00BE; #100;
A = 16'h007D; B = 16'h00BF; #100;
A = 16'h007D; B = 16'h00C0; #100;
A = 16'h007D; B = 16'h00C1; #100;
A = 16'h007D; B = 16'h00C2; #100;
A = 16'h007D; B = 16'h00C3; #100;
A = 16'h007D; B = 16'h00C4; #100;
A = 16'h007D; B = 16'h00C5; #100;
A = 16'h007D; B = 16'h00C6; #100;
A = 16'h007D; B = 16'h00C7; #100;
A = 16'h007D; B = 16'h00C8; #100;
A = 16'h007D; B = 16'h00C9; #100;
A = 16'h007D; B = 16'h00CA; #100;
A = 16'h007D; B = 16'h00CB; #100;
A = 16'h007D; B = 16'h00CC; #100;
A = 16'h007D; B = 16'h00CD; #100;
A = 16'h007D; B = 16'h00CE; #100;
A = 16'h007D; B = 16'h00CF; #100;
A = 16'h007D; B = 16'h00D0; #100;
A = 16'h007D; B = 16'h00D1; #100;
A = 16'h007D; B = 16'h00D2; #100;
A = 16'h007D; B = 16'h00D3; #100;
A = 16'h007D; B = 16'h00D4; #100;
A = 16'h007D; B = 16'h00D5; #100;
A = 16'h007D; B = 16'h00D6; #100;
A = 16'h007D; B = 16'h00D7; #100;
A = 16'h007D; B = 16'h00D8; #100;
A = 16'h007D; B = 16'h00D9; #100;
A = 16'h007D; B = 16'h00DA; #100;
A = 16'h007D; B = 16'h00DB; #100;
A = 16'h007D; B = 16'h00DC; #100;
A = 16'h007D; B = 16'h00DD; #100;
A = 16'h007D; B = 16'h00DE; #100;
A = 16'h007D; B = 16'h00DF; #100;
A = 16'h007D; B = 16'h00E0; #100;
A = 16'h007D; B = 16'h00E1; #100;
A = 16'h007D; B = 16'h00E2; #100;
A = 16'h007D; B = 16'h00E3; #100;
A = 16'h007D; B = 16'h00E4; #100;
A = 16'h007D; B = 16'h00E5; #100;
A = 16'h007D; B = 16'h00E6; #100;
A = 16'h007D; B = 16'h00E7; #100;
A = 16'h007D; B = 16'h00E8; #100;
A = 16'h007D; B = 16'h00E9; #100;
A = 16'h007D; B = 16'h00EA; #100;
A = 16'h007D; B = 16'h00EB; #100;
A = 16'h007D; B = 16'h00EC; #100;
A = 16'h007D; B = 16'h00ED; #100;
A = 16'h007D; B = 16'h00EE; #100;
A = 16'h007D; B = 16'h00EF; #100;
A = 16'h007D; B = 16'h00F0; #100;
A = 16'h007D; B = 16'h00F1; #100;
A = 16'h007D; B = 16'h00F2; #100;
A = 16'h007D; B = 16'h00F3; #100;
A = 16'h007D; B = 16'h00F4; #100;
A = 16'h007D; B = 16'h00F5; #100;
A = 16'h007D; B = 16'h00F6; #100;
A = 16'h007D; B = 16'h00F7; #100;
A = 16'h007D; B = 16'h00F8; #100;
A = 16'h007D; B = 16'h00F9; #100;
A = 16'h007D; B = 16'h00FA; #100;
A = 16'h007D; B = 16'h00FB; #100;
A = 16'h007D; B = 16'h00FC; #100;
A = 16'h007D; B = 16'h00FD; #100;
A = 16'h007D; B = 16'h00FE; #100;
A = 16'h007D; B = 16'h00FF; #100;
A = 16'h007E; B = 16'h000; #100;
A = 16'h007E; B = 16'h001; #100;
A = 16'h007E; B = 16'h002; #100;
A = 16'h007E; B = 16'h003; #100;
A = 16'h007E; B = 16'h004; #100;
A = 16'h007E; B = 16'h005; #100;
A = 16'h007E; B = 16'h006; #100;
A = 16'h007E; B = 16'h007; #100;
A = 16'h007E; B = 16'h008; #100;
A = 16'h007E; B = 16'h009; #100;
A = 16'h007E; B = 16'h00A; #100;
A = 16'h007E; B = 16'h00B; #100;
A = 16'h007E; B = 16'h00C; #100;
A = 16'h007E; B = 16'h00D; #100;
A = 16'h007E; B = 16'h00E; #100;
A = 16'h007E; B = 16'h00F; #100;
A = 16'h007E; B = 16'h0010; #100;
A = 16'h007E; B = 16'h0011; #100;
A = 16'h007E; B = 16'h0012; #100;
A = 16'h007E; B = 16'h0013; #100;
A = 16'h007E; B = 16'h0014; #100;
A = 16'h007E; B = 16'h0015; #100;
A = 16'h007E; B = 16'h0016; #100;
A = 16'h007E; B = 16'h0017; #100;
A = 16'h007E; B = 16'h0018; #100;
A = 16'h007E; B = 16'h0019; #100;
A = 16'h007E; B = 16'h001A; #100;
A = 16'h007E; B = 16'h001B; #100;
A = 16'h007E; B = 16'h001C; #100;
A = 16'h007E; B = 16'h001D; #100;
A = 16'h007E; B = 16'h001E; #100;
A = 16'h007E; B = 16'h001F; #100;
A = 16'h007E; B = 16'h0020; #100;
A = 16'h007E; B = 16'h0021; #100;
A = 16'h007E; B = 16'h0022; #100;
A = 16'h007E; B = 16'h0023; #100;
A = 16'h007E; B = 16'h0024; #100;
A = 16'h007E; B = 16'h0025; #100;
A = 16'h007E; B = 16'h0026; #100;
A = 16'h007E; B = 16'h0027; #100;
A = 16'h007E; B = 16'h0028; #100;
A = 16'h007E; B = 16'h0029; #100;
A = 16'h007E; B = 16'h002A; #100;
A = 16'h007E; B = 16'h002B; #100;
A = 16'h007E; B = 16'h002C; #100;
A = 16'h007E; B = 16'h002D; #100;
A = 16'h007E; B = 16'h002E; #100;
A = 16'h007E; B = 16'h002F; #100;
A = 16'h007E; B = 16'h0030; #100;
A = 16'h007E; B = 16'h0031; #100;
A = 16'h007E; B = 16'h0032; #100;
A = 16'h007E; B = 16'h0033; #100;
A = 16'h007E; B = 16'h0034; #100;
A = 16'h007E; B = 16'h0035; #100;
A = 16'h007E; B = 16'h0036; #100;
A = 16'h007E; B = 16'h0037; #100;
A = 16'h007E; B = 16'h0038; #100;
A = 16'h007E; B = 16'h0039; #100;
A = 16'h007E; B = 16'h003A; #100;
A = 16'h007E; B = 16'h003B; #100;
A = 16'h007E; B = 16'h003C; #100;
A = 16'h007E; B = 16'h003D; #100;
A = 16'h007E; B = 16'h003E; #100;
A = 16'h007E; B = 16'h003F; #100;
A = 16'h007E; B = 16'h0040; #100;
A = 16'h007E; B = 16'h0041; #100;
A = 16'h007E; B = 16'h0042; #100;
A = 16'h007E; B = 16'h0043; #100;
A = 16'h007E; B = 16'h0044; #100;
A = 16'h007E; B = 16'h0045; #100;
A = 16'h007E; B = 16'h0046; #100;
A = 16'h007E; B = 16'h0047; #100;
A = 16'h007E; B = 16'h0048; #100;
A = 16'h007E; B = 16'h0049; #100;
A = 16'h007E; B = 16'h004A; #100;
A = 16'h007E; B = 16'h004B; #100;
A = 16'h007E; B = 16'h004C; #100;
A = 16'h007E; B = 16'h004D; #100;
A = 16'h007E; B = 16'h004E; #100;
A = 16'h007E; B = 16'h004F; #100;
A = 16'h007E; B = 16'h0050; #100;
A = 16'h007E; B = 16'h0051; #100;
A = 16'h007E; B = 16'h0052; #100;
A = 16'h007E; B = 16'h0053; #100;
A = 16'h007E; B = 16'h0054; #100;
A = 16'h007E; B = 16'h0055; #100;
A = 16'h007E; B = 16'h0056; #100;
A = 16'h007E; B = 16'h0057; #100;
A = 16'h007E; B = 16'h0058; #100;
A = 16'h007E; B = 16'h0059; #100;
A = 16'h007E; B = 16'h005A; #100;
A = 16'h007E; B = 16'h005B; #100;
A = 16'h007E; B = 16'h005C; #100;
A = 16'h007E; B = 16'h005D; #100;
A = 16'h007E; B = 16'h005E; #100;
A = 16'h007E; B = 16'h005F; #100;
A = 16'h007E; B = 16'h0060; #100;
A = 16'h007E; B = 16'h0061; #100;
A = 16'h007E; B = 16'h0062; #100;
A = 16'h007E; B = 16'h0063; #100;
A = 16'h007E; B = 16'h0064; #100;
A = 16'h007E; B = 16'h0065; #100;
A = 16'h007E; B = 16'h0066; #100;
A = 16'h007E; B = 16'h0067; #100;
A = 16'h007E; B = 16'h0068; #100;
A = 16'h007E; B = 16'h0069; #100;
A = 16'h007E; B = 16'h006A; #100;
A = 16'h007E; B = 16'h006B; #100;
A = 16'h007E; B = 16'h006C; #100;
A = 16'h007E; B = 16'h006D; #100;
A = 16'h007E; B = 16'h006E; #100;
A = 16'h007E; B = 16'h006F; #100;
A = 16'h007E; B = 16'h0070; #100;
A = 16'h007E; B = 16'h0071; #100;
A = 16'h007E; B = 16'h0072; #100;
A = 16'h007E; B = 16'h0073; #100;
A = 16'h007E; B = 16'h0074; #100;
A = 16'h007E; B = 16'h0075; #100;
A = 16'h007E; B = 16'h0076; #100;
A = 16'h007E; B = 16'h0077; #100;
A = 16'h007E; B = 16'h0078; #100;
A = 16'h007E; B = 16'h0079; #100;
A = 16'h007E; B = 16'h007A; #100;
A = 16'h007E; B = 16'h007B; #100;
A = 16'h007E; B = 16'h007C; #100;
A = 16'h007E; B = 16'h007D; #100;
A = 16'h007E; B = 16'h007E; #100;
A = 16'h007E; B = 16'h007F; #100;
A = 16'h007E; B = 16'h0080; #100;
A = 16'h007E; B = 16'h0081; #100;
A = 16'h007E; B = 16'h0082; #100;
A = 16'h007E; B = 16'h0083; #100;
A = 16'h007E; B = 16'h0084; #100;
A = 16'h007E; B = 16'h0085; #100;
A = 16'h007E; B = 16'h0086; #100;
A = 16'h007E; B = 16'h0087; #100;
A = 16'h007E; B = 16'h0088; #100;
A = 16'h007E; B = 16'h0089; #100;
A = 16'h007E; B = 16'h008A; #100;
A = 16'h007E; B = 16'h008B; #100;
A = 16'h007E; B = 16'h008C; #100;
A = 16'h007E; B = 16'h008D; #100;
A = 16'h007E; B = 16'h008E; #100;
A = 16'h007E; B = 16'h008F; #100;
A = 16'h007E; B = 16'h0090; #100;
A = 16'h007E; B = 16'h0091; #100;
A = 16'h007E; B = 16'h0092; #100;
A = 16'h007E; B = 16'h0093; #100;
A = 16'h007E; B = 16'h0094; #100;
A = 16'h007E; B = 16'h0095; #100;
A = 16'h007E; B = 16'h0096; #100;
A = 16'h007E; B = 16'h0097; #100;
A = 16'h007E; B = 16'h0098; #100;
A = 16'h007E; B = 16'h0099; #100;
A = 16'h007E; B = 16'h009A; #100;
A = 16'h007E; B = 16'h009B; #100;
A = 16'h007E; B = 16'h009C; #100;
A = 16'h007E; B = 16'h009D; #100;
A = 16'h007E; B = 16'h009E; #100;
A = 16'h007E; B = 16'h009F; #100;
A = 16'h007E; B = 16'h00A0; #100;
A = 16'h007E; B = 16'h00A1; #100;
A = 16'h007E; B = 16'h00A2; #100;
A = 16'h007E; B = 16'h00A3; #100;
A = 16'h007E; B = 16'h00A4; #100;
A = 16'h007E; B = 16'h00A5; #100;
A = 16'h007E; B = 16'h00A6; #100;
A = 16'h007E; B = 16'h00A7; #100;
A = 16'h007E; B = 16'h00A8; #100;
A = 16'h007E; B = 16'h00A9; #100;
A = 16'h007E; B = 16'h00AA; #100;
A = 16'h007E; B = 16'h00AB; #100;
A = 16'h007E; B = 16'h00AC; #100;
A = 16'h007E; B = 16'h00AD; #100;
A = 16'h007E; B = 16'h00AE; #100;
A = 16'h007E; B = 16'h00AF; #100;
A = 16'h007E; B = 16'h00B0; #100;
A = 16'h007E; B = 16'h00B1; #100;
A = 16'h007E; B = 16'h00B2; #100;
A = 16'h007E; B = 16'h00B3; #100;
A = 16'h007E; B = 16'h00B4; #100;
A = 16'h007E; B = 16'h00B5; #100;
A = 16'h007E; B = 16'h00B6; #100;
A = 16'h007E; B = 16'h00B7; #100;
A = 16'h007E; B = 16'h00B8; #100;
A = 16'h007E; B = 16'h00B9; #100;
A = 16'h007E; B = 16'h00BA; #100;
A = 16'h007E; B = 16'h00BB; #100;
A = 16'h007E; B = 16'h00BC; #100;
A = 16'h007E; B = 16'h00BD; #100;
A = 16'h007E; B = 16'h00BE; #100;
A = 16'h007E; B = 16'h00BF; #100;
A = 16'h007E; B = 16'h00C0; #100;
A = 16'h007E; B = 16'h00C1; #100;
A = 16'h007E; B = 16'h00C2; #100;
A = 16'h007E; B = 16'h00C3; #100;
A = 16'h007E; B = 16'h00C4; #100;
A = 16'h007E; B = 16'h00C5; #100;
A = 16'h007E; B = 16'h00C6; #100;
A = 16'h007E; B = 16'h00C7; #100;
A = 16'h007E; B = 16'h00C8; #100;
A = 16'h007E; B = 16'h00C9; #100;
A = 16'h007E; B = 16'h00CA; #100;
A = 16'h007E; B = 16'h00CB; #100;
A = 16'h007E; B = 16'h00CC; #100;
A = 16'h007E; B = 16'h00CD; #100;
A = 16'h007E; B = 16'h00CE; #100;
A = 16'h007E; B = 16'h00CF; #100;
A = 16'h007E; B = 16'h00D0; #100;
A = 16'h007E; B = 16'h00D1; #100;
A = 16'h007E; B = 16'h00D2; #100;
A = 16'h007E; B = 16'h00D3; #100;
A = 16'h007E; B = 16'h00D4; #100;
A = 16'h007E; B = 16'h00D5; #100;
A = 16'h007E; B = 16'h00D6; #100;
A = 16'h007E; B = 16'h00D7; #100;
A = 16'h007E; B = 16'h00D8; #100;
A = 16'h007E; B = 16'h00D9; #100;
A = 16'h007E; B = 16'h00DA; #100;
A = 16'h007E; B = 16'h00DB; #100;
A = 16'h007E; B = 16'h00DC; #100;
A = 16'h007E; B = 16'h00DD; #100;
A = 16'h007E; B = 16'h00DE; #100;
A = 16'h007E; B = 16'h00DF; #100;
A = 16'h007E; B = 16'h00E0; #100;
A = 16'h007E; B = 16'h00E1; #100;
A = 16'h007E; B = 16'h00E2; #100;
A = 16'h007E; B = 16'h00E3; #100;
A = 16'h007E; B = 16'h00E4; #100;
A = 16'h007E; B = 16'h00E5; #100;
A = 16'h007E; B = 16'h00E6; #100;
A = 16'h007E; B = 16'h00E7; #100;
A = 16'h007E; B = 16'h00E8; #100;
A = 16'h007E; B = 16'h00E9; #100;
A = 16'h007E; B = 16'h00EA; #100;
A = 16'h007E; B = 16'h00EB; #100;
A = 16'h007E; B = 16'h00EC; #100;
A = 16'h007E; B = 16'h00ED; #100;
A = 16'h007E; B = 16'h00EE; #100;
A = 16'h007E; B = 16'h00EF; #100;
A = 16'h007E; B = 16'h00F0; #100;
A = 16'h007E; B = 16'h00F1; #100;
A = 16'h007E; B = 16'h00F2; #100;
A = 16'h007E; B = 16'h00F3; #100;
A = 16'h007E; B = 16'h00F4; #100;
A = 16'h007E; B = 16'h00F5; #100;
A = 16'h007E; B = 16'h00F6; #100;
A = 16'h007E; B = 16'h00F7; #100;
A = 16'h007E; B = 16'h00F8; #100;
A = 16'h007E; B = 16'h00F9; #100;
A = 16'h007E; B = 16'h00FA; #100;
A = 16'h007E; B = 16'h00FB; #100;
A = 16'h007E; B = 16'h00FC; #100;
A = 16'h007E; B = 16'h00FD; #100;
A = 16'h007E; B = 16'h00FE; #100;
A = 16'h007E; B = 16'h00FF; #100;
A = 16'h007F; B = 16'h000; #100;
A = 16'h007F; B = 16'h001; #100;
A = 16'h007F; B = 16'h002; #100;
A = 16'h007F; B = 16'h003; #100;
A = 16'h007F; B = 16'h004; #100;
A = 16'h007F; B = 16'h005; #100;
A = 16'h007F; B = 16'h006; #100;
A = 16'h007F; B = 16'h007; #100;
A = 16'h007F; B = 16'h008; #100;
A = 16'h007F; B = 16'h009; #100;
A = 16'h007F; B = 16'h00A; #100;
A = 16'h007F; B = 16'h00B; #100;
A = 16'h007F; B = 16'h00C; #100;
A = 16'h007F; B = 16'h00D; #100;
A = 16'h007F; B = 16'h00E; #100;
A = 16'h007F; B = 16'h00F; #100;
A = 16'h007F; B = 16'h0010; #100;
A = 16'h007F; B = 16'h0011; #100;
A = 16'h007F; B = 16'h0012; #100;
A = 16'h007F; B = 16'h0013; #100;
A = 16'h007F; B = 16'h0014; #100;
A = 16'h007F; B = 16'h0015; #100;
A = 16'h007F; B = 16'h0016; #100;
A = 16'h007F; B = 16'h0017; #100;
A = 16'h007F; B = 16'h0018; #100;
A = 16'h007F; B = 16'h0019; #100;
A = 16'h007F; B = 16'h001A; #100;
A = 16'h007F; B = 16'h001B; #100;
A = 16'h007F; B = 16'h001C; #100;
A = 16'h007F; B = 16'h001D; #100;
A = 16'h007F; B = 16'h001E; #100;
A = 16'h007F; B = 16'h001F; #100;
A = 16'h007F; B = 16'h0020; #100;
A = 16'h007F; B = 16'h0021; #100;
A = 16'h007F; B = 16'h0022; #100;
A = 16'h007F; B = 16'h0023; #100;
A = 16'h007F; B = 16'h0024; #100;
A = 16'h007F; B = 16'h0025; #100;
A = 16'h007F; B = 16'h0026; #100;
A = 16'h007F; B = 16'h0027; #100;
A = 16'h007F; B = 16'h0028; #100;
A = 16'h007F; B = 16'h0029; #100;
A = 16'h007F; B = 16'h002A; #100;
A = 16'h007F; B = 16'h002B; #100;
A = 16'h007F; B = 16'h002C; #100;
A = 16'h007F; B = 16'h002D; #100;
A = 16'h007F; B = 16'h002E; #100;
A = 16'h007F; B = 16'h002F; #100;
A = 16'h007F; B = 16'h0030; #100;
A = 16'h007F; B = 16'h0031; #100;
A = 16'h007F; B = 16'h0032; #100;
A = 16'h007F; B = 16'h0033; #100;
A = 16'h007F; B = 16'h0034; #100;
A = 16'h007F; B = 16'h0035; #100;
A = 16'h007F; B = 16'h0036; #100;
A = 16'h007F; B = 16'h0037; #100;
A = 16'h007F; B = 16'h0038; #100;
A = 16'h007F; B = 16'h0039; #100;
A = 16'h007F; B = 16'h003A; #100;
A = 16'h007F; B = 16'h003B; #100;
A = 16'h007F; B = 16'h003C; #100;
A = 16'h007F; B = 16'h003D; #100;
A = 16'h007F; B = 16'h003E; #100;
A = 16'h007F; B = 16'h003F; #100;
A = 16'h007F; B = 16'h0040; #100;
A = 16'h007F; B = 16'h0041; #100;
A = 16'h007F; B = 16'h0042; #100;
A = 16'h007F; B = 16'h0043; #100;
A = 16'h007F; B = 16'h0044; #100;
A = 16'h007F; B = 16'h0045; #100;
A = 16'h007F; B = 16'h0046; #100;
A = 16'h007F; B = 16'h0047; #100;
A = 16'h007F; B = 16'h0048; #100;
A = 16'h007F; B = 16'h0049; #100;
A = 16'h007F; B = 16'h004A; #100;
A = 16'h007F; B = 16'h004B; #100;
A = 16'h007F; B = 16'h004C; #100;
A = 16'h007F; B = 16'h004D; #100;
A = 16'h007F; B = 16'h004E; #100;
A = 16'h007F; B = 16'h004F; #100;
A = 16'h007F; B = 16'h0050; #100;
A = 16'h007F; B = 16'h0051; #100;
A = 16'h007F; B = 16'h0052; #100;
A = 16'h007F; B = 16'h0053; #100;
A = 16'h007F; B = 16'h0054; #100;
A = 16'h007F; B = 16'h0055; #100;
A = 16'h007F; B = 16'h0056; #100;
A = 16'h007F; B = 16'h0057; #100;
A = 16'h007F; B = 16'h0058; #100;
A = 16'h007F; B = 16'h0059; #100;
A = 16'h007F; B = 16'h005A; #100;
A = 16'h007F; B = 16'h005B; #100;
A = 16'h007F; B = 16'h005C; #100;
A = 16'h007F; B = 16'h005D; #100;
A = 16'h007F; B = 16'h005E; #100;
A = 16'h007F; B = 16'h005F; #100;
A = 16'h007F; B = 16'h0060; #100;
A = 16'h007F; B = 16'h0061; #100;
A = 16'h007F; B = 16'h0062; #100;
A = 16'h007F; B = 16'h0063; #100;
A = 16'h007F; B = 16'h0064; #100;
A = 16'h007F; B = 16'h0065; #100;
A = 16'h007F; B = 16'h0066; #100;
A = 16'h007F; B = 16'h0067; #100;
A = 16'h007F; B = 16'h0068; #100;
A = 16'h007F; B = 16'h0069; #100;
A = 16'h007F; B = 16'h006A; #100;
A = 16'h007F; B = 16'h006B; #100;
A = 16'h007F; B = 16'h006C; #100;
A = 16'h007F; B = 16'h006D; #100;
A = 16'h007F; B = 16'h006E; #100;
A = 16'h007F; B = 16'h006F; #100;
A = 16'h007F; B = 16'h0070; #100;
A = 16'h007F; B = 16'h0071; #100;
A = 16'h007F; B = 16'h0072; #100;
A = 16'h007F; B = 16'h0073; #100;
A = 16'h007F; B = 16'h0074; #100;
A = 16'h007F; B = 16'h0075; #100;
A = 16'h007F; B = 16'h0076; #100;
A = 16'h007F; B = 16'h0077; #100;
A = 16'h007F; B = 16'h0078; #100;
A = 16'h007F; B = 16'h0079; #100;
A = 16'h007F; B = 16'h007A; #100;
A = 16'h007F; B = 16'h007B; #100;
A = 16'h007F; B = 16'h007C; #100;
A = 16'h007F; B = 16'h007D; #100;
A = 16'h007F; B = 16'h007E; #100;
A = 16'h007F; B = 16'h007F; #100;
A = 16'h007F; B = 16'h0080; #100;
A = 16'h007F; B = 16'h0081; #100;
A = 16'h007F; B = 16'h0082; #100;
A = 16'h007F; B = 16'h0083; #100;
A = 16'h007F; B = 16'h0084; #100;
A = 16'h007F; B = 16'h0085; #100;
A = 16'h007F; B = 16'h0086; #100;
A = 16'h007F; B = 16'h0087; #100;
A = 16'h007F; B = 16'h0088; #100;
A = 16'h007F; B = 16'h0089; #100;
A = 16'h007F; B = 16'h008A; #100;
A = 16'h007F; B = 16'h008B; #100;
A = 16'h007F; B = 16'h008C; #100;
A = 16'h007F; B = 16'h008D; #100;
A = 16'h007F; B = 16'h008E; #100;
A = 16'h007F; B = 16'h008F; #100;
A = 16'h007F; B = 16'h0090; #100;
A = 16'h007F; B = 16'h0091; #100;
A = 16'h007F; B = 16'h0092; #100;
A = 16'h007F; B = 16'h0093; #100;
A = 16'h007F; B = 16'h0094; #100;
A = 16'h007F; B = 16'h0095; #100;
A = 16'h007F; B = 16'h0096; #100;
A = 16'h007F; B = 16'h0097; #100;
A = 16'h007F; B = 16'h0098; #100;
A = 16'h007F; B = 16'h0099; #100;
A = 16'h007F; B = 16'h009A; #100;
A = 16'h007F; B = 16'h009B; #100;
A = 16'h007F; B = 16'h009C; #100;
A = 16'h007F; B = 16'h009D; #100;
A = 16'h007F; B = 16'h009E; #100;
A = 16'h007F; B = 16'h009F; #100;
A = 16'h007F; B = 16'h00A0; #100;
A = 16'h007F; B = 16'h00A1; #100;
A = 16'h007F; B = 16'h00A2; #100;
A = 16'h007F; B = 16'h00A3; #100;
A = 16'h007F; B = 16'h00A4; #100;
A = 16'h007F; B = 16'h00A5; #100;
A = 16'h007F; B = 16'h00A6; #100;
A = 16'h007F; B = 16'h00A7; #100;
A = 16'h007F; B = 16'h00A8; #100;
A = 16'h007F; B = 16'h00A9; #100;
A = 16'h007F; B = 16'h00AA; #100;
A = 16'h007F; B = 16'h00AB; #100;
A = 16'h007F; B = 16'h00AC; #100;
A = 16'h007F; B = 16'h00AD; #100;
A = 16'h007F; B = 16'h00AE; #100;
A = 16'h007F; B = 16'h00AF; #100;
A = 16'h007F; B = 16'h00B0; #100;
A = 16'h007F; B = 16'h00B1; #100;
A = 16'h007F; B = 16'h00B2; #100;
A = 16'h007F; B = 16'h00B3; #100;
A = 16'h007F; B = 16'h00B4; #100;
A = 16'h007F; B = 16'h00B5; #100;
A = 16'h007F; B = 16'h00B6; #100;
A = 16'h007F; B = 16'h00B7; #100;
A = 16'h007F; B = 16'h00B8; #100;
A = 16'h007F; B = 16'h00B9; #100;
A = 16'h007F; B = 16'h00BA; #100;
A = 16'h007F; B = 16'h00BB; #100;
A = 16'h007F; B = 16'h00BC; #100;
A = 16'h007F; B = 16'h00BD; #100;
A = 16'h007F; B = 16'h00BE; #100;
A = 16'h007F; B = 16'h00BF; #100;
A = 16'h007F; B = 16'h00C0; #100;
A = 16'h007F; B = 16'h00C1; #100;
A = 16'h007F; B = 16'h00C2; #100;
A = 16'h007F; B = 16'h00C3; #100;
A = 16'h007F; B = 16'h00C4; #100;
A = 16'h007F; B = 16'h00C5; #100;
A = 16'h007F; B = 16'h00C6; #100;
A = 16'h007F; B = 16'h00C7; #100;
A = 16'h007F; B = 16'h00C8; #100;
A = 16'h007F; B = 16'h00C9; #100;
A = 16'h007F; B = 16'h00CA; #100;
A = 16'h007F; B = 16'h00CB; #100;
A = 16'h007F; B = 16'h00CC; #100;
A = 16'h007F; B = 16'h00CD; #100;
A = 16'h007F; B = 16'h00CE; #100;
A = 16'h007F; B = 16'h00CF; #100;
A = 16'h007F; B = 16'h00D0; #100;
A = 16'h007F; B = 16'h00D1; #100;
A = 16'h007F; B = 16'h00D2; #100;
A = 16'h007F; B = 16'h00D3; #100;
A = 16'h007F; B = 16'h00D4; #100;
A = 16'h007F; B = 16'h00D5; #100;
A = 16'h007F; B = 16'h00D6; #100;
A = 16'h007F; B = 16'h00D7; #100;
A = 16'h007F; B = 16'h00D8; #100;
A = 16'h007F; B = 16'h00D9; #100;
A = 16'h007F; B = 16'h00DA; #100;
A = 16'h007F; B = 16'h00DB; #100;
A = 16'h007F; B = 16'h00DC; #100;
A = 16'h007F; B = 16'h00DD; #100;
A = 16'h007F; B = 16'h00DE; #100;
A = 16'h007F; B = 16'h00DF; #100;
A = 16'h007F; B = 16'h00E0; #100;
A = 16'h007F; B = 16'h00E1; #100;
A = 16'h007F; B = 16'h00E2; #100;
A = 16'h007F; B = 16'h00E3; #100;
A = 16'h007F; B = 16'h00E4; #100;
A = 16'h007F; B = 16'h00E5; #100;
A = 16'h007F; B = 16'h00E6; #100;
A = 16'h007F; B = 16'h00E7; #100;
A = 16'h007F; B = 16'h00E8; #100;
A = 16'h007F; B = 16'h00E9; #100;
A = 16'h007F; B = 16'h00EA; #100;
A = 16'h007F; B = 16'h00EB; #100;
A = 16'h007F; B = 16'h00EC; #100;
A = 16'h007F; B = 16'h00ED; #100;
A = 16'h007F; B = 16'h00EE; #100;
A = 16'h007F; B = 16'h00EF; #100;
A = 16'h007F; B = 16'h00F0; #100;
A = 16'h007F; B = 16'h00F1; #100;
A = 16'h007F; B = 16'h00F2; #100;
A = 16'h007F; B = 16'h00F3; #100;
A = 16'h007F; B = 16'h00F4; #100;
A = 16'h007F; B = 16'h00F5; #100;
A = 16'h007F; B = 16'h00F6; #100;
A = 16'h007F; B = 16'h00F7; #100;
A = 16'h007F; B = 16'h00F8; #100;
A = 16'h007F; B = 16'h00F9; #100;
A = 16'h007F; B = 16'h00FA; #100;
A = 16'h007F; B = 16'h00FB; #100;
A = 16'h007F; B = 16'h00FC; #100;
A = 16'h007F; B = 16'h00FD; #100;
A = 16'h007F; B = 16'h00FE; #100;
A = 16'h007F; B = 16'h00FF; #100;
A = 16'h0080; B = 16'h000; #100;
A = 16'h0080; B = 16'h001; #100;
A = 16'h0080; B = 16'h002; #100;
A = 16'h0080; B = 16'h003; #100;
A = 16'h0080; B = 16'h004; #100;
A = 16'h0080; B = 16'h005; #100;
A = 16'h0080; B = 16'h006; #100;
A = 16'h0080; B = 16'h007; #100;
A = 16'h0080; B = 16'h008; #100;
A = 16'h0080; B = 16'h009; #100;
A = 16'h0080; B = 16'h00A; #100;
A = 16'h0080; B = 16'h00B; #100;
A = 16'h0080; B = 16'h00C; #100;
A = 16'h0080; B = 16'h00D; #100;
A = 16'h0080; B = 16'h00E; #100;
A = 16'h0080; B = 16'h00F; #100;
A = 16'h0080; B = 16'h0010; #100;
A = 16'h0080; B = 16'h0011; #100;
A = 16'h0080; B = 16'h0012; #100;
A = 16'h0080; B = 16'h0013; #100;
A = 16'h0080; B = 16'h0014; #100;
A = 16'h0080; B = 16'h0015; #100;
A = 16'h0080; B = 16'h0016; #100;
A = 16'h0080; B = 16'h0017; #100;
A = 16'h0080; B = 16'h0018; #100;
A = 16'h0080; B = 16'h0019; #100;
A = 16'h0080; B = 16'h001A; #100;
A = 16'h0080; B = 16'h001B; #100;
A = 16'h0080; B = 16'h001C; #100;
A = 16'h0080; B = 16'h001D; #100;
A = 16'h0080; B = 16'h001E; #100;
A = 16'h0080; B = 16'h001F; #100;
A = 16'h0080; B = 16'h0020; #100;
A = 16'h0080; B = 16'h0021; #100;
A = 16'h0080; B = 16'h0022; #100;
A = 16'h0080; B = 16'h0023; #100;
A = 16'h0080; B = 16'h0024; #100;
A = 16'h0080; B = 16'h0025; #100;
A = 16'h0080; B = 16'h0026; #100;
A = 16'h0080; B = 16'h0027; #100;
A = 16'h0080; B = 16'h0028; #100;
A = 16'h0080; B = 16'h0029; #100;
A = 16'h0080; B = 16'h002A; #100;
A = 16'h0080; B = 16'h002B; #100;
A = 16'h0080; B = 16'h002C; #100;
A = 16'h0080; B = 16'h002D; #100;
A = 16'h0080; B = 16'h002E; #100;
A = 16'h0080; B = 16'h002F; #100;
A = 16'h0080; B = 16'h0030; #100;
A = 16'h0080; B = 16'h0031; #100;
A = 16'h0080; B = 16'h0032; #100;
A = 16'h0080; B = 16'h0033; #100;
A = 16'h0080; B = 16'h0034; #100;
A = 16'h0080; B = 16'h0035; #100;
A = 16'h0080; B = 16'h0036; #100;
A = 16'h0080; B = 16'h0037; #100;
A = 16'h0080; B = 16'h0038; #100;
A = 16'h0080; B = 16'h0039; #100;
A = 16'h0080; B = 16'h003A; #100;
A = 16'h0080; B = 16'h003B; #100;
A = 16'h0080; B = 16'h003C; #100;
A = 16'h0080; B = 16'h003D; #100;
A = 16'h0080; B = 16'h003E; #100;
A = 16'h0080; B = 16'h003F; #100;
A = 16'h0080; B = 16'h0040; #100;
A = 16'h0080; B = 16'h0041; #100;
A = 16'h0080; B = 16'h0042; #100;
A = 16'h0080; B = 16'h0043; #100;
A = 16'h0080; B = 16'h0044; #100;
A = 16'h0080; B = 16'h0045; #100;
A = 16'h0080; B = 16'h0046; #100;
A = 16'h0080; B = 16'h0047; #100;
A = 16'h0080; B = 16'h0048; #100;
A = 16'h0080; B = 16'h0049; #100;
A = 16'h0080; B = 16'h004A; #100;
A = 16'h0080; B = 16'h004B; #100;
A = 16'h0080; B = 16'h004C; #100;
A = 16'h0080; B = 16'h004D; #100;
A = 16'h0080; B = 16'h004E; #100;
A = 16'h0080; B = 16'h004F; #100;
A = 16'h0080; B = 16'h0050; #100;
A = 16'h0080; B = 16'h0051; #100;
A = 16'h0080; B = 16'h0052; #100;
A = 16'h0080; B = 16'h0053; #100;
A = 16'h0080; B = 16'h0054; #100;
A = 16'h0080; B = 16'h0055; #100;
A = 16'h0080; B = 16'h0056; #100;
A = 16'h0080; B = 16'h0057; #100;
A = 16'h0080; B = 16'h0058; #100;
A = 16'h0080; B = 16'h0059; #100;
A = 16'h0080; B = 16'h005A; #100;
A = 16'h0080; B = 16'h005B; #100;
A = 16'h0080; B = 16'h005C; #100;
A = 16'h0080; B = 16'h005D; #100;
A = 16'h0080; B = 16'h005E; #100;
A = 16'h0080; B = 16'h005F; #100;
A = 16'h0080; B = 16'h0060; #100;
A = 16'h0080; B = 16'h0061; #100;
A = 16'h0080; B = 16'h0062; #100;
A = 16'h0080; B = 16'h0063; #100;
A = 16'h0080; B = 16'h0064; #100;
A = 16'h0080; B = 16'h0065; #100;
A = 16'h0080; B = 16'h0066; #100;
A = 16'h0080; B = 16'h0067; #100;
A = 16'h0080; B = 16'h0068; #100;
A = 16'h0080; B = 16'h0069; #100;
A = 16'h0080; B = 16'h006A; #100;
A = 16'h0080; B = 16'h006B; #100;
A = 16'h0080; B = 16'h006C; #100;
A = 16'h0080; B = 16'h006D; #100;
A = 16'h0080; B = 16'h006E; #100;
A = 16'h0080; B = 16'h006F; #100;
A = 16'h0080; B = 16'h0070; #100;
A = 16'h0080; B = 16'h0071; #100;
A = 16'h0080; B = 16'h0072; #100;
A = 16'h0080; B = 16'h0073; #100;
A = 16'h0080; B = 16'h0074; #100;
A = 16'h0080; B = 16'h0075; #100;
A = 16'h0080; B = 16'h0076; #100;
A = 16'h0080; B = 16'h0077; #100;
A = 16'h0080; B = 16'h0078; #100;
A = 16'h0080; B = 16'h0079; #100;
A = 16'h0080; B = 16'h007A; #100;
A = 16'h0080; B = 16'h007B; #100;
A = 16'h0080; B = 16'h007C; #100;
A = 16'h0080; B = 16'h007D; #100;
A = 16'h0080; B = 16'h007E; #100;
A = 16'h0080; B = 16'h007F; #100;
A = 16'h0080; B = 16'h0080; #100;
A = 16'h0080; B = 16'h0081; #100;
A = 16'h0080; B = 16'h0082; #100;
A = 16'h0080; B = 16'h0083; #100;
A = 16'h0080; B = 16'h0084; #100;
A = 16'h0080; B = 16'h0085; #100;
A = 16'h0080; B = 16'h0086; #100;
A = 16'h0080; B = 16'h0087; #100;
A = 16'h0080; B = 16'h0088; #100;
A = 16'h0080; B = 16'h0089; #100;
A = 16'h0080; B = 16'h008A; #100;
A = 16'h0080; B = 16'h008B; #100;
A = 16'h0080; B = 16'h008C; #100;
A = 16'h0080; B = 16'h008D; #100;
A = 16'h0080; B = 16'h008E; #100;
A = 16'h0080; B = 16'h008F; #100;
A = 16'h0080; B = 16'h0090; #100;
A = 16'h0080; B = 16'h0091; #100;
A = 16'h0080; B = 16'h0092; #100;
A = 16'h0080; B = 16'h0093; #100;
A = 16'h0080; B = 16'h0094; #100;
A = 16'h0080; B = 16'h0095; #100;
A = 16'h0080; B = 16'h0096; #100;
A = 16'h0080; B = 16'h0097; #100;
A = 16'h0080; B = 16'h0098; #100;
A = 16'h0080; B = 16'h0099; #100;
A = 16'h0080; B = 16'h009A; #100;
A = 16'h0080; B = 16'h009B; #100;
A = 16'h0080; B = 16'h009C; #100;
A = 16'h0080; B = 16'h009D; #100;
A = 16'h0080; B = 16'h009E; #100;
A = 16'h0080; B = 16'h009F; #100;
A = 16'h0080; B = 16'h00A0; #100;
A = 16'h0080; B = 16'h00A1; #100;
A = 16'h0080; B = 16'h00A2; #100;
A = 16'h0080; B = 16'h00A3; #100;
A = 16'h0080; B = 16'h00A4; #100;
A = 16'h0080; B = 16'h00A5; #100;
A = 16'h0080; B = 16'h00A6; #100;
A = 16'h0080; B = 16'h00A7; #100;
A = 16'h0080; B = 16'h00A8; #100;
A = 16'h0080; B = 16'h00A9; #100;
A = 16'h0080; B = 16'h00AA; #100;
A = 16'h0080; B = 16'h00AB; #100;
A = 16'h0080; B = 16'h00AC; #100;
A = 16'h0080; B = 16'h00AD; #100;
A = 16'h0080; B = 16'h00AE; #100;
A = 16'h0080; B = 16'h00AF; #100;
A = 16'h0080; B = 16'h00B0; #100;
A = 16'h0080; B = 16'h00B1; #100;
A = 16'h0080; B = 16'h00B2; #100;
A = 16'h0080; B = 16'h00B3; #100;
A = 16'h0080; B = 16'h00B4; #100;
A = 16'h0080; B = 16'h00B5; #100;
A = 16'h0080; B = 16'h00B6; #100;
A = 16'h0080; B = 16'h00B7; #100;
A = 16'h0080; B = 16'h00B8; #100;
A = 16'h0080; B = 16'h00B9; #100;
A = 16'h0080; B = 16'h00BA; #100;
A = 16'h0080; B = 16'h00BB; #100;
A = 16'h0080; B = 16'h00BC; #100;
A = 16'h0080; B = 16'h00BD; #100;
A = 16'h0080; B = 16'h00BE; #100;
A = 16'h0080; B = 16'h00BF; #100;
A = 16'h0080; B = 16'h00C0; #100;
A = 16'h0080; B = 16'h00C1; #100;
A = 16'h0080; B = 16'h00C2; #100;
A = 16'h0080; B = 16'h00C3; #100;
A = 16'h0080; B = 16'h00C4; #100;
A = 16'h0080; B = 16'h00C5; #100;
A = 16'h0080; B = 16'h00C6; #100;
A = 16'h0080; B = 16'h00C7; #100;
A = 16'h0080; B = 16'h00C8; #100;
A = 16'h0080; B = 16'h00C9; #100;
A = 16'h0080; B = 16'h00CA; #100;
A = 16'h0080; B = 16'h00CB; #100;
A = 16'h0080; B = 16'h00CC; #100;
A = 16'h0080; B = 16'h00CD; #100;
A = 16'h0080; B = 16'h00CE; #100;
A = 16'h0080; B = 16'h00CF; #100;
A = 16'h0080; B = 16'h00D0; #100;
A = 16'h0080; B = 16'h00D1; #100;
A = 16'h0080; B = 16'h00D2; #100;
A = 16'h0080; B = 16'h00D3; #100;
A = 16'h0080; B = 16'h00D4; #100;
A = 16'h0080; B = 16'h00D5; #100;
A = 16'h0080; B = 16'h00D6; #100;
A = 16'h0080; B = 16'h00D7; #100;
A = 16'h0080; B = 16'h00D8; #100;
A = 16'h0080; B = 16'h00D9; #100;
A = 16'h0080; B = 16'h00DA; #100;
A = 16'h0080; B = 16'h00DB; #100;
A = 16'h0080; B = 16'h00DC; #100;
A = 16'h0080; B = 16'h00DD; #100;
A = 16'h0080; B = 16'h00DE; #100;
A = 16'h0080; B = 16'h00DF; #100;
A = 16'h0080; B = 16'h00E0; #100;
A = 16'h0080; B = 16'h00E1; #100;
A = 16'h0080; B = 16'h00E2; #100;
A = 16'h0080; B = 16'h00E3; #100;
A = 16'h0080; B = 16'h00E4; #100;
A = 16'h0080; B = 16'h00E5; #100;
A = 16'h0080; B = 16'h00E6; #100;
A = 16'h0080; B = 16'h00E7; #100;
A = 16'h0080; B = 16'h00E8; #100;
A = 16'h0080; B = 16'h00E9; #100;
A = 16'h0080; B = 16'h00EA; #100;
A = 16'h0080; B = 16'h00EB; #100;
A = 16'h0080; B = 16'h00EC; #100;
A = 16'h0080; B = 16'h00ED; #100;
A = 16'h0080; B = 16'h00EE; #100;
A = 16'h0080; B = 16'h00EF; #100;
A = 16'h0080; B = 16'h00F0; #100;
A = 16'h0080; B = 16'h00F1; #100;
A = 16'h0080; B = 16'h00F2; #100;
A = 16'h0080; B = 16'h00F3; #100;
A = 16'h0080; B = 16'h00F4; #100;
A = 16'h0080; B = 16'h00F5; #100;
A = 16'h0080; B = 16'h00F6; #100;
A = 16'h0080; B = 16'h00F7; #100;
A = 16'h0080; B = 16'h00F8; #100;
A = 16'h0080; B = 16'h00F9; #100;
A = 16'h0080; B = 16'h00FA; #100;
A = 16'h0080; B = 16'h00FB; #100;
A = 16'h0080; B = 16'h00FC; #100;
A = 16'h0080; B = 16'h00FD; #100;
A = 16'h0080; B = 16'h00FE; #100;
A = 16'h0080; B = 16'h00FF; #100;
A = 16'h0081; B = 16'h000; #100;
A = 16'h0081; B = 16'h001; #100;
A = 16'h0081; B = 16'h002; #100;
A = 16'h0081; B = 16'h003; #100;
A = 16'h0081; B = 16'h004; #100;
A = 16'h0081; B = 16'h005; #100;
A = 16'h0081; B = 16'h006; #100;
A = 16'h0081; B = 16'h007; #100;
A = 16'h0081; B = 16'h008; #100;
A = 16'h0081; B = 16'h009; #100;
A = 16'h0081; B = 16'h00A; #100;
A = 16'h0081; B = 16'h00B; #100;
A = 16'h0081; B = 16'h00C; #100;
A = 16'h0081; B = 16'h00D; #100;
A = 16'h0081; B = 16'h00E; #100;
A = 16'h0081; B = 16'h00F; #100;
A = 16'h0081; B = 16'h0010; #100;
A = 16'h0081; B = 16'h0011; #100;
A = 16'h0081; B = 16'h0012; #100;
A = 16'h0081; B = 16'h0013; #100;
A = 16'h0081; B = 16'h0014; #100;
A = 16'h0081; B = 16'h0015; #100;
A = 16'h0081; B = 16'h0016; #100;
A = 16'h0081; B = 16'h0017; #100;
A = 16'h0081; B = 16'h0018; #100;
A = 16'h0081; B = 16'h0019; #100;
A = 16'h0081; B = 16'h001A; #100;
A = 16'h0081; B = 16'h001B; #100;
A = 16'h0081; B = 16'h001C; #100;
A = 16'h0081; B = 16'h001D; #100;
A = 16'h0081; B = 16'h001E; #100;
A = 16'h0081; B = 16'h001F; #100;
A = 16'h0081; B = 16'h0020; #100;
A = 16'h0081; B = 16'h0021; #100;
A = 16'h0081; B = 16'h0022; #100;
A = 16'h0081; B = 16'h0023; #100;
A = 16'h0081; B = 16'h0024; #100;
A = 16'h0081; B = 16'h0025; #100;
A = 16'h0081; B = 16'h0026; #100;
A = 16'h0081; B = 16'h0027; #100;
A = 16'h0081; B = 16'h0028; #100;
A = 16'h0081; B = 16'h0029; #100;
A = 16'h0081; B = 16'h002A; #100;
A = 16'h0081; B = 16'h002B; #100;
A = 16'h0081; B = 16'h002C; #100;
A = 16'h0081; B = 16'h002D; #100;
A = 16'h0081; B = 16'h002E; #100;
A = 16'h0081; B = 16'h002F; #100;
A = 16'h0081; B = 16'h0030; #100;
A = 16'h0081; B = 16'h0031; #100;
A = 16'h0081; B = 16'h0032; #100;
A = 16'h0081; B = 16'h0033; #100;
A = 16'h0081; B = 16'h0034; #100;
A = 16'h0081; B = 16'h0035; #100;
A = 16'h0081; B = 16'h0036; #100;
A = 16'h0081; B = 16'h0037; #100;
A = 16'h0081; B = 16'h0038; #100;
A = 16'h0081; B = 16'h0039; #100;
A = 16'h0081; B = 16'h003A; #100;
A = 16'h0081; B = 16'h003B; #100;
A = 16'h0081; B = 16'h003C; #100;
A = 16'h0081; B = 16'h003D; #100;
A = 16'h0081; B = 16'h003E; #100;
A = 16'h0081; B = 16'h003F; #100;
A = 16'h0081; B = 16'h0040; #100;
A = 16'h0081; B = 16'h0041; #100;
A = 16'h0081; B = 16'h0042; #100;
A = 16'h0081; B = 16'h0043; #100;
A = 16'h0081; B = 16'h0044; #100;
A = 16'h0081; B = 16'h0045; #100;
A = 16'h0081; B = 16'h0046; #100;
A = 16'h0081; B = 16'h0047; #100;
A = 16'h0081; B = 16'h0048; #100;
A = 16'h0081; B = 16'h0049; #100;
A = 16'h0081; B = 16'h004A; #100;
A = 16'h0081; B = 16'h004B; #100;
A = 16'h0081; B = 16'h004C; #100;
A = 16'h0081; B = 16'h004D; #100;
A = 16'h0081; B = 16'h004E; #100;
A = 16'h0081; B = 16'h004F; #100;
A = 16'h0081; B = 16'h0050; #100;
A = 16'h0081; B = 16'h0051; #100;
A = 16'h0081; B = 16'h0052; #100;
A = 16'h0081; B = 16'h0053; #100;
A = 16'h0081; B = 16'h0054; #100;
A = 16'h0081; B = 16'h0055; #100;
A = 16'h0081; B = 16'h0056; #100;
A = 16'h0081; B = 16'h0057; #100;
A = 16'h0081; B = 16'h0058; #100;
A = 16'h0081; B = 16'h0059; #100;
A = 16'h0081; B = 16'h005A; #100;
A = 16'h0081; B = 16'h005B; #100;
A = 16'h0081; B = 16'h005C; #100;
A = 16'h0081; B = 16'h005D; #100;
A = 16'h0081; B = 16'h005E; #100;
A = 16'h0081; B = 16'h005F; #100;
A = 16'h0081; B = 16'h0060; #100;
A = 16'h0081; B = 16'h0061; #100;
A = 16'h0081; B = 16'h0062; #100;
A = 16'h0081; B = 16'h0063; #100;
A = 16'h0081; B = 16'h0064; #100;
A = 16'h0081; B = 16'h0065; #100;
A = 16'h0081; B = 16'h0066; #100;
A = 16'h0081; B = 16'h0067; #100;
A = 16'h0081; B = 16'h0068; #100;
A = 16'h0081; B = 16'h0069; #100;
A = 16'h0081; B = 16'h006A; #100;
A = 16'h0081; B = 16'h006B; #100;
A = 16'h0081; B = 16'h006C; #100;
A = 16'h0081; B = 16'h006D; #100;
A = 16'h0081; B = 16'h006E; #100;
A = 16'h0081; B = 16'h006F; #100;
A = 16'h0081; B = 16'h0070; #100;
A = 16'h0081; B = 16'h0071; #100;
A = 16'h0081; B = 16'h0072; #100;
A = 16'h0081; B = 16'h0073; #100;
A = 16'h0081; B = 16'h0074; #100;
A = 16'h0081; B = 16'h0075; #100;
A = 16'h0081; B = 16'h0076; #100;
A = 16'h0081; B = 16'h0077; #100;
A = 16'h0081; B = 16'h0078; #100;
A = 16'h0081; B = 16'h0079; #100;
A = 16'h0081; B = 16'h007A; #100;
A = 16'h0081; B = 16'h007B; #100;
A = 16'h0081; B = 16'h007C; #100;
A = 16'h0081; B = 16'h007D; #100;
A = 16'h0081; B = 16'h007E; #100;
A = 16'h0081; B = 16'h007F; #100;
A = 16'h0081; B = 16'h0080; #100;
A = 16'h0081; B = 16'h0081; #100;
A = 16'h0081; B = 16'h0082; #100;
A = 16'h0081; B = 16'h0083; #100;
A = 16'h0081; B = 16'h0084; #100;
A = 16'h0081; B = 16'h0085; #100;
A = 16'h0081; B = 16'h0086; #100;
A = 16'h0081; B = 16'h0087; #100;
A = 16'h0081; B = 16'h0088; #100;
A = 16'h0081; B = 16'h0089; #100;
A = 16'h0081; B = 16'h008A; #100;
A = 16'h0081; B = 16'h008B; #100;
A = 16'h0081; B = 16'h008C; #100;
A = 16'h0081; B = 16'h008D; #100;
A = 16'h0081; B = 16'h008E; #100;
A = 16'h0081; B = 16'h008F; #100;
A = 16'h0081; B = 16'h0090; #100;
A = 16'h0081; B = 16'h0091; #100;
A = 16'h0081; B = 16'h0092; #100;
A = 16'h0081; B = 16'h0093; #100;
A = 16'h0081; B = 16'h0094; #100;
A = 16'h0081; B = 16'h0095; #100;
A = 16'h0081; B = 16'h0096; #100;
A = 16'h0081; B = 16'h0097; #100;
A = 16'h0081; B = 16'h0098; #100;
A = 16'h0081; B = 16'h0099; #100;
A = 16'h0081; B = 16'h009A; #100;
A = 16'h0081; B = 16'h009B; #100;
A = 16'h0081; B = 16'h009C; #100;
A = 16'h0081; B = 16'h009D; #100;
A = 16'h0081; B = 16'h009E; #100;
A = 16'h0081; B = 16'h009F; #100;
A = 16'h0081; B = 16'h00A0; #100;
A = 16'h0081; B = 16'h00A1; #100;
A = 16'h0081; B = 16'h00A2; #100;
A = 16'h0081; B = 16'h00A3; #100;
A = 16'h0081; B = 16'h00A4; #100;
A = 16'h0081; B = 16'h00A5; #100;
A = 16'h0081; B = 16'h00A6; #100;
A = 16'h0081; B = 16'h00A7; #100;
A = 16'h0081; B = 16'h00A8; #100;
A = 16'h0081; B = 16'h00A9; #100;
A = 16'h0081; B = 16'h00AA; #100;
A = 16'h0081; B = 16'h00AB; #100;
A = 16'h0081; B = 16'h00AC; #100;
A = 16'h0081; B = 16'h00AD; #100;
A = 16'h0081; B = 16'h00AE; #100;
A = 16'h0081; B = 16'h00AF; #100;
A = 16'h0081; B = 16'h00B0; #100;
A = 16'h0081; B = 16'h00B1; #100;
A = 16'h0081; B = 16'h00B2; #100;
A = 16'h0081; B = 16'h00B3; #100;
A = 16'h0081; B = 16'h00B4; #100;
A = 16'h0081; B = 16'h00B5; #100;
A = 16'h0081; B = 16'h00B6; #100;
A = 16'h0081; B = 16'h00B7; #100;
A = 16'h0081; B = 16'h00B8; #100;
A = 16'h0081; B = 16'h00B9; #100;
A = 16'h0081; B = 16'h00BA; #100;
A = 16'h0081; B = 16'h00BB; #100;
A = 16'h0081; B = 16'h00BC; #100;
A = 16'h0081; B = 16'h00BD; #100;
A = 16'h0081; B = 16'h00BE; #100;
A = 16'h0081; B = 16'h00BF; #100;
A = 16'h0081; B = 16'h00C0; #100;
A = 16'h0081; B = 16'h00C1; #100;
A = 16'h0081; B = 16'h00C2; #100;
A = 16'h0081; B = 16'h00C3; #100;
A = 16'h0081; B = 16'h00C4; #100;
A = 16'h0081; B = 16'h00C5; #100;
A = 16'h0081; B = 16'h00C6; #100;
A = 16'h0081; B = 16'h00C7; #100;
A = 16'h0081; B = 16'h00C8; #100;
A = 16'h0081; B = 16'h00C9; #100;
A = 16'h0081; B = 16'h00CA; #100;
A = 16'h0081; B = 16'h00CB; #100;
A = 16'h0081; B = 16'h00CC; #100;
A = 16'h0081; B = 16'h00CD; #100;
A = 16'h0081; B = 16'h00CE; #100;
A = 16'h0081; B = 16'h00CF; #100;
A = 16'h0081; B = 16'h00D0; #100;
A = 16'h0081; B = 16'h00D1; #100;
A = 16'h0081; B = 16'h00D2; #100;
A = 16'h0081; B = 16'h00D3; #100;
A = 16'h0081; B = 16'h00D4; #100;
A = 16'h0081; B = 16'h00D5; #100;
A = 16'h0081; B = 16'h00D6; #100;
A = 16'h0081; B = 16'h00D7; #100;
A = 16'h0081; B = 16'h00D8; #100;
A = 16'h0081; B = 16'h00D9; #100;
A = 16'h0081; B = 16'h00DA; #100;
A = 16'h0081; B = 16'h00DB; #100;
A = 16'h0081; B = 16'h00DC; #100;
A = 16'h0081; B = 16'h00DD; #100;
A = 16'h0081; B = 16'h00DE; #100;
A = 16'h0081; B = 16'h00DF; #100;
A = 16'h0081; B = 16'h00E0; #100;
A = 16'h0081; B = 16'h00E1; #100;
A = 16'h0081; B = 16'h00E2; #100;
A = 16'h0081; B = 16'h00E3; #100;
A = 16'h0081; B = 16'h00E4; #100;
A = 16'h0081; B = 16'h00E5; #100;
A = 16'h0081; B = 16'h00E6; #100;
A = 16'h0081; B = 16'h00E7; #100;
A = 16'h0081; B = 16'h00E8; #100;
A = 16'h0081; B = 16'h00E9; #100;
A = 16'h0081; B = 16'h00EA; #100;
A = 16'h0081; B = 16'h00EB; #100;
A = 16'h0081; B = 16'h00EC; #100;
A = 16'h0081; B = 16'h00ED; #100;
A = 16'h0081; B = 16'h00EE; #100;
A = 16'h0081; B = 16'h00EF; #100;
A = 16'h0081; B = 16'h00F0; #100;
A = 16'h0081; B = 16'h00F1; #100;
A = 16'h0081; B = 16'h00F2; #100;
A = 16'h0081; B = 16'h00F3; #100;
A = 16'h0081; B = 16'h00F4; #100;
A = 16'h0081; B = 16'h00F5; #100;
A = 16'h0081; B = 16'h00F6; #100;
A = 16'h0081; B = 16'h00F7; #100;
A = 16'h0081; B = 16'h00F8; #100;
A = 16'h0081; B = 16'h00F9; #100;
A = 16'h0081; B = 16'h00FA; #100;
A = 16'h0081; B = 16'h00FB; #100;
A = 16'h0081; B = 16'h00FC; #100;
A = 16'h0081; B = 16'h00FD; #100;
A = 16'h0081; B = 16'h00FE; #100;
A = 16'h0081; B = 16'h00FF; #100;
A = 16'h0082; B = 16'h000; #100;
A = 16'h0082; B = 16'h001; #100;
A = 16'h0082; B = 16'h002; #100;
A = 16'h0082; B = 16'h003; #100;
A = 16'h0082; B = 16'h004; #100;
A = 16'h0082; B = 16'h005; #100;
A = 16'h0082; B = 16'h006; #100;
A = 16'h0082; B = 16'h007; #100;
A = 16'h0082; B = 16'h008; #100;
A = 16'h0082; B = 16'h009; #100;
A = 16'h0082; B = 16'h00A; #100;
A = 16'h0082; B = 16'h00B; #100;
A = 16'h0082; B = 16'h00C; #100;
A = 16'h0082; B = 16'h00D; #100;
A = 16'h0082; B = 16'h00E; #100;
A = 16'h0082; B = 16'h00F; #100;
A = 16'h0082; B = 16'h0010; #100;
A = 16'h0082; B = 16'h0011; #100;
A = 16'h0082; B = 16'h0012; #100;
A = 16'h0082; B = 16'h0013; #100;
A = 16'h0082; B = 16'h0014; #100;
A = 16'h0082; B = 16'h0015; #100;
A = 16'h0082; B = 16'h0016; #100;
A = 16'h0082; B = 16'h0017; #100;
A = 16'h0082; B = 16'h0018; #100;
A = 16'h0082; B = 16'h0019; #100;
A = 16'h0082; B = 16'h001A; #100;
A = 16'h0082; B = 16'h001B; #100;
A = 16'h0082; B = 16'h001C; #100;
A = 16'h0082; B = 16'h001D; #100;
A = 16'h0082; B = 16'h001E; #100;
A = 16'h0082; B = 16'h001F; #100;
A = 16'h0082; B = 16'h0020; #100;
A = 16'h0082; B = 16'h0021; #100;
A = 16'h0082; B = 16'h0022; #100;
A = 16'h0082; B = 16'h0023; #100;
A = 16'h0082; B = 16'h0024; #100;
A = 16'h0082; B = 16'h0025; #100;
A = 16'h0082; B = 16'h0026; #100;
A = 16'h0082; B = 16'h0027; #100;
A = 16'h0082; B = 16'h0028; #100;
A = 16'h0082; B = 16'h0029; #100;
A = 16'h0082; B = 16'h002A; #100;
A = 16'h0082; B = 16'h002B; #100;
A = 16'h0082; B = 16'h002C; #100;
A = 16'h0082; B = 16'h002D; #100;
A = 16'h0082; B = 16'h002E; #100;
A = 16'h0082; B = 16'h002F; #100;
A = 16'h0082; B = 16'h0030; #100;
A = 16'h0082; B = 16'h0031; #100;
A = 16'h0082; B = 16'h0032; #100;
A = 16'h0082; B = 16'h0033; #100;
A = 16'h0082; B = 16'h0034; #100;
A = 16'h0082; B = 16'h0035; #100;
A = 16'h0082; B = 16'h0036; #100;
A = 16'h0082; B = 16'h0037; #100;
A = 16'h0082; B = 16'h0038; #100;
A = 16'h0082; B = 16'h0039; #100;
A = 16'h0082; B = 16'h003A; #100;
A = 16'h0082; B = 16'h003B; #100;
A = 16'h0082; B = 16'h003C; #100;
A = 16'h0082; B = 16'h003D; #100;
A = 16'h0082; B = 16'h003E; #100;
A = 16'h0082; B = 16'h003F; #100;
A = 16'h0082; B = 16'h0040; #100;
A = 16'h0082; B = 16'h0041; #100;
A = 16'h0082; B = 16'h0042; #100;
A = 16'h0082; B = 16'h0043; #100;
A = 16'h0082; B = 16'h0044; #100;
A = 16'h0082; B = 16'h0045; #100;
A = 16'h0082; B = 16'h0046; #100;
A = 16'h0082; B = 16'h0047; #100;
A = 16'h0082; B = 16'h0048; #100;
A = 16'h0082; B = 16'h0049; #100;
A = 16'h0082; B = 16'h004A; #100;
A = 16'h0082; B = 16'h004B; #100;
A = 16'h0082; B = 16'h004C; #100;
A = 16'h0082; B = 16'h004D; #100;
A = 16'h0082; B = 16'h004E; #100;
A = 16'h0082; B = 16'h004F; #100;
A = 16'h0082; B = 16'h0050; #100;
A = 16'h0082; B = 16'h0051; #100;
A = 16'h0082; B = 16'h0052; #100;
A = 16'h0082; B = 16'h0053; #100;
A = 16'h0082; B = 16'h0054; #100;
A = 16'h0082; B = 16'h0055; #100;
A = 16'h0082; B = 16'h0056; #100;
A = 16'h0082; B = 16'h0057; #100;
A = 16'h0082; B = 16'h0058; #100;
A = 16'h0082; B = 16'h0059; #100;
A = 16'h0082; B = 16'h005A; #100;
A = 16'h0082; B = 16'h005B; #100;
A = 16'h0082; B = 16'h005C; #100;
A = 16'h0082; B = 16'h005D; #100;
A = 16'h0082; B = 16'h005E; #100;
A = 16'h0082; B = 16'h005F; #100;
A = 16'h0082; B = 16'h0060; #100;
A = 16'h0082; B = 16'h0061; #100;
A = 16'h0082; B = 16'h0062; #100;
A = 16'h0082; B = 16'h0063; #100;
A = 16'h0082; B = 16'h0064; #100;
A = 16'h0082; B = 16'h0065; #100;
A = 16'h0082; B = 16'h0066; #100;
A = 16'h0082; B = 16'h0067; #100;
A = 16'h0082; B = 16'h0068; #100;
A = 16'h0082; B = 16'h0069; #100;
A = 16'h0082; B = 16'h006A; #100;
A = 16'h0082; B = 16'h006B; #100;
A = 16'h0082; B = 16'h006C; #100;
A = 16'h0082; B = 16'h006D; #100;
A = 16'h0082; B = 16'h006E; #100;
A = 16'h0082; B = 16'h006F; #100;
A = 16'h0082; B = 16'h0070; #100;
A = 16'h0082; B = 16'h0071; #100;
A = 16'h0082; B = 16'h0072; #100;
A = 16'h0082; B = 16'h0073; #100;
A = 16'h0082; B = 16'h0074; #100;
A = 16'h0082; B = 16'h0075; #100;
A = 16'h0082; B = 16'h0076; #100;
A = 16'h0082; B = 16'h0077; #100;
A = 16'h0082; B = 16'h0078; #100;
A = 16'h0082; B = 16'h0079; #100;
A = 16'h0082; B = 16'h007A; #100;
A = 16'h0082; B = 16'h007B; #100;
A = 16'h0082; B = 16'h007C; #100;
A = 16'h0082; B = 16'h007D; #100;
A = 16'h0082; B = 16'h007E; #100;
A = 16'h0082; B = 16'h007F; #100;
A = 16'h0082; B = 16'h0080; #100;
A = 16'h0082; B = 16'h0081; #100;
A = 16'h0082; B = 16'h0082; #100;
A = 16'h0082; B = 16'h0083; #100;
A = 16'h0082; B = 16'h0084; #100;
A = 16'h0082; B = 16'h0085; #100;
A = 16'h0082; B = 16'h0086; #100;
A = 16'h0082; B = 16'h0087; #100;
A = 16'h0082; B = 16'h0088; #100;
A = 16'h0082; B = 16'h0089; #100;
A = 16'h0082; B = 16'h008A; #100;
A = 16'h0082; B = 16'h008B; #100;
A = 16'h0082; B = 16'h008C; #100;
A = 16'h0082; B = 16'h008D; #100;
A = 16'h0082; B = 16'h008E; #100;
A = 16'h0082; B = 16'h008F; #100;
A = 16'h0082; B = 16'h0090; #100;
A = 16'h0082; B = 16'h0091; #100;
A = 16'h0082; B = 16'h0092; #100;
A = 16'h0082; B = 16'h0093; #100;
A = 16'h0082; B = 16'h0094; #100;
A = 16'h0082; B = 16'h0095; #100;
A = 16'h0082; B = 16'h0096; #100;
A = 16'h0082; B = 16'h0097; #100;
A = 16'h0082; B = 16'h0098; #100;
A = 16'h0082; B = 16'h0099; #100;
A = 16'h0082; B = 16'h009A; #100;
A = 16'h0082; B = 16'h009B; #100;
A = 16'h0082; B = 16'h009C; #100;
A = 16'h0082; B = 16'h009D; #100;
A = 16'h0082; B = 16'h009E; #100;
A = 16'h0082; B = 16'h009F; #100;
A = 16'h0082; B = 16'h00A0; #100;
A = 16'h0082; B = 16'h00A1; #100;
A = 16'h0082; B = 16'h00A2; #100;
A = 16'h0082; B = 16'h00A3; #100;
A = 16'h0082; B = 16'h00A4; #100;
A = 16'h0082; B = 16'h00A5; #100;
A = 16'h0082; B = 16'h00A6; #100;
A = 16'h0082; B = 16'h00A7; #100;
A = 16'h0082; B = 16'h00A8; #100;
A = 16'h0082; B = 16'h00A9; #100;
A = 16'h0082; B = 16'h00AA; #100;
A = 16'h0082; B = 16'h00AB; #100;
A = 16'h0082; B = 16'h00AC; #100;
A = 16'h0082; B = 16'h00AD; #100;
A = 16'h0082; B = 16'h00AE; #100;
A = 16'h0082; B = 16'h00AF; #100;
A = 16'h0082; B = 16'h00B0; #100;
A = 16'h0082; B = 16'h00B1; #100;
A = 16'h0082; B = 16'h00B2; #100;
A = 16'h0082; B = 16'h00B3; #100;
A = 16'h0082; B = 16'h00B4; #100;
A = 16'h0082; B = 16'h00B5; #100;
A = 16'h0082; B = 16'h00B6; #100;
A = 16'h0082; B = 16'h00B7; #100;
A = 16'h0082; B = 16'h00B8; #100;
A = 16'h0082; B = 16'h00B9; #100;
A = 16'h0082; B = 16'h00BA; #100;
A = 16'h0082; B = 16'h00BB; #100;
A = 16'h0082; B = 16'h00BC; #100;
A = 16'h0082; B = 16'h00BD; #100;
A = 16'h0082; B = 16'h00BE; #100;
A = 16'h0082; B = 16'h00BF; #100;
A = 16'h0082; B = 16'h00C0; #100;
A = 16'h0082; B = 16'h00C1; #100;
A = 16'h0082; B = 16'h00C2; #100;
A = 16'h0082; B = 16'h00C3; #100;
A = 16'h0082; B = 16'h00C4; #100;
A = 16'h0082; B = 16'h00C5; #100;
A = 16'h0082; B = 16'h00C6; #100;
A = 16'h0082; B = 16'h00C7; #100;
A = 16'h0082; B = 16'h00C8; #100;
A = 16'h0082; B = 16'h00C9; #100;
A = 16'h0082; B = 16'h00CA; #100;
A = 16'h0082; B = 16'h00CB; #100;
A = 16'h0082; B = 16'h00CC; #100;
A = 16'h0082; B = 16'h00CD; #100;
A = 16'h0082; B = 16'h00CE; #100;
A = 16'h0082; B = 16'h00CF; #100;
A = 16'h0082; B = 16'h00D0; #100;
A = 16'h0082; B = 16'h00D1; #100;
A = 16'h0082; B = 16'h00D2; #100;
A = 16'h0082; B = 16'h00D3; #100;
A = 16'h0082; B = 16'h00D4; #100;
A = 16'h0082; B = 16'h00D5; #100;
A = 16'h0082; B = 16'h00D6; #100;
A = 16'h0082; B = 16'h00D7; #100;
A = 16'h0082; B = 16'h00D8; #100;
A = 16'h0082; B = 16'h00D9; #100;
A = 16'h0082; B = 16'h00DA; #100;
A = 16'h0082; B = 16'h00DB; #100;
A = 16'h0082; B = 16'h00DC; #100;
A = 16'h0082; B = 16'h00DD; #100;
A = 16'h0082; B = 16'h00DE; #100;
A = 16'h0082; B = 16'h00DF; #100;
A = 16'h0082; B = 16'h00E0; #100;
A = 16'h0082; B = 16'h00E1; #100;
A = 16'h0082; B = 16'h00E2; #100;
A = 16'h0082; B = 16'h00E3; #100;
A = 16'h0082; B = 16'h00E4; #100;
A = 16'h0082; B = 16'h00E5; #100;
A = 16'h0082; B = 16'h00E6; #100;
A = 16'h0082; B = 16'h00E7; #100;
A = 16'h0082; B = 16'h00E8; #100;
A = 16'h0082; B = 16'h00E9; #100;
A = 16'h0082; B = 16'h00EA; #100;
A = 16'h0082; B = 16'h00EB; #100;
A = 16'h0082; B = 16'h00EC; #100;
A = 16'h0082; B = 16'h00ED; #100;
A = 16'h0082; B = 16'h00EE; #100;
A = 16'h0082; B = 16'h00EF; #100;
A = 16'h0082; B = 16'h00F0; #100;
A = 16'h0082; B = 16'h00F1; #100;
A = 16'h0082; B = 16'h00F2; #100;
A = 16'h0082; B = 16'h00F3; #100;
A = 16'h0082; B = 16'h00F4; #100;
A = 16'h0082; B = 16'h00F5; #100;
A = 16'h0082; B = 16'h00F6; #100;
A = 16'h0082; B = 16'h00F7; #100;
A = 16'h0082; B = 16'h00F8; #100;
A = 16'h0082; B = 16'h00F9; #100;
A = 16'h0082; B = 16'h00FA; #100;
A = 16'h0082; B = 16'h00FB; #100;
A = 16'h0082; B = 16'h00FC; #100;
A = 16'h0082; B = 16'h00FD; #100;
A = 16'h0082; B = 16'h00FE; #100;
A = 16'h0082; B = 16'h00FF; #100;
A = 16'h0083; B = 16'h000; #100;
A = 16'h0083; B = 16'h001; #100;
A = 16'h0083; B = 16'h002; #100;
A = 16'h0083; B = 16'h003; #100;
A = 16'h0083; B = 16'h004; #100;
A = 16'h0083; B = 16'h005; #100;
A = 16'h0083; B = 16'h006; #100;
A = 16'h0083; B = 16'h007; #100;
A = 16'h0083; B = 16'h008; #100;
A = 16'h0083; B = 16'h009; #100;
A = 16'h0083; B = 16'h00A; #100;
A = 16'h0083; B = 16'h00B; #100;
A = 16'h0083; B = 16'h00C; #100;
A = 16'h0083; B = 16'h00D; #100;
A = 16'h0083; B = 16'h00E; #100;
A = 16'h0083; B = 16'h00F; #100;
A = 16'h0083; B = 16'h0010; #100;
A = 16'h0083; B = 16'h0011; #100;
A = 16'h0083; B = 16'h0012; #100;
A = 16'h0083; B = 16'h0013; #100;
A = 16'h0083; B = 16'h0014; #100;
A = 16'h0083; B = 16'h0015; #100;
A = 16'h0083; B = 16'h0016; #100;
A = 16'h0083; B = 16'h0017; #100;
A = 16'h0083; B = 16'h0018; #100;
A = 16'h0083; B = 16'h0019; #100;
A = 16'h0083; B = 16'h001A; #100;
A = 16'h0083; B = 16'h001B; #100;
A = 16'h0083; B = 16'h001C; #100;
A = 16'h0083; B = 16'h001D; #100;
A = 16'h0083; B = 16'h001E; #100;
A = 16'h0083; B = 16'h001F; #100;
A = 16'h0083; B = 16'h0020; #100;
A = 16'h0083; B = 16'h0021; #100;
A = 16'h0083; B = 16'h0022; #100;
A = 16'h0083; B = 16'h0023; #100;
A = 16'h0083; B = 16'h0024; #100;
A = 16'h0083; B = 16'h0025; #100;
A = 16'h0083; B = 16'h0026; #100;
A = 16'h0083; B = 16'h0027; #100;
A = 16'h0083; B = 16'h0028; #100;
A = 16'h0083; B = 16'h0029; #100;
A = 16'h0083; B = 16'h002A; #100;
A = 16'h0083; B = 16'h002B; #100;
A = 16'h0083; B = 16'h002C; #100;
A = 16'h0083; B = 16'h002D; #100;
A = 16'h0083; B = 16'h002E; #100;
A = 16'h0083; B = 16'h002F; #100;
A = 16'h0083; B = 16'h0030; #100;
A = 16'h0083; B = 16'h0031; #100;
A = 16'h0083; B = 16'h0032; #100;
A = 16'h0083; B = 16'h0033; #100;
A = 16'h0083; B = 16'h0034; #100;
A = 16'h0083; B = 16'h0035; #100;
A = 16'h0083; B = 16'h0036; #100;
A = 16'h0083; B = 16'h0037; #100;
A = 16'h0083; B = 16'h0038; #100;
A = 16'h0083; B = 16'h0039; #100;
A = 16'h0083; B = 16'h003A; #100;
A = 16'h0083; B = 16'h003B; #100;
A = 16'h0083; B = 16'h003C; #100;
A = 16'h0083; B = 16'h003D; #100;
A = 16'h0083; B = 16'h003E; #100;
A = 16'h0083; B = 16'h003F; #100;
A = 16'h0083; B = 16'h0040; #100;
A = 16'h0083; B = 16'h0041; #100;
A = 16'h0083; B = 16'h0042; #100;
A = 16'h0083; B = 16'h0043; #100;
A = 16'h0083; B = 16'h0044; #100;
A = 16'h0083; B = 16'h0045; #100;
A = 16'h0083; B = 16'h0046; #100;
A = 16'h0083; B = 16'h0047; #100;
A = 16'h0083; B = 16'h0048; #100;
A = 16'h0083; B = 16'h0049; #100;
A = 16'h0083; B = 16'h004A; #100;
A = 16'h0083; B = 16'h004B; #100;
A = 16'h0083; B = 16'h004C; #100;
A = 16'h0083; B = 16'h004D; #100;
A = 16'h0083; B = 16'h004E; #100;
A = 16'h0083; B = 16'h004F; #100;
A = 16'h0083; B = 16'h0050; #100;
A = 16'h0083; B = 16'h0051; #100;
A = 16'h0083; B = 16'h0052; #100;
A = 16'h0083; B = 16'h0053; #100;
A = 16'h0083; B = 16'h0054; #100;
A = 16'h0083; B = 16'h0055; #100;
A = 16'h0083; B = 16'h0056; #100;
A = 16'h0083; B = 16'h0057; #100;
A = 16'h0083; B = 16'h0058; #100;
A = 16'h0083; B = 16'h0059; #100;
A = 16'h0083; B = 16'h005A; #100;
A = 16'h0083; B = 16'h005B; #100;
A = 16'h0083; B = 16'h005C; #100;
A = 16'h0083; B = 16'h005D; #100;
A = 16'h0083; B = 16'h005E; #100;
A = 16'h0083; B = 16'h005F; #100;
A = 16'h0083; B = 16'h0060; #100;
A = 16'h0083; B = 16'h0061; #100;
A = 16'h0083; B = 16'h0062; #100;
A = 16'h0083; B = 16'h0063; #100;
A = 16'h0083; B = 16'h0064; #100;
A = 16'h0083; B = 16'h0065; #100;
A = 16'h0083; B = 16'h0066; #100;
A = 16'h0083; B = 16'h0067; #100;
A = 16'h0083; B = 16'h0068; #100;
A = 16'h0083; B = 16'h0069; #100;
A = 16'h0083; B = 16'h006A; #100;
A = 16'h0083; B = 16'h006B; #100;
A = 16'h0083; B = 16'h006C; #100;
A = 16'h0083; B = 16'h006D; #100;
A = 16'h0083; B = 16'h006E; #100;
A = 16'h0083; B = 16'h006F; #100;
A = 16'h0083; B = 16'h0070; #100;
A = 16'h0083; B = 16'h0071; #100;
A = 16'h0083; B = 16'h0072; #100;
A = 16'h0083; B = 16'h0073; #100;
A = 16'h0083; B = 16'h0074; #100;
A = 16'h0083; B = 16'h0075; #100;
A = 16'h0083; B = 16'h0076; #100;
A = 16'h0083; B = 16'h0077; #100;
A = 16'h0083; B = 16'h0078; #100;
A = 16'h0083; B = 16'h0079; #100;
A = 16'h0083; B = 16'h007A; #100;
A = 16'h0083; B = 16'h007B; #100;
A = 16'h0083; B = 16'h007C; #100;
A = 16'h0083; B = 16'h007D; #100;
A = 16'h0083; B = 16'h007E; #100;
A = 16'h0083; B = 16'h007F; #100;
A = 16'h0083; B = 16'h0080; #100;
A = 16'h0083; B = 16'h0081; #100;
A = 16'h0083; B = 16'h0082; #100;
A = 16'h0083; B = 16'h0083; #100;
A = 16'h0083; B = 16'h0084; #100;
A = 16'h0083; B = 16'h0085; #100;
A = 16'h0083; B = 16'h0086; #100;
A = 16'h0083; B = 16'h0087; #100;
A = 16'h0083; B = 16'h0088; #100;
A = 16'h0083; B = 16'h0089; #100;
A = 16'h0083; B = 16'h008A; #100;
A = 16'h0083; B = 16'h008B; #100;
A = 16'h0083; B = 16'h008C; #100;
A = 16'h0083; B = 16'h008D; #100;
A = 16'h0083; B = 16'h008E; #100;
A = 16'h0083; B = 16'h008F; #100;
A = 16'h0083; B = 16'h0090; #100;
A = 16'h0083; B = 16'h0091; #100;
A = 16'h0083; B = 16'h0092; #100;
A = 16'h0083; B = 16'h0093; #100;
A = 16'h0083; B = 16'h0094; #100;
A = 16'h0083; B = 16'h0095; #100;
A = 16'h0083; B = 16'h0096; #100;
A = 16'h0083; B = 16'h0097; #100;
A = 16'h0083; B = 16'h0098; #100;
A = 16'h0083; B = 16'h0099; #100;
A = 16'h0083; B = 16'h009A; #100;
A = 16'h0083; B = 16'h009B; #100;
A = 16'h0083; B = 16'h009C; #100;
A = 16'h0083; B = 16'h009D; #100;
A = 16'h0083; B = 16'h009E; #100;
A = 16'h0083; B = 16'h009F; #100;
A = 16'h0083; B = 16'h00A0; #100;
A = 16'h0083; B = 16'h00A1; #100;
A = 16'h0083; B = 16'h00A2; #100;
A = 16'h0083; B = 16'h00A3; #100;
A = 16'h0083; B = 16'h00A4; #100;
A = 16'h0083; B = 16'h00A5; #100;
A = 16'h0083; B = 16'h00A6; #100;
A = 16'h0083; B = 16'h00A7; #100;
A = 16'h0083; B = 16'h00A8; #100;
A = 16'h0083; B = 16'h00A9; #100;
A = 16'h0083; B = 16'h00AA; #100;
A = 16'h0083; B = 16'h00AB; #100;
A = 16'h0083; B = 16'h00AC; #100;
A = 16'h0083; B = 16'h00AD; #100;
A = 16'h0083; B = 16'h00AE; #100;
A = 16'h0083; B = 16'h00AF; #100;
A = 16'h0083; B = 16'h00B0; #100;
A = 16'h0083; B = 16'h00B1; #100;
A = 16'h0083; B = 16'h00B2; #100;
A = 16'h0083; B = 16'h00B3; #100;
A = 16'h0083; B = 16'h00B4; #100;
A = 16'h0083; B = 16'h00B5; #100;
A = 16'h0083; B = 16'h00B6; #100;
A = 16'h0083; B = 16'h00B7; #100;
A = 16'h0083; B = 16'h00B8; #100;
A = 16'h0083; B = 16'h00B9; #100;
A = 16'h0083; B = 16'h00BA; #100;
A = 16'h0083; B = 16'h00BB; #100;
A = 16'h0083; B = 16'h00BC; #100;
A = 16'h0083; B = 16'h00BD; #100;
A = 16'h0083; B = 16'h00BE; #100;
A = 16'h0083; B = 16'h00BF; #100;
A = 16'h0083; B = 16'h00C0; #100;
A = 16'h0083; B = 16'h00C1; #100;
A = 16'h0083; B = 16'h00C2; #100;
A = 16'h0083; B = 16'h00C3; #100;
A = 16'h0083; B = 16'h00C4; #100;
A = 16'h0083; B = 16'h00C5; #100;
A = 16'h0083; B = 16'h00C6; #100;
A = 16'h0083; B = 16'h00C7; #100;
A = 16'h0083; B = 16'h00C8; #100;
A = 16'h0083; B = 16'h00C9; #100;
A = 16'h0083; B = 16'h00CA; #100;
A = 16'h0083; B = 16'h00CB; #100;
A = 16'h0083; B = 16'h00CC; #100;
A = 16'h0083; B = 16'h00CD; #100;
A = 16'h0083; B = 16'h00CE; #100;
A = 16'h0083; B = 16'h00CF; #100;
A = 16'h0083; B = 16'h00D0; #100;
A = 16'h0083; B = 16'h00D1; #100;
A = 16'h0083; B = 16'h00D2; #100;
A = 16'h0083; B = 16'h00D3; #100;
A = 16'h0083; B = 16'h00D4; #100;
A = 16'h0083; B = 16'h00D5; #100;
A = 16'h0083; B = 16'h00D6; #100;
A = 16'h0083; B = 16'h00D7; #100;
A = 16'h0083; B = 16'h00D8; #100;
A = 16'h0083; B = 16'h00D9; #100;
A = 16'h0083; B = 16'h00DA; #100;
A = 16'h0083; B = 16'h00DB; #100;
A = 16'h0083; B = 16'h00DC; #100;
A = 16'h0083; B = 16'h00DD; #100;
A = 16'h0083; B = 16'h00DE; #100;
A = 16'h0083; B = 16'h00DF; #100;
A = 16'h0083; B = 16'h00E0; #100;
A = 16'h0083; B = 16'h00E1; #100;
A = 16'h0083; B = 16'h00E2; #100;
A = 16'h0083; B = 16'h00E3; #100;
A = 16'h0083; B = 16'h00E4; #100;
A = 16'h0083; B = 16'h00E5; #100;
A = 16'h0083; B = 16'h00E6; #100;
A = 16'h0083; B = 16'h00E7; #100;
A = 16'h0083; B = 16'h00E8; #100;
A = 16'h0083; B = 16'h00E9; #100;
A = 16'h0083; B = 16'h00EA; #100;
A = 16'h0083; B = 16'h00EB; #100;
A = 16'h0083; B = 16'h00EC; #100;
A = 16'h0083; B = 16'h00ED; #100;
A = 16'h0083; B = 16'h00EE; #100;
A = 16'h0083; B = 16'h00EF; #100;
A = 16'h0083; B = 16'h00F0; #100;
A = 16'h0083; B = 16'h00F1; #100;
A = 16'h0083; B = 16'h00F2; #100;
A = 16'h0083; B = 16'h00F3; #100;
A = 16'h0083; B = 16'h00F4; #100;
A = 16'h0083; B = 16'h00F5; #100;
A = 16'h0083; B = 16'h00F6; #100;
A = 16'h0083; B = 16'h00F7; #100;
A = 16'h0083; B = 16'h00F8; #100;
A = 16'h0083; B = 16'h00F9; #100;
A = 16'h0083; B = 16'h00FA; #100;
A = 16'h0083; B = 16'h00FB; #100;
A = 16'h0083; B = 16'h00FC; #100;
A = 16'h0083; B = 16'h00FD; #100;
A = 16'h0083; B = 16'h00FE; #100;
A = 16'h0083; B = 16'h00FF; #100;
A = 16'h0084; B = 16'h000; #100;
A = 16'h0084; B = 16'h001; #100;
A = 16'h0084; B = 16'h002; #100;
A = 16'h0084; B = 16'h003; #100;
A = 16'h0084; B = 16'h004; #100;
A = 16'h0084; B = 16'h005; #100;
A = 16'h0084; B = 16'h006; #100;
A = 16'h0084; B = 16'h007; #100;
A = 16'h0084; B = 16'h008; #100;
A = 16'h0084; B = 16'h009; #100;
A = 16'h0084; B = 16'h00A; #100;
A = 16'h0084; B = 16'h00B; #100;
A = 16'h0084; B = 16'h00C; #100;
A = 16'h0084; B = 16'h00D; #100;
A = 16'h0084; B = 16'h00E; #100;
A = 16'h0084; B = 16'h00F; #100;
A = 16'h0084; B = 16'h0010; #100;
A = 16'h0084; B = 16'h0011; #100;
A = 16'h0084; B = 16'h0012; #100;
A = 16'h0084; B = 16'h0013; #100;
A = 16'h0084; B = 16'h0014; #100;
A = 16'h0084; B = 16'h0015; #100;
A = 16'h0084; B = 16'h0016; #100;
A = 16'h0084; B = 16'h0017; #100;
A = 16'h0084; B = 16'h0018; #100;
A = 16'h0084; B = 16'h0019; #100;
A = 16'h0084; B = 16'h001A; #100;
A = 16'h0084; B = 16'h001B; #100;
A = 16'h0084; B = 16'h001C; #100;
A = 16'h0084; B = 16'h001D; #100;
A = 16'h0084; B = 16'h001E; #100;
A = 16'h0084; B = 16'h001F; #100;
A = 16'h0084; B = 16'h0020; #100;
A = 16'h0084; B = 16'h0021; #100;
A = 16'h0084; B = 16'h0022; #100;
A = 16'h0084; B = 16'h0023; #100;
A = 16'h0084; B = 16'h0024; #100;
A = 16'h0084; B = 16'h0025; #100;
A = 16'h0084; B = 16'h0026; #100;
A = 16'h0084; B = 16'h0027; #100;
A = 16'h0084; B = 16'h0028; #100;
A = 16'h0084; B = 16'h0029; #100;
A = 16'h0084; B = 16'h002A; #100;
A = 16'h0084; B = 16'h002B; #100;
A = 16'h0084; B = 16'h002C; #100;
A = 16'h0084; B = 16'h002D; #100;
A = 16'h0084; B = 16'h002E; #100;
A = 16'h0084; B = 16'h002F; #100;
A = 16'h0084; B = 16'h0030; #100;
A = 16'h0084; B = 16'h0031; #100;
A = 16'h0084; B = 16'h0032; #100;
A = 16'h0084; B = 16'h0033; #100;
A = 16'h0084; B = 16'h0034; #100;
A = 16'h0084; B = 16'h0035; #100;
A = 16'h0084; B = 16'h0036; #100;
A = 16'h0084; B = 16'h0037; #100;
A = 16'h0084; B = 16'h0038; #100;
A = 16'h0084; B = 16'h0039; #100;
A = 16'h0084; B = 16'h003A; #100;
A = 16'h0084; B = 16'h003B; #100;
A = 16'h0084; B = 16'h003C; #100;
A = 16'h0084; B = 16'h003D; #100;
A = 16'h0084; B = 16'h003E; #100;
A = 16'h0084; B = 16'h003F; #100;
A = 16'h0084; B = 16'h0040; #100;
A = 16'h0084; B = 16'h0041; #100;
A = 16'h0084; B = 16'h0042; #100;
A = 16'h0084; B = 16'h0043; #100;
A = 16'h0084; B = 16'h0044; #100;
A = 16'h0084; B = 16'h0045; #100;
A = 16'h0084; B = 16'h0046; #100;
A = 16'h0084; B = 16'h0047; #100;
A = 16'h0084; B = 16'h0048; #100;
A = 16'h0084; B = 16'h0049; #100;
A = 16'h0084; B = 16'h004A; #100;
A = 16'h0084; B = 16'h004B; #100;
A = 16'h0084; B = 16'h004C; #100;
A = 16'h0084; B = 16'h004D; #100;
A = 16'h0084; B = 16'h004E; #100;
A = 16'h0084; B = 16'h004F; #100;
A = 16'h0084; B = 16'h0050; #100;
A = 16'h0084; B = 16'h0051; #100;
A = 16'h0084; B = 16'h0052; #100;
A = 16'h0084; B = 16'h0053; #100;
A = 16'h0084; B = 16'h0054; #100;
A = 16'h0084; B = 16'h0055; #100;
A = 16'h0084; B = 16'h0056; #100;
A = 16'h0084; B = 16'h0057; #100;
A = 16'h0084; B = 16'h0058; #100;
A = 16'h0084; B = 16'h0059; #100;
A = 16'h0084; B = 16'h005A; #100;
A = 16'h0084; B = 16'h005B; #100;
A = 16'h0084; B = 16'h005C; #100;
A = 16'h0084; B = 16'h005D; #100;
A = 16'h0084; B = 16'h005E; #100;
A = 16'h0084; B = 16'h005F; #100;
A = 16'h0084; B = 16'h0060; #100;
A = 16'h0084; B = 16'h0061; #100;
A = 16'h0084; B = 16'h0062; #100;
A = 16'h0084; B = 16'h0063; #100;
A = 16'h0084; B = 16'h0064; #100;
A = 16'h0084; B = 16'h0065; #100;
A = 16'h0084; B = 16'h0066; #100;
A = 16'h0084; B = 16'h0067; #100;
A = 16'h0084; B = 16'h0068; #100;
A = 16'h0084; B = 16'h0069; #100;
A = 16'h0084; B = 16'h006A; #100;
A = 16'h0084; B = 16'h006B; #100;
A = 16'h0084; B = 16'h006C; #100;
A = 16'h0084; B = 16'h006D; #100;
A = 16'h0084; B = 16'h006E; #100;
A = 16'h0084; B = 16'h006F; #100;
A = 16'h0084; B = 16'h0070; #100;
A = 16'h0084; B = 16'h0071; #100;
A = 16'h0084; B = 16'h0072; #100;
A = 16'h0084; B = 16'h0073; #100;
A = 16'h0084; B = 16'h0074; #100;
A = 16'h0084; B = 16'h0075; #100;
A = 16'h0084; B = 16'h0076; #100;
A = 16'h0084; B = 16'h0077; #100;
A = 16'h0084; B = 16'h0078; #100;
A = 16'h0084; B = 16'h0079; #100;
A = 16'h0084; B = 16'h007A; #100;
A = 16'h0084; B = 16'h007B; #100;
A = 16'h0084; B = 16'h007C; #100;
A = 16'h0084; B = 16'h007D; #100;
A = 16'h0084; B = 16'h007E; #100;
A = 16'h0084; B = 16'h007F; #100;
A = 16'h0084; B = 16'h0080; #100;
A = 16'h0084; B = 16'h0081; #100;
A = 16'h0084; B = 16'h0082; #100;
A = 16'h0084; B = 16'h0083; #100;
A = 16'h0084; B = 16'h0084; #100;
A = 16'h0084; B = 16'h0085; #100;
A = 16'h0084; B = 16'h0086; #100;
A = 16'h0084; B = 16'h0087; #100;
A = 16'h0084; B = 16'h0088; #100;
A = 16'h0084; B = 16'h0089; #100;
A = 16'h0084; B = 16'h008A; #100;
A = 16'h0084; B = 16'h008B; #100;
A = 16'h0084; B = 16'h008C; #100;
A = 16'h0084; B = 16'h008D; #100;
A = 16'h0084; B = 16'h008E; #100;
A = 16'h0084; B = 16'h008F; #100;
A = 16'h0084; B = 16'h0090; #100;
A = 16'h0084; B = 16'h0091; #100;
A = 16'h0084; B = 16'h0092; #100;
A = 16'h0084; B = 16'h0093; #100;
A = 16'h0084; B = 16'h0094; #100;
A = 16'h0084; B = 16'h0095; #100;
A = 16'h0084; B = 16'h0096; #100;
A = 16'h0084; B = 16'h0097; #100;
A = 16'h0084; B = 16'h0098; #100;
A = 16'h0084; B = 16'h0099; #100;
A = 16'h0084; B = 16'h009A; #100;
A = 16'h0084; B = 16'h009B; #100;
A = 16'h0084; B = 16'h009C; #100;
A = 16'h0084; B = 16'h009D; #100;
A = 16'h0084; B = 16'h009E; #100;
A = 16'h0084; B = 16'h009F; #100;
A = 16'h0084; B = 16'h00A0; #100;
A = 16'h0084; B = 16'h00A1; #100;
A = 16'h0084; B = 16'h00A2; #100;
A = 16'h0084; B = 16'h00A3; #100;
A = 16'h0084; B = 16'h00A4; #100;
A = 16'h0084; B = 16'h00A5; #100;
A = 16'h0084; B = 16'h00A6; #100;
A = 16'h0084; B = 16'h00A7; #100;
A = 16'h0084; B = 16'h00A8; #100;
A = 16'h0084; B = 16'h00A9; #100;
A = 16'h0084; B = 16'h00AA; #100;
A = 16'h0084; B = 16'h00AB; #100;
A = 16'h0084; B = 16'h00AC; #100;
A = 16'h0084; B = 16'h00AD; #100;
A = 16'h0084; B = 16'h00AE; #100;
A = 16'h0084; B = 16'h00AF; #100;
A = 16'h0084; B = 16'h00B0; #100;
A = 16'h0084; B = 16'h00B1; #100;
A = 16'h0084; B = 16'h00B2; #100;
A = 16'h0084; B = 16'h00B3; #100;
A = 16'h0084; B = 16'h00B4; #100;
A = 16'h0084; B = 16'h00B5; #100;
A = 16'h0084; B = 16'h00B6; #100;
A = 16'h0084; B = 16'h00B7; #100;
A = 16'h0084; B = 16'h00B8; #100;
A = 16'h0084; B = 16'h00B9; #100;
A = 16'h0084; B = 16'h00BA; #100;
A = 16'h0084; B = 16'h00BB; #100;
A = 16'h0084; B = 16'h00BC; #100;
A = 16'h0084; B = 16'h00BD; #100;
A = 16'h0084; B = 16'h00BE; #100;
A = 16'h0084; B = 16'h00BF; #100;
A = 16'h0084; B = 16'h00C0; #100;
A = 16'h0084; B = 16'h00C1; #100;
A = 16'h0084; B = 16'h00C2; #100;
A = 16'h0084; B = 16'h00C3; #100;
A = 16'h0084; B = 16'h00C4; #100;
A = 16'h0084; B = 16'h00C5; #100;
A = 16'h0084; B = 16'h00C6; #100;
A = 16'h0084; B = 16'h00C7; #100;
A = 16'h0084; B = 16'h00C8; #100;
A = 16'h0084; B = 16'h00C9; #100;
A = 16'h0084; B = 16'h00CA; #100;
A = 16'h0084; B = 16'h00CB; #100;
A = 16'h0084; B = 16'h00CC; #100;
A = 16'h0084; B = 16'h00CD; #100;
A = 16'h0084; B = 16'h00CE; #100;
A = 16'h0084; B = 16'h00CF; #100;
A = 16'h0084; B = 16'h00D0; #100;
A = 16'h0084; B = 16'h00D1; #100;
A = 16'h0084; B = 16'h00D2; #100;
A = 16'h0084; B = 16'h00D3; #100;
A = 16'h0084; B = 16'h00D4; #100;
A = 16'h0084; B = 16'h00D5; #100;
A = 16'h0084; B = 16'h00D6; #100;
A = 16'h0084; B = 16'h00D7; #100;
A = 16'h0084; B = 16'h00D8; #100;
A = 16'h0084; B = 16'h00D9; #100;
A = 16'h0084; B = 16'h00DA; #100;
A = 16'h0084; B = 16'h00DB; #100;
A = 16'h0084; B = 16'h00DC; #100;
A = 16'h0084; B = 16'h00DD; #100;
A = 16'h0084; B = 16'h00DE; #100;
A = 16'h0084; B = 16'h00DF; #100;
A = 16'h0084; B = 16'h00E0; #100;
A = 16'h0084; B = 16'h00E1; #100;
A = 16'h0084; B = 16'h00E2; #100;
A = 16'h0084; B = 16'h00E3; #100;
A = 16'h0084; B = 16'h00E4; #100;
A = 16'h0084; B = 16'h00E5; #100;
A = 16'h0084; B = 16'h00E6; #100;
A = 16'h0084; B = 16'h00E7; #100;
A = 16'h0084; B = 16'h00E8; #100;
A = 16'h0084; B = 16'h00E9; #100;
A = 16'h0084; B = 16'h00EA; #100;
A = 16'h0084; B = 16'h00EB; #100;
A = 16'h0084; B = 16'h00EC; #100;
A = 16'h0084; B = 16'h00ED; #100;
A = 16'h0084; B = 16'h00EE; #100;
A = 16'h0084; B = 16'h00EF; #100;
A = 16'h0084; B = 16'h00F0; #100;
A = 16'h0084; B = 16'h00F1; #100;
A = 16'h0084; B = 16'h00F2; #100;
A = 16'h0084; B = 16'h00F3; #100;
A = 16'h0084; B = 16'h00F4; #100;
A = 16'h0084; B = 16'h00F5; #100;
A = 16'h0084; B = 16'h00F6; #100;
A = 16'h0084; B = 16'h00F7; #100;
A = 16'h0084; B = 16'h00F8; #100;
A = 16'h0084; B = 16'h00F9; #100;
A = 16'h0084; B = 16'h00FA; #100;
A = 16'h0084; B = 16'h00FB; #100;
A = 16'h0084; B = 16'h00FC; #100;
A = 16'h0084; B = 16'h00FD; #100;
A = 16'h0084; B = 16'h00FE; #100;
A = 16'h0084; B = 16'h00FF; #100;
A = 16'h0085; B = 16'h000; #100;
A = 16'h0085; B = 16'h001; #100;
A = 16'h0085; B = 16'h002; #100;
A = 16'h0085; B = 16'h003; #100;
A = 16'h0085; B = 16'h004; #100;
A = 16'h0085; B = 16'h005; #100;
A = 16'h0085; B = 16'h006; #100;
A = 16'h0085; B = 16'h007; #100;
A = 16'h0085; B = 16'h008; #100;
A = 16'h0085; B = 16'h009; #100;
A = 16'h0085; B = 16'h00A; #100;
A = 16'h0085; B = 16'h00B; #100;
A = 16'h0085; B = 16'h00C; #100;
A = 16'h0085; B = 16'h00D; #100;
A = 16'h0085; B = 16'h00E; #100;
A = 16'h0085; B = 16'h00F; #100;
A = 16'h0085; B = 16'h0010; #100;
A = 16'h0085; B = 16'h0011; #100;
A = 16'h0085; B = 16'h0012; #100;
A = 16'h0085; B = 16'h0013; #100;
A = 16'h0085; B = 16'h0014; #100;
A = 16'h0085; B = 16'h0015; #100;
A = 16'h0085; B = 16'h0016; #100;
A = 16'h0085; B = 16'h0017; #100;
A = 16'h0085; B = 16'h0018; #100;
A = 16'h0085; B = 16'h0019; #100;
A = 16'h0085; B = 16'h001A; #100;
A = 16'h0085; B = 16'h001B; #100;
A = 16'h0085; B = 16'h001C; #100;
A = 16'h0085; B = 16'h001D; #100;
A = 16'h0085; B = 16'h001E; #100;
A = 16'h0085; B = 16'h001F; #100;
A = 16'h0085; B = 16'h0020; #100;
A = 16'h0085; B = 16'h0021; #100;
A = 16'h0085; B = 16'h0022; #100;
A = 16'h0085; B = 16'h0023; #100;
A = 16'h0085; B = 16'h0024; #100;
A = 16'h0085; B = 16'h0025; #100;
A = 16'h0085; B = 16'h0026; #100;
A = 16'h0085; B = 16'h0027; #100;
A = 16'h0085; B = 16'h0028; #100;
A = 16'h0085; B = 16'h0029; #100;
A = 16'h0085; B = 16'h002A; #100;
A = 16'h0085; B = 16'h002B; #100;
A = 16'h0085; B = 16'h002C; #100;
A = 16'h0085; B = 16'h002D; #100;
A = 16'h0085; B = 16'h002E; #100;
A = 16'h0085; B = 16'h002F; #100;
A = 16'h0085; B = 16'h0030; #100;
A = 16'h0085; B = 16'h0031; #100;
A = 16'h0085; B = 16'h0032; #100;
A = 16'h0085; B = 16'h0033; #100;
A = 16'h0085; B = 16'h0034; #100;
A = 16'h0085; B = 16'h0035; #100;
A = 16'h0085; B = 16'h0036; #100;
A = 16'h0085; B = 16'h0037; #100;
A = 16'h0085; B = 16'h0038; #100;
A = 16'h0085; B = 16'h0039; #100;
A = 16'h0085; B = 16'h003A; #100;
A = 16'h0085; B = 16'h003B; #100;
A = 16'h0085; B = 16'h003C; #100;
A = 16'h0085; B = 16'h003D; #100;
A = 16'h0085; B = 16'h003E; #100;
A = 16'h0085; B = 16'h003F; #100;
A = 16'h0085; B = 16'h0040; #100;
A = 16'h0085; B = 16'h0041; #100;
A = 16'h0085; B = 16'h0042; #100;
A = 16'h0085; B = 16'h0043; #100;
A = 16'h0085; B = 16'h0044; #100;
A = 16'h0085; B = 16'h0045; #100;
A = 16'h0085; B = 16'h0046; #100;
A = 16'h0085; B = 16'h0047; #100;
A = 16'h0085; B = 16'h0048; #100;
A = 16'h0085; B = 16'h0049; #100;
A = 16'h0085; B = 16'h004A; #100;
A = 16'h0085; B = 16'h004B; #100;
A = 16'h0085; B = 16'h004C; #100;
A = 16'h0085; B = 16'h004D; #100;
A = 16'h0085; B = 16'h004E; #100;
A = 16'h0085; B = 16'h004F; #100;
A = 16'h0085; B = 16'h0050; #100;
A = 16'h0085; B = 16'h0051; #100;
A = 16'h0085; B = 16'h0052; #100;
A = 16'h0085; B = 16'h0053; #100;
A = 16'h0085; B = 16'h0054; #100;
A = 16'h0085; B = 16'h0055; #100;
A = 16'h0085; B = 16'h0056; #100;
A = 16'h0085; B = 16'h0057; #100;
A = 16'h0085; B = 16'h0058; #100;
A = 16'h0085; B = 16'h0059; #100;
A = 16'h0085; B = 16'h005A; #100;
A = 16'h0085; B = 16'h005B; #100;
A = 16'h0085; B = 16'h005C; #100;
A = 16'h0085; B = 16'h005D; #100;
A = 16'h0085; B = 16'h005E; #100;
A = 16'h0085; B = 16'h005F; #100;
A = 16'h0085; B = 16'h0060; #100;
A = 16'h0085; B = 16'h0061; #100;
A = 16'h0085; B = 16'h0062; #100;
A = 16'h0085; B = 16'h0063; #100;
A = 16'h0085; B = 16'h0064; #100;
A = 16'h0085; B = 16'h0065; #100;
A = 16'h0085; B = 16'h0066; #100;
A = 16'h0085; B = 16'h0067; #100;
A = 16'h0085; B = 16'h0068; #100;
A = 16'h0085; B = 16'h0069; #100;
A = 16'h0085; B = 16'h006A; #100;
A = 16'h0085; B = 16'h006B; #100;
A = 16'h0085; B = 16'h006C; #100;
A = 16'h0085; B = 16'h006D; #100;
A = 16'h0085; B = 16'h006E; #100;
A = 16'h0085; B = 16'h006F; #100;
A = 16'h0085; B = 16'h0070; #100;
A = 16'h0085; B = 16'h0071; #100;
A = 16'h0085; B = 16'h0072; #100;
A = 16'h0085; B = 16'h0073; #100;
A = 16'h0085; B = 16'h0074; #100;
A = 16'h0085; B = 16'h0075; #100;
A = 16'h0085; B = 16'h0076; #100;
A = 16'h0085; B = 16'h0077; #100;
A = 16'h0085; B = 16'h0078; #100;
A = 16'h0085; B = 16'h0079; #100;
A = 16'h0085; B = 16'h007A; #100;
A = 16'h0085; B = 16'h007B; #100;
A = 16'h0085; B = 16'h007C; #100;
A = 16'h0085; B = 16'h007D; #100;
A = 16'h0085; B = 16'h007E; #100;
A = 16'h0085; B = 16'h007F; #100;
A = 16'h0085; B = 16'h0080; #100;
A = 16'h0085; B = 16'h0081; #100;
A = 16'h0085; B = 16'h0082; #100;
A = 16'h0085; B = 16'h0083; #100;
A = 16'h0085; B = 16'h0084; #100;
A = 16'h0085; B = 16'h0085; #100;
A = 16'h0085; B = 16'h0086; #100;
A = 16'h0085; B = 16'h0087; #100;
A = 16'h0085; B = 16'h0088; #100;
A = 16'h0085; B = 16'h0089; #100;
A = 16'h0085; B = 16'h008A; #100;
A = 16'h0085; B = 16'h008B; #100;
A = 16'h0085; B = 16'h008C; #100;
A = 16'h0085; B = 16'h008D; #100;
A = 16'h0085; B = 16'h008E; #100;
A = 16'h0085; B = 16'h008F; #100;
A = 16'h0085; B = 16'h0090; #100;
A = 16'h0085; B = 16'h0091; #100;
A = 16'h0085; B = 16'h0092; #100;
A = 16'h0085; B = 16'h0093; #100;
A = 16'h0085; B = 16'h0094; #100;
A = 16'h0085; B = 16'h0095; #100;
A = 16'h0085; B = 16'h0096; #100;
A = 16'h0085; B = 16'h0097; #100;
A = 16'h0085; B = 16'h0098; #100;
A = 16'h0085; B = 16'h0099; #100;
A = 16'h0085; B = 16'h009A; #100;
A = 16'h0085; B = 16'h009B; #100;
A = 16'h0085; B = 16'h009C; #100;
A = 16'h0085; B = 16'h009D; #100;
A = 16'h0085; B = 16'h009E; #100;
A = 16'h0085; B = 16'h009F; #100;
A = 16'h0085; B = 16'h00A0; #100;
A = 16'h0085; B = 16'h00A1; #100;
A = 16'h0085; B = 16'h00A2; #100;
A = 16'h0085; B = 16'h00A3; #100;
A = 16'h0085; B = 16'h00A4; #100;
A = 16'h0085; B = 16'h00A5; #100;
A = 16'h0085; B = 16'h00A6; #100;
A = 16'h0085; B = 16'h00A7; #100;
A = 16'h0085; B = 16'h00A8; #100;
A = 16'h0085; B = 16'h00A9; #100;
A = 16'h0085; B = 16'h00AA; #100;
A = 16'h0085; B = 16'h00AB; #100;
A = 16'h0085; B = 16'h00AC; #100;
A = 16'h0085; B = 16'h00AD; #100;
A = 16'h0085; B = 16'h00AE; #100;
A = 16'h0085; B = 16'h00AF; #100;
A = 16'h0085; B = 16'h00B0; #100;
A = 16'h0085; B = 16'h00B1; #100;
A = 16'h0085; B = 16'h00B2; #100;
A = 16'h0085; B = 16'h00B3; #100;
A = 16'h0085; B = 16'h00B4; #100;
A = 16'h0085; B = 16'h00B5; #100;
A = 16'h0085; B = 16'h00B6; #100;
A = 16'h0085; B = 16'h00B7; #100;
A = 16'h0085; B = 16'h00B8; #100;
A = 16'h0085; B = 16'h00B9; #100;
A = 16'h0085; B = 16'h00BA; #100;
A = 16'h0085; B = 16'h00BB; #100;
A = 16'h0085; B = 16'h00BC; #100;
A = 16'h0085; B = 16'h00BD; #100;
A = 16'h0085; B = 16'h00BE; #100;
A = 16'h0085; B = 16'h00BF; #100;
A = 16'h0085; B = 16'h00C0; #100;
A = 16'h0085; B = 16'h00C1; #100;
A = 16'h0085; B = 16'h00C2; #100;
A = 16'h0085; B = 16'h00C3; #100;
A = 16'h0085; B = 16'h00C4; #100;
A = 16'h0085; B = 16'h00C5; #100;
A = 16'h0085; B = 16'h00C6; #100;
A = 16'h0085; B = 16'h00C7; #100;
A = 16'h0085; B = 16'h00C8; #100;
A = 16'h0085; B = 16'h00C9; #100;
A = 16'h0085; B = 16'h00CA; #100;
A = 16'h0085; B = 16'h00CB; #100;
A = 16'h0085; B = 16'h00CC; #100;
A = 16'h0085; B = 16'h00CD; #100;
A = 16'h0085; B = 16'h00CE; #100;
A = 16'h0085; B = 16'h00CF; #100;
A = 16'h0085; B = 16'h00D0; #100;
A = 16'h0085; B = 16'h00D1; #100;
A = 16'h0085; B = 16'h00D2; #100;
A = 16'h0085; B = 16'h00D3; #100;
A = 16'h0085; B = 16'h00D4; #100;
A = 16'h0085; B = 16'h00D5; #100;
A = 16'h0085; B = 16'h00D6; #100;
A = 16'h0085; B = 16'h00D7; #100;
A = 16'h0085; B = 16'h00D8; #100;
A = 16'h0085; B = 16'h00D9; #100;
A = 16'h0085; B = 16'h00DA; #100;
A = 16'h0085; B = 16'h00DB; #100;
A = 16'h0085; B = 16'h00DC; #100;
A = 16'h0085; B = 16'h00DD; #100;
A = 16'h0085; B = 16'h00DE; #100;
A = 16'h0085; B = 16'h00DF; #100;
A = 16'h0085; B = 16'h00E0; #100;
A = 16'h0085; B = 16'h00E1; #100;
A = 16'h0085; B = 16'h00E2; #100;
A = 16'h0085; B = 16'h00E3; #100;
A = 16'h0085; B = 16'h00E4; #100;
A = 16'h0085; B = 16'h00E5; #100;
A = 16'h0085; B = 16'h00E6; #100;
A = 16'h0085; B = 16'h00E7; #100;
A = 16'h0085; B = 16'h00E8; #100;
A = 16'h0085; B = 16'h00E9; #100;
A = 16'h0085; B = 16'h00EA; #100;
A = 16'h0085; B = 16'h00EB; #100;
A = 16'h0085; B = 16'h00EC; #100;
A = 16'h0085; B = 16'h00ED; #100;
A = 16'h0085; B = 16'h00EE; #100;
A = 16'h0085; B = 16'h00EF; #100;
A = 16'h0085; B = 16'h00F0; #100;
A = 16'h0085; B = 16'h00F1; #100;
A = 16'h0085; B = 16'h00F2; #100;
A = 16'h0085; B = 16'h00F3; #100;
A = 16'h0085; B = 16'h00F4; #100;
A = 16'h0085; B = 16'h00F5; #100;
A = 16'h0085; B = 16'h00F6; #100;
A = 16'h0085; B = 16'h00F7; #100;
A = 16'h0085; B = 16'h00F8; #100;
A = 16'h0085; B = 16'h00F9; #100;
A = 16'h0085; B = 16'h00FA; #100;
A = 16'h0085; B = 16'h00FB; #100;
A = 16'h0085; B = 16'h00FC; #100;
A = 16'h0085; B = 16'h00FD; #100;
A = 16'h0085; B = 16'h00FE; #100;
A = 16'h0085; B = 16'h00FF; #100;
A = 16'h0086; B = 16'h000; #100;
A = 16'h0086; B = 16'h001; #100;
A = 16'h0086; B = 16'h002; #100;
A = 16'h0086; B = 16'h003; #100;
A = 16'h0086; B = 16'h004; #100;
A = 16'h0086; B = 16'h005; #100;
A = 16'h0086; B = 16'h006; #100;
A = 16'h0086; B = 16'h007; #100;
A = 16'h0086; B = 16'h008; #100;
A = 16'h0086; B = 16'h009; #100;
A = 16'h0086; B = 16'h00A; #100;
A = 16'h0086; B = 16'h00B; #100;
A = 16'h0086; B = 16'h00C; #100;
A = 16'h0086; B = 16'h00D; #100;
A = 16'h0086; B = 16'h00E; #100;
A = 16'h0086; B = 16'h00F; #100;
A = 16'h0086; B = 16'h0010; #100;
A = 16'h0086; B = 16'h0011; #100;
A = 16'h0086; B = 16'h0012; #100;
A = 16'h0086; B = 16'h0013; #100;
A = 16'h0086; B = 16'h0014; #100;
A = 16'h0086; B = 16'h0015; #100;
A = 16'h0086; B = 16'h0016; #100;
A = 16'h0086; B = 16'h0017; #100;
A = 16'h0086; B = 16'h0018; #100;
A = 16'h0086; B = 16'h0019; #100;
A = 16'h0086; B = 16'h001A; #100;
A = 16'h0086; B = 16'h001B; #100;
A = 16'h0086; B = 16'h001C; #100;
A = 16'h0086; B = 16'h001D; #100;
A = 16'h0086; B = 16'h001E; #100;
A = 16'h0086; B = 16'h001F; #100;
A = 16'h0086; B = 16'h0020; #100;
A = 16'h0086; B = 16'h0021; #100;
A = 16'h0086; B = 16'h0022; #100;
A = 16'h0086; B = 16'h0023; #100;
A = 16'h0086; B = 16'h0024; #100;
A = 16'h0086; B = 16'h0025; #100;
A = 16'h0086; B = 16'h0026; #100;
A = 16'h0086; B = 16'h0027; #100;
A = 16'h0086; B = 16'h0028; #100;
A = 16'h0086; B = 16'h0029; #100;
A = 16'h0086; B = 16'h002A; #100;
A = 16'h0086; B = 16'h002B; #100;
A = 16'h0086; B = 16'h002C; #100;
A = 16'h0086; B = 16'h002D; #100;
A = 16'h0086; B = 16'h002E; #100;
A = 16'h0086; B = 16'h002F; #100;
A = 16'h0086; B = 16'h0030; #100;
A = 16'h0086; B = 16'h0031; #100;
A = 16'h0086; B = 16'h0032; #100;
A = 16'h0086; B = 16'h0033; #100;
A = 16'h0086; B = 16'h0034; #100;
A = 16'h0086; B = 16'h0035; #100;
A = 16'h0086; B = 16'h0036; #100;
A = 16'h0086; B = 16'h0037; #100;
A = 16'h0086; B = 16'h0038; #100;
A = 16'h0086; B = 16'h0039; #100;
A = 16'h0086; B = 16'h003A; #100;
A = 16'h0086; B = 16'h003B; #100;
A = 16'h0086; B = 16'h003C; #100;
A = 16'h0086; B = 16'h003D; #100;
A = 16'h0086; B = 16'h003E; #100;
A = 16'h0086; B = 16'h003F; #100;
A = 16'h0086; B = 16'h0040; #100;
A = 16'h0086; B = 16'h0041; #100;
A = 16'h0086; B = 16'h0042; #100;
A = 16'h0086; B = 16'h0043; #100;
A = 16'h0086; B = 16'h0044; #100;
A = 16'h0086; B = 16'h0045; #100;
A = 16'h0086; B = 16'h0046; #100;
A = 16'h0086; B = 16'h0047; #100;
A = 16'h0086; B = 16'h0048; #100;
A = 16'h0086; B = 16'h0049; #100;
A = 16'h0086; B = 16'h004A; #100;
A = 16'h0086; B = 16'h004B; #100;
A = 16'h0086; B = 16'h004C; #100;
A = 16'h0086; B = 16'h004D; #100;
A = 16'h0086; B = 16'h004E; #100;
A = 16'h0086; B = 16'h004F; #100;
A = 16'h0086; B = 16'h0050; #100;
A = 16'h0086; B = 16'h0051; #100;
A = 16'h0086; B = 16'h0052; #100;
A = 16'h0086; B = 16'h0053; #100;
A = 16'h0086; B = 16'h0054; #100;
A = 16'h0086; B = 16'h0055; #100;
A = 16'h0086; B = 16'h0056; #100;
A = 16'h0086; B = 16'h0057; #100;
A = 16'h0086; B = 16'h0058; #100;
A = 16'h0086; B = 16'h0059; #100;
A = 16'h0086; B = 16'h005A; #100;
A = 16'h0086; B = 16'h005B; #100;
A = 16'h0086; B = 16'h005C; #100;
A = 16'h0086; B = 16'h005D; #100;
A = 16'h0086; B = 16'h005E; #100;
A = 16'h0086; B = 16'h005F; #100;
A = 16'h0086; B = 16'h0060; #100;
A = 16'h0086; B = 16'h0061; #100;
A = 16'h0086; B = 16'h0062; #100;
A = 16'h0086; B = 16'h0063; #100;
A = 16'h0086; B = 16'h0064; #100;
A = 16'h0086; B = 16'h0065; #100;
A = 16'h0086; B = 16'h0066; #100;
A = 16'h0086; B = 16'h0067; #100;
A = 16'h0086; B = 16'h0068; #100;
A = 16'h0086; B = 16'h0069; #100;
A = 16'h0086; B = 16'h006A; #100;
A = 16'h0086; B = 16'h006B; #100;
A = 16'h0086; B = 16'h006C; #100;
A = 16'h0086; B = 16'h006D; #100;
A = 16'h0086; B = 16'h006E; #100;
A = 16'h0086; B = 16'h006F; #100;
A = 16'h0086; B = 16'h0070; #100;
A = 16'h0086; B = 16'h0071; #100;
A = 16'h0086; B = 16'h0072; #100;
A = 16'h0086; B = 16'h0073; #100;
A = 16'h0086; B = 16'h0074; #100;
A = 16'h0086; B = 16'h0075; #100;
A = 16'h0086; B = 16'h0076; #100;
A = 16'h0086; B = 16'h0077; #100;
A = 16'h0086; B = 16'h0078; #100;
A = 16'h0086; B = 16'h0079; #100;
A = 16'h0086; B = 16'h007A; #100;
A = 16'h0086; B = 16'h007B; #100;
A = 16'h0086; B = 16'h007C; #100;
A = 16'h0086; B = 16'h007D; #100;
A = 16'h0086; B = 16'h007E; #100;
A = 16'h0086; B = 16'h007F; #100;
A = 16'h0086; B = 16'h0080; #100;
A = 16'h0086; B = 16'h0081; #100;
A = 16'h0086; B = 16'h0082; #100;
A = 16'h0086; B = 16'h0083; #100;
A = 16'h0086; B = 16'h0084; #100;
A = 16'h0086; B = 16'h0085; #100;
A = 16'h0086; B = 16'h0086; #100;
A = 16'h0086; B = 16'h0087; #100;
A = 16'h0086; B = 16'h0088; #100;
A = 16'h0086; B = 16'h0089; #100;
A = 16'h0086; B = 16'h008A; #100;
A = 16'h0086; B = 16'h008B; #100;
A = 16'h0086; B = 16'h008C; #100;
A = 16'h0086; B = 16'h008D; #100;
A = 16'h0086; B = 16'h008E; #100;
A = 16'h0086; B = 16'h008F; #100;
A = 16'h0086; B = 16'h0090; #100;
A = 16'h0086; B = 16'h0091; #100;
A = 16'h0086; B = 16'h0092; #100;
A = 16'h0086; B = 16'h0093; #100;
A = 16'h0086; B = 16'h0094; #100;
A = 16'h0086; B = 16'h0095; #100;
A = 16'h0086; B = 16'h0096; #100;
A = 16'h0086; B = 16'h0097; #100;
A = 16'h0086; B = 16'h0098; #100;
A = 16'h0086; B = 16'h0099; #100;
A = 16'h0086; B = 16'h009A; #100;
A = 16'h0086; B = 16'h009B; #100;
A = 16'h0086; B = 16'h009C; #100;
A = 16'h0086; B = 16'h009D; #100;
A = 16'h0086; B = 16'h009E; #100;
A = 16'h0086; B = 16'h009F; #100;
A = 16'h0086; B = 16'h00A0; #100;
A = 16'h0086; B = 16'h00A1; #100;
A = 16'h0086; B = 16'h00A2; #100;
A = 16'h0086; B = 16'h00A3; #100;
A = 16'h0086; B = 16'h00A4; #100;
A = 16'h0086; B = 16'h00A5; #100;
A = 16'h0086; B = 16'h00A6; #100;
A = 16'h0086; B = 16'h00A7; #100;
A = 16'h0086; B = 16'h00A8; #100;
A = 16'h0086; B = 16'h00A9; #100;
A = 16'h0086; B = 16'h00AA; #100;
A = 16'h0086; B = 16'h00AB; #100;
A = 16'h0086; B = 16'h00AC; #100;
A = 16'h0086; B = 16'h00AD; #100;
A = 16'h0086; B = 16'h00AE; #100;
A = 16'h0086; B = 16'h00AF; #100;
A = 16'h0086; B = 16'h00B0; #100;
A = 16'h0086; B = 16'h00B1; #100;
A = 16'h0086; B = 16'h00B2; #100;
A = 16'h0086; B = 16'h00B3; #100;
A = 16'h0086; B = 16'h00B4; #100;
A = 16'h0086; B = 16'h00B5; #100;
A = 16'h0086; B = 16'h00B6; #100;
A = 16'h0086; B = 16'h00B7; #100;
A = 16'h0086; B = 16'h00B8; #100;
A = 16'h0086; B = 16'h00B9; #100;
A = 16'h0086; B = 16'h00BA; #100;
A = 16'h0086; B = 16'h00BB; #100;
A = 16'h0086; B = 16'h00BC; #100;
A = 16'h0086; B = 16'h00BD; #100;
A = 16'h0086; B = 16'h00BE; #100;
A = 16'h0086; B = 16'h00BF; #100;
A = 16'h0086; B = 16'h00C0; #100;
A = 16'h0086; B = 16'h00C1; #100;
A = 16'h0086; B = 16'h00C2; #100;
A = 16'h0086; B = 16'h00C3; #100;
A = 16'h0086; B = 16'h00C4; #100;
A = 16'h0086; B = 16'h00C5; #100;
A = 16'h0086; B = 16'h00C6; #100;
A = 16'h0086; B = 16'h00C7; #100;
A = 16'h0086; B = 16'h00C8; #100;
A = 16'h0086; B = 16'h00C9; #100;
A = 16'h0086; B = 16'h00CA; #100;
A = 16'h0086; B = 16'h00CB; #100;
A = 16'h0086; B = 16'h00CC; #100;
A = 16'h0086; B = 16'h00CD; #100;
A = 16'h0086; B = 16'h00CE; #100;
A = 16'h0086; B = 16'h00CF; #100;
A = 16'h0086; B = 16'h00D0; #100;
A = 16'h0086; B = 16'h00D1; #100;
A = 16'h0086; B = 16'h00D2; #100;
A = 16'h0086; B = 16'h00D3; #100;
A = 16'h0086; B = 16'h00D4; #100;
A = 16'h0086; B = 16'h00D5; #100;
A = 16'h0086; B = 16'h00D6; #100;
A = 16'h0086; B = 16'h00D7; #100;
A = 16'h0086; B = 16'h00D8; #100;
A = 16'h0086; B = 16'h00D9; #100;
A = 16'h0086; B = 16'h00DA; #100;
A = 16'h0086; B = 16'h00DB; #100;
A = 16'h0086; B = 16'h00DC; #100;
A = 16'h0086; B = 16'h00DD; #100;
A = 16'h0086; B = 16'h00DE; #100;
A = 16'h0086; B = 16'h00DF; #100;
A = 16'h0086; B = 16'h00E0; #100;
A = 16'h0086; B = 16'h00E1; #100;
A = 16'h0086; B = 16'h00E2; #100;
A = 16'h0086; B = 16'h00E3; #100;
A = 16'h0086; B = 16'h00E4; #100;
A = 16'h0086; B = 16'h00E5; #100;
A = 16'h0086; B = 16'h00E6; #100;
A = 16'h0086; B = 16'h00E7; #100;
A = 16'h0086; B = 16'h00E8; #100;
A = 16'h0086; B = 16'h00E9; #100;
A = 16'h0086; B = 16'h00EA; #100;
A = 16'h0086; B = 16'h00EB; #100;
A = 16'h0086; B = 16'h00EC; #100;
A = 16'h0086; B = 16'h00ED; #100;
A = 16'h0086; B = 16'h00EE; #100;
A = 16'h0086; B = 16'h00EF; #100;
A = 16'h0086; B = 16'h00F0; #100;
A = 16'h0086; B = 16'h00F1; #100;
A = 16'h0086; B = 16'h00F2; #100;
A = 16'h0086; B = 16'h00F3; #100;
A = 16'h0086; B = 16'h00F4; #100;
A = 16'h0086; B = 16'h00F5; #100;
A = 16'h0086; B = 16'h00F6; #100;
A = 16'h0086; B = 16'h00F7; #100;
A = 16'h0086; B = 16'h00F8; #100;
A = 16'h0086; B = 16'h00F9; #100;
A = 16'h0086; B = 16'h00FA; #100;
A = 16'h0086; B = 16'h00FB; #100;
A = 16'h0086; B = 16'h00FC; #100;
A = 16'h0086; B = 16'h00FD; #100;
A = 16'h0086; B = 16'h00FE; #100;
A = 16'h0086; B = 16'h00FF; #100;
A = 16'h0087; B = 16'h000; #100;
A = 16'h0087; B = 16'h001; #100;
A = 16'h0087; B = 16'h002; #100;
A = 16'h0087; B = 16'h003; #100;
A = 16'h0087; B = 16'h004; #100;
A = 16'h0087; B = 16'h005; #100;
A = 16'h0087; B = 16'h006; #100;
A = 16'h0087; B = 16'h007; #100;
A = 16'h0087; B = 16'h008; #100;
A = 16'h0087; B = 16'h009; #100;
A = 16'h0087; B = 16'h00A; #100;
A = 16'h0087; B = 16'h00B; #100;
A = 16'h0087; B = 16'h00C; #100;
A = 16'h0087; B = 16'h00D; #100;
A = 16'h0087; B = 16'h00E; #100;
A = 16'h0087; B = 16'h00F; #100;
A = 16'h0087; B = 16'h0010; #100;
A = 16'h0087; B = 16'h0011; #100;
A = 16'h0087; B = 16'h0012; #100;
A = 16'h0087; B = 16'h0013; #100;
A = 16'h0087; B = 16'h0014; #100;
A = 16'h0087; B = 16'h0015; #100;
A = 16'h0087; B = 16'h0016; #100;
A = 16'h0087; B = 16'h0017; #100;
A = 16'h0087; B = 16'h0018; #100;
A = 16'h0087; B = 16'h0019; #100;
A = 16'h0087; B = 16'h001A; #100;
A = 16'h0087; B = 16'h001B; #100;
A = 16'h0087; B = 16'h001C; #100;
A = 16'h0087; B = 16'h001D; #100;
A = 16'h0087; B = 16'h001E; #100;
A = 16'h0087; B = 16'h001F; #100;
A = 16'h0087; B = 16'h0020; #100;
A = 16'h0087; B = 16'h0021; #100;
A = 16'h0087; B = 16'h0022; #100;
A = 16'h0087; B = 16'h0023; #100;
A = 16'h0087; B = 16'h0024; #100;
A = 16'h0087; B = 16'h0025; #100;
A = 16'h0087; B = 16'h0026; #100;
A = 16'h0087; B = 16'h0027; #100;
A = 16'h0087; B = 16'h0028; #100;
A = 16'h0087; B = 16'h0029; #100;
A = 16'h0087; B = 16'h002A; #100;
A = 16'h0087; B = 16'h002B; #100;
A = 16'h0087; B = 16'h002C; #100;
A = 16'h0087; B = 16'h002D; #100;
A = 16'h0087; B = 16'h002E; #100;
A = 16'h0087; B = 16'h002F; #100;
A = 16'h0087; B = 16'h0030; #100;
A = 16'h0087; B = 16'h0031; #100;
A = 16'h0087; B = 16'h0032; #100;
A = 16'h0087; B = 16'h0033; #100;
A = 16'h0087; B = 16'h0034; #100;
A = 16'h0087; B = 16'h0035; #100;
A = 16'h0087; B = 16'h0036; #100;
A = 16'h0087; B = 16'h0037; #100;
A = 16'h0087; B = 16'h0038; #100;
A = 16'h0087; B = 16'h0039; #100;
A = 16'h0087; B = 16'h003A; #100;
A = 16'h0087; B = 16'h003B; #100;
A = 16'h0087; B = 16'h003C; #100;
A = 16'h0087; B = 16'h003D; #100;
A = 16'h0087; B = 16'h003E; #100;
A = 16'h0087; B = 16'h003F; #100;
A = 16'h0087; B = 16'h0040; #100;
A = 16'h0087; B = 16'h0041; #100;
A = 16'h0087; B = 16'h0042; #100;
A = 16'h0087; B = 16'h0043; #100;
A = 16'h0087; B = 16'h0044; #100;
A = 16'h0087; B = 16'h0045; #100;
A = 16'h0087; B = 16'h0046; #100;
A = 16'h0087; B = 16'h0047; #100;
A = 16'h0087; B = 16'h0048; #100;
A = 16'h0087; B = 16'h0049; #100;
A = 16'h0087; B = 16'h004A; #100;
A = 16'h0087; B = 16'h004B; #100;
A = 16'h0087; B = 16'h004C; #100;
A = 16'h0087; B = 16'h004D; #100;
A = 16'h0087; B = 16'h004E; #100;
A = 16'h0087; B = 16'h004F; #100;
A = 16'h0087; B = 16'h0050; #100;
A = 16'h0087; B = 16'h0051; #100;
A = 16'h0087; B = 16'h0052; #100;
A = 16'h0087; B = 16'h0053; #100;
A = 16'h0087; B = 16'h0054; #100;
A = 16'h0087; B = 16'h0055; #100;
A = 16'h0087; B = 16'h0056; #100;
A = 16'h0087; B = 16'h0057; #100;
A = 16'h0087; B = 16'h0058; #100;
A = 16'h0087; B = 16'h0059; #100;
A = 16'h0087; B = 16'h005A; #100;
A = 16'h0087; B = 16'h005B; #100;
A = 16'h0087; B = 16'h005C; #100;
A = 16'h0087; B = 16'h005D; #100;
A = 16'h0087; B = 16'h005E; #100;
A = 16'h0087; B = 16'h005F; #100;
A = 16'h0087; B = 16'h0060; #100;
A = 16'h0087; B = 16'h0061; #100;
A = 16'h0087; B = 16'h0062; #100;
A = 16'h0087; B = 16'h0063; #100;
A = 16'h0087; B = 16'h0064; #100;
A = 16'h0087; B = 16'h0065; #100;
A = 16'h0087; B = 16'h0066; #100;
A = 16'h0087; B = 16'h0067; #100;
A = 16'h0087; B = 16'h0068; #100;
A = 16'h0087; B = 16'h0069; #100;
A = 16'h0087; B = 16'h006A; #100;
A = 16'h0087; B = 16'h006B; #100;
A = 16'h0087; B = 16'h006C; #100;
A = 16'h0087; B = 16'h006D; #100;
A = 16'h0087; B = 16'h006E; #100;
A = 16'h0087; B = 16'h006F; #100;
A = 16'h0087; B = 16'h0070; #100;
A = 16'h0087; B = 16'h0071; #100;
A = 16'h0087; B = 16'h0072; #100;
A = 16'h0087; B = 16'h0073; #100;
A = 16'h0087; B = 16'h0074; #100;
A = 16'h0087; B = 16'h0075; #100;
A = 16'h0087; B = 16'h0076; #100;
A = 16'h0087; B = 16'h0077; #100;
A = 16'h0087; B = 16'h0078; #100;
A = 16'h0087; B = 16'h0079; #100;
A = 16'h0087; B = 16'h007A; #100;
A = 16'h0087; B = 16'h007B; #100;
A = 16'h0087; B = 16'h007C; #100;
A = 16'h0087; B = 16'h007D; #100;
A = 16'h0087; B = 16'h007E; #100;
A = 16'h0087; B = 16'h007F; #100;
A = 16'h0087; B = 16'h0080; #100;
A = 16'h0087; B = 16'h0081; #100;
A = 16'h0087; B = 16'h0082; #100;
A = 16'h0087; B = 16'h0083; #100;
A = 16'h0087; B = 16'h0084; #100;
A = 16'h0087; B = 16'h0085; #100;
A = 16'h0087; B = 16'h0086; #100;
A = 16'h0087; B = 16'h0087; #100;
A = 16'h0087; B = 16'h0088; #100;
A = 16'h0087; B = 16'h0089; #100;
A = 16'h0087; B = 16'h008A; #100;
A = 16'h0087; B = 16'h008B; #100;
A = 16'h0087; B = 16'h008C; #100;
A = 16'h0087; B = 16'h008D; #100;
A = 16'h0087; B = 16'h008E; #100;
A = 16'h0087; B = 16'h008F; #100;
A = 16'h0087; B = 16'h0090; #100;
A = 16'h0087; B = 16'h0091; #100;
A = 16'h0087; B = 16'h0092; #100;
A = 16'h0087; B = 16'h0093; #100;
A = 16'h0087; B = 16'h0094; #100;
A = 16'h0087; B = 16'h0095; #100;
A = 16'h0087; B = 16'h0096; #100;
A = 16'h0087; B = 16'h0097; #100;
A = 16'h0087; B = 16'h0098; #100;
A = 16'h0087; B = 16'h0099; #100;
A = 16'h0087; B = 16'h009A; #100;
A = 16'h0087; B = 16'h009B; #100;
A = 16'h0087; B = 16'h009C; #100;
A = 16'h0087; B = 16'h009D; #100;
A = 16'h0087; B = 16'h009E; #100;
A = 16'h0087; B = 16'h009F; #100;
A = 16'h0087; B = 16'h00A0; #100;
A = 16'h0087; B = 16'h00A1; #100;
A = 16'h0087; B = 16'h00A2; #100;
A = 16'h0087; B = 16'h00A3; #100;
A = 16'h0087; B = 16'h00A4; #100;
A = 16'h0087; B = 16'h00A5; #100;
A = 16'h0087; B = 16'h00A6; #100;
A = 16'h0087; B = 16'h00A7; #100;
A = 16'h0087; B = 16'h00A8; #100;
A = 16'h0087; B = 16'h00A9; #100;
A = 16'h0087; B = 16'h00AA; #100;
A = 16'h0087; B = 16'h00AB; #100;
A = 16'h0087; B = 16'h00AC; #100;
A = 16'h0087; B = 16'h00AD; #100;
A = 16'h0087; B = 16'h00AE; #100;
A = 16'h0087; B = 16'h00AF; #100;
A = 16'h0087; B = 16'h00B0; #100;
A = 16'h0087; B = 16'h00B1; #100;
A = 16'h0087; B = 16'h00B2; #100;
A = 16'h0087; B = 16'h00B3; #100;
A = 16'h0087; B = 16'h00B4; #100;
A = 16'h0087; B = 16'h00B5; #100;
A = 16'h0087; B = 16'h00B6; #100;
A = 16'h0087; B = 16'h00B7; #100;
A = 16'h0087; B = 16'h00B8; #100;
A = 16'h0087; B = 16'h00B9; #100;
A = 16'h0087; B = 16'h00BA; #100;
A = 16'h0087; B = 16'h00BB; #100;
A = 16'h0087; B = 16'h00BC; #100;
A = 16'h0087; B = 16'h00BD; #100;
A = 16'h0087; B = 16'h00BE; #100;
A = 16'h0087; B = 16'h00BF; #100;
A = 16'h0087; B = 16'h00C0; #100;
A = 16'h0087; B = 16'h00C1; #100;
A = 16'h0087; B = 16'h00C2; #100;
A = 16'h0087; B = 16'h00C3; #100;
A = 16'h0087; B = 16'h00C4; #100;
A = 16'h0087; B = 16'h00C5; #100;
A = 16'h0087; B = 16'h00C6; #100;
A = 16'h0087; B = 16'h00C7; #100;
A = 16'h0087; B = 16'h00C8; #100;
A = 16'h0087; B = 16'h00C9; #100;
A = 16'h0087; B = 16'h00CA; #100;
A = 16'h0087; B = 16'h00CB; #100;
A = 16'h0087; B = 16'h00CC; #100;
A = 16'h0087; B = 16'h00CD; #100;
A = 16'h0087; B = 16'h00CE; #100;
A = 16'h0087; B = 16'h00CF; #100;
A = 16'h0087; B = 16'h00D0; #100;
A = 16'h0087; B = 16'h00D1; #100;
A = 16'h0087; B = 16'h00D2; #100;
A = 16'h0087; B = 16'h00D3; #100;
A = 16'h0087; B = 16'h00D4; #100;
A = 16'h0087; B = 16'h00D5; #100;
A = 16'h0087; B = 16'h00D6; #100;
A = 16'h0087; B = 16'h00D7; #100;
A = 16'h0087; B = 16'h00D8; #100;
A = 16'h0087; B = 16'h00D9; #100;
A = 16'h0087; B = 16'h00DA; #100;
A = 16'h0087; B = 16'h00DB; #100;
A = 16'h0087; B = 16'h00DC; #100;
A = 16'h0087; B = 16'h00DD; #100;
A = 16'h0087; B = 16'h00DE; #100;
A = 16'h0087; B = 16'h00DF; #100;
A = 16'h0087; B = 16'h00E0; #100;
A = 16'h0087; B = 16'h00E1; #100;
A = 16'h0087; B = 16'h00E2; #100;
A = 16'h0087; B = 16'h00E3; #100;
A = 16'h0087; B = 16'h00E4; #100;
A = 16'h0087; B = 16'h00E5; #100;
A = 16'h0087; B = 16'h00E6; #100;
A = 16'h0087; B = 16'h00E7; #100;
A = 16'h0087; B = 16'h00E8; #100;
A = 16'h0087; B = 16'h00E9; #100;
A = 16'h0087; B = 16'h00EA; #100;
A = 16'h0087; B = 16'h00EB; #100;
A = 16'h0087; B = 16'h00EC; #100;
A = 16'h0087; B = 16'h00ED; #100;
A = 16'h0087; B = 16'h00EE; #100;
A = 16'h0087; B = 16'h00EF; #100;
A = 16'h0087; B = 16'h00F0; #100;
A = 16'h0087; B = 16'h00F1; #100;
A = 16'h0087; B = 16'h00F2; #100;
A = 16'h0087; B = 16'h00F3; #100;
A = 16'h0087; B = 16'h00F4; #100;
A = 16'h0087; B = 16'h00F5; #100;
A = 16'h0087; B = 16'h00F6; #100;
A = 16'h0087; B = 16'h00F7; #100;
A = 16'h0087; B = 16'h00F8; #100;
A = 16'h0087; B = 16'h00F9; #100;
A = 16'h0087; B = 16'h00FA; #100;
A = 16'h0087; B = 16'h00FB; #100;
A = 16'h0087; B = 16'h00FC; #100;
A = 16'h0087; B = 16'h00FD; #100;
A = 16'h0087; B = 16'h00FE; #100;
A = 16'h0087; B = 16'h00FF; #100;
A = 16'h0088; B = 16'h000; #100;
A = 16'h0088; B = 16'h001; #100;
A = 16'h0088; B = 16'h002; #100;
A = 16'h0088; B = 16'h003; #100;
A = 16'h0088; B = 16'h004; #100;
A = 16'h0088; B = 16'h005; #100;
A = 16'h0088; B = 16'h006; #100;
A = 16'h0088; B = 16'h007; #100;
A = 16'h0088; B = 16'h008; #100;
A = 16'h0088; B = 16'h009; #100;
A = 16'h0088; B = 16'h00A; #100;
A = 16'h0088; B = 16'h00B; #100;
A = 16'h0088; B = 16'h00C; #100;
A = 16'h0088; B = 16'h00D; #100;
A = 16'h0088; B = 16'h00E; #100;
A = 16'h0088; B = 16'h00F; #100;
A = 16'h0088; B = 16'h0010; #100;
A = 16'h0088; B = 16'h0011; #100;
A = 16'h0088; B = 16'h0012; #100;
A = 16'h0088; B = 16'h0013; #100;
A = 16'h0088; B = 16'h0014; #100;
A = 16'h0088; B = 16'h0015; #100;
A = 16'h0088; B = 16'h0016; #100;
A = 16'h0088; B = 16'h0017; #100;
A = 16'h0088; B = 16'h0018; #100;
A = 16'h0088; B = 16'h0019; #100;
A = 16'h0088; B = 16'h001A; #100;
A = 16'h0088; B = 16'h001B; #100;
A = 16'h0088; B = 16'h001C; #100;
A = 16'h0088; B = 16'h001D; #100;
A = 16'h0088; B = 16'h001E; #100;
A = 16'h0088; B = 16'h001F; #100;
A = 16'h0088; B = 16'h0020; #100;
A = 16'h0088; B = 16'h0021; #100;
A = 16'h0088; B = 16'h0022; #100;
A = 16'h0088; B = 16'h0023; #100;
A = 16'h0088; B = 16'h0024; #100;
A = 16'h0088; B = 16'h0025; #100;
A = 16'h0088; B = 16'h0026; #100;
A = 16'h0088; B = 16'h0027; #100;
A = 16'h0088; B = 16'h0028; #100;
A = 16'h0088; B = 16'h0029; #100;
A = 16'h0088; B = 16'h002A; #100;
A = 16'h0088; B = 16'h002B; #100;
A = 16'h0088; B = 16'h002C; #100;
A = 16'h0088; B = 16'h002D; #100;
A = 16'h0088; B = 16'h002E; #100;
A = 16'h0088; B = 16'h002F; #100;
A = 16'h0088; B = 16'h0030; #100;
A = 16'h0088; B = 16'h0031; #100;
A = 16'h0088; B = 16'h0032; #100;
A = 16'h0088; B = 16'h0033; #100;
A = 16'h0088; B = 16'h0034; #100;
A = 16'h0088; B = 16'h0035; #100;
A = 16'h0088; B = 16'h0036; #100;
A = 16'h0088; B = 16'h0037; #100;
A = 16'h0088; B = 16'h0038; #100;
A = 16'h0088; B = 16'h0039; #100;
A = 16'h0088; B = 16'h003A; #100;
A = 16'h0088; B = 16'h003B; #100;
A = 16'h0088; B = 16'h003C; #100;
A = 16'h0088; B = 16'h003D; #100;
A = 16'h0088; B = 16'h003E; #100;
A = 16'h0088; B = 16'h003F; #100;
A = 16'h0088; B = 16'h0040; #100;
A = 16'h0088; B = 16'h0041; #100;
A = 16'h0088; B = 16'h0042; #100;
A = 16'h0088; B = 16'h0043; #100;
A = 16'h0088; B = 16'h0044; #100;
A = 16'h0088; B = 16'h0045; #100;
A = 16'h0088; B = 16'h0046; #100;
A = 16'h0088; B = 16'h0047; #100;
A = 16'h0088; B = 16'h0048; #100;
A = 16'h0088; B = 16'h0049; #100;
A = 16'h0088; B = 16'h004A; #100;
A = 16'h0088; B = 16'h004B; #100;
A = 16'h0088; B = 16'h004C; #100;
A = 16'h0088; B = 16'h004D; #100;
A = 16'h0088; B = 16'h004E; #100;
A = 16'h0088; B = 16'h004F; #100;
A = 16'h0088; B = 16'h0050; #100;
A = 16'h0088; B = 16'h0051; #100;
A = 16'h0088; B = 16'h0052; #100;
A = 16'h0088; B = 16'h0053; #100;
A = 16'h0088; B = 16'h0054; #100;
A = 16'h0088; B = 16'h0055; #100;
A = 16'h0088; B = 16'h0056; #100;
A = 16'h0088; B = 16'h0057; #100;
A = 16'h0088; B = 16'h0058; #100;
A = 16'h0088; B = 16'h0059; #100;
A = 16'h0088; B = 16'h005A; #100;
A = 16'h0088; B = 16'h005B; #100;
A = 16'h0088; B = 16'h005C; #100;
A = 16'h0088; B = 16'h005D; #100;
A = 16'h0088; B = 16'h005E; #100;
A = 16'h0088; B = 16'h005F; #100;
A = 16'h0088; B = 16'h0060; #100;
A = 16'h0088; B = 16'h0061; #100;
A = 16'h0088; B = 16'h0062; #100;
A = 16'h0088; B = 16'h0063; #100;
A = 16'h0088; B = 16'h0064; #100;
A = 16'h0088; B = 16'h0065; #100;
A = 16'h0088; B = 16'h0066; #100;
A = 16'h0088; B = 16'h0067; #100;
A = 16'h0088; B = 16'h0068; #100;
A = 16'h0088; B = 16'h0069; #100;
A = 16'h0088; B = 16'h006A; #100;
A = 16'h0088; B = 16'h006B; #100;
A = 16'h0088; B = 16'h006C; #100;
A = 16'h0088; B = 16'h006D; #100;
A = 16'h0088; B = 16'h006E; #100;
A = 16'h0088; B = 16'h006F; #100;
A = 16'h0088; B = 16'h0070; #100;
A = 16'h0088; B = 16'h0071; #100;
A = 16'h0088; B = 16'h0072; #100;
A = 16'h0088; B = 16'h0073; #100;
A = 16'h0088; B = 16'h0074; #100;
A = 16'h0088; B = 16'h0075; #100;
A = 16'h0088; B = 16'h0076; #100;
A = 16'h0088; B = 16'h0077; #100;
A = 16'h0088; B = 16'h0078; #100;
A = 16'h0088; B = 16'h0079; #100;
A = 16'h0088; B = 16'h007A; #100;
A = 16'h0088; B = 16'h007B; #100;
A = 16'h0088; B = 16'h007C; #100;
A = 16'h0088; B = 16'h007D; #100;
A = 16'h0088; B = 16'h007E; #100;
A = 16'h0088; B = 16'h007F; #100;
A = 16'h0088; B = 16'h0080; #100;
A = 16'h0088; B = 16'h0081; #100;
A = 16'h0088; B = 16'h0082; #100;
A = 16'h0088; B = 16'h0083; #100;
A = 16'h0088; B = 16'h0084; #100;
A = 16'h0088; B = 16'h0085; #100;
A = 16'h0088; B = 16'h0086; #100;
A = 16'h0088; B = 16'h0087; #100;
A = 16'h0088; B = 16'h0088; #100;
A = 16'h0088; B = 16'h0089; #100;
A = 16'h0088; B = 16'h008A; #100;
A = 16'h0088; B = 16'h008B; #100;
A = 16'h0088; B = 16'h008C; #100;
A = 16'h0088; B = 16'h008D; #100;
A = 16'h0088; B = 16'h008E; #100;
A = 16'h0088; B = 16'h008F; #100;
A = 16'h0088; B = 16'h0090; #100;
A = 16'h0088; B = 16'h0091; #100;
A = 16'h0088; B = 16'h0092; #100;
A = 16'h0088; B = 16'h0093; #100;
A = 16'h0088; B = 16'h0094; #100;
A = 16'h0088; B = 16'h0095; #100;
A = 16'h0088; B = 16'h0096; #100;
A = 16'h0088; B = 16'h0097; #100;
A = 16'h0088; B = 16'h0098; #100;
A = 16'h0088; B = 16'h0099; #100;
A = 16'h0088; B = 16'h009A; #100;
A = 16'h0088; B = 16'h009B; #100;
A = 16'h0088; B = 16'h009C; #100;
A = 16'h0088; B = 16'h009D; #100;
A = 16'h0088; B = 16'h009E; #100;
A = 16'h0088; B = 16'h009F; #100;
A = 16'h0088; B = 16'h00A0; #100;
A = 16'h0088; B = 16'h00A1; #100;
A = 16'h0088; B = 16'h00A2; #100;
A = 16'h0088; B = 16'h00A3; #100;
A = 16'h0088; B = 16'h00A4; #100;
A = 16'h0088; B = 16'h00A5; #100;
A = 16'h0088; B = 16'h00A6; #100;
A = 16'h0088; B = 16'h00A7; #100;
A = 16'h0088; B = 16'h00A8; #100;
A = 16'h0088; B = 16'h00A9; #100;
A = 16'h0088; B = 16'h00AA; #100;
A = 16'h0088; B = 16'h00AB; #100;
A = 16'h0088; B = 16'h00AC; #100;
A = 16'h0088; B = 16'h00AD; #100;
A = 16'h0088; B = 16'h00AE; #100;
A = 16'h0088; B = 16'h00AF; #100;
A = 16'h0088; B = 16'h00B0; #100;
A = 16'h0088; B = 16'h00B1; #100;
A = 16'h0088; B = 16'h00B2; #100;
A = 16'h0088; B = 16'h00B3; #100;
A = 16'h0088; B = 16'h00B4; #100;
A = 16'h0088; B = 16'h00B5; #100;
A = 16'h0088; B = 16'h00B6; #100;
A = 16'h0088; B = 16'h00B7; #100;
A = 16'h0088; B = 16'h00B8; #100;
A = 16'h0088; B = 16'h00B9; #100;
A = 16'h0088; B = 16'h00BA; #100;
A = 16'h0088; B = 16'h00BB; #100;
A = 16'h0088; B = 16'h00BC; #100;
A = 16'h0088; B = 16'h00BD; #100;
A = 16'h0088; B = 16'h00BE; #100;
A = 16'h0088; B = 16'h00BF; #100;
A = 16'h0088; B = 16'h00C0; #100;
A = 16'h0088; B = 16'h00C1; #100;
A = 16'h0088; B = 16'h00C2; #100;
A = 16'h0088; B = 16'h00C3; #100;
A = 16'h0088; B = 16'h00C4; #100;
A = 16'h0088; B = 16'h00C5; #100;
A = 16'h0088; B = 16'h00C6; #100;
A = 16'h0088; B = 16'h00C7; #100;
A = 16'h0088; B = 16'h00C8; #100;
A = 16'h0088; B = 16'h00C9; #100;
A = 16'h0088; B = 16'h00CA; #100;
A = 16'h0088; B = 16'h00CB; #100;
A = 16'h0088; B = 16'h00CC; #100;
A = 16'h0088; B = 16'h00CD; #100;
A = 16'h0088; B = 16'h00CE; #100;
A = 16'h0088; B = 16'h00CF; #100;
A = 16'h0088; B = 16'h00D0; #100;
A = 16'h0088; B = 16'h00D1; #100;
A = 16'h0088; B = 16'h00D2; #100;
A = 16'h0088; B = 16'h00D3; #100;
A = 16'h0088; B = 16'h00D4; #100;
A = 16'h0088; B = 16'h00D5; #100;
A = 16'h0088; B = 16'h00D6; #100;
A = 16'h0088; B = 16'h00D7; #100;
A = 16'h0088; B = 16'h00D8; #100;
A = 16'h0088; B = 16'h00D9; #100;
A = 16'h0088; B = 16'h00DA; #100;
A = 16'h0088; B = 16'h00DB; #100;
A = 16'h0088; B = 16'h00DC; #100;
A = 16'h0088; B = 16'h00DD; #100;
A = 16'h0088; B = 16'h00DE; #100;
A = 16'h0088; B = 16'h00DF; #100;
A = 16'h0088; B = 16'h00E0; #100;
A = 16'h0088; B = 16'h00E1; #100;
A = 16'h0088; B = 16'h00E2; #100;
A = 16'h0088; B = 16'h00E3; #100;
A = 16'h0088; B = 16'h00E4; #100;
A = 16'h0088; B = 16'h00E5; #100;
A = 16'h0088; B = 16'h00E6; #100;
A = 16'h0088; B = 16'h00E7; #100;
A = 16'h0088; B = 16'h00E8; #100;
A = 16'h0088; B = 16'h00E9; #100;
A = 16'h0088; B = 16'h00EA; #100;
A = 16'h0088; B = 16'h00EB; #100;
A = 16'h0088; B = 16'h00EC; #100;
A = 16'h0088; B = 16'h00ED; #100;
A = 16'h0088; B = 16'h00EE; #100;
A = 16'h0088; B = 16'h00EF; #100;
A = 16'h0088; B = 16'h00F0; #100;
A = 16'h0088; B = 16'h00F1; #100;
A = 16'h0088; B = 16'h00F2; #100;
A = 16'h0088; B = 16'h00F3; #100;
A = 16'h0088; B = 16'h00F4; #100;
A = 16'h0088; B = 16'h00F5; #100;
A = 16'h0088; B = 16'h00F6; #100;
A = 16'h0088; B = 16'h00F7; #100;
A = 16'h0088; B = 16'h00F8; #100;
A = 16'h0088; B = 16'h00F9; #100;
A = 16'h0088; B = 16'h00FA; #100;
A = 16'h0088; B = 16'h00FB; #100;
A = 16'h0088; B = 16'h00FC; #100;
A = 16'h0088; B = 16'h00FD; #100;
A = 16'h0088; B = 16'h00FE; #100;
A = 16'h0088; B = 16'h00FF; #100;
A = 16'h0089; B = 16'h000; #100;
A = 16'h0089; B = 16'h001; #100;
A = 16'h0089; B = 16'h002; #100;
A = 16'h0089; B = 16'h003; #100;
A = 16'h0089; B = 16'h004; #100;
A = 16'h0089; B = 16'h005; #100;
A = 16'h0089; B = 16'h006; #100;
A = 16'h0089; B = 16'h007; #100;
A = 16'h0089; B = 16'h008; #100;
A = 16'h0089; B = 16'h009; #100;
A = 16'h0089; B = 16'h00A; #100;
A = 16'h0089; B = 16'h00B; #100;
A = 16'h0089; B = 16'h00C; #100;
A = 16'h0089; B = 16'h00D; #100;
A = 16'h0089; B = 16'h00E; #100;
A = 16'h0089; B = 16'h00F; #100;
A = 16'h0089; B = 16'h0010; #100;
A = 16'h0089; B = 16'h0011; #100;
A = 16'h0089; B = 16'h0012; #100;
A = 16'h0089; B = 16'h0013; #100;
A = 16'h0089; B = 16'h0014; #100;
A = 16'h0089; B = 16'h0015; #100;
A = 16'h0089; B = 16'h0016; #100;
A = 16'h0089; B = 16'h0017; #100;
A = 16'h0089; B = 16'h0018; #100;
A = 16'h0089; B = 16'h0019; #100;
A = 16'h0089; B = 16'h001A; #100;
A = 16'h0089; B = 16'h001B; #100;
A = 16'h0089; B = 16'h001C; #100;
A = 16'h0089; B = 16'h001D; #100;
A = 16'h0089; B = 16'h001E; #100;
A = 16'h0089; B = 16'h001F; #100;
A = 16'h0089; B = 16'h0020; #100;
A = 16'h0089; B = 16'h0021; #100;
A = 16'h0089; B = 16'h0022; #100;
A = 16'h0089; B = 16'h0023; #100;
A = 16'h0089; B = 16'h0024; #100;
A = 16'h0089; B = 16'h0025; #100;
A = 16'h0089; B = 16'h0026; #100;
A = 16'h0089; B = 16'h0027; #100;
A = 16'h0089; B = 16'h0028; #100;
A = 16'h0089; B = 16'h0029; #100;
A = 16'h0089; B = 16'h002A; #100;
A = 16'h0089; B = 16'h002B; #100;
A = 16'h0089; B = 16'h002C; #100;
A = 16'h0089; B = 16'h002D; #100;
A = 16'h0089; B = 16'h002E; #100;
A = 16'h0089; B = 16'h002F; #100;
A = 16'h0089; B = 16'h0030; #100;
A = 16'h0089; B = 16'h0031; #100;
A = 16'h0089; B = 16'h0032; #100;
A = 16'h0089; B = 16'h0033; #100;
A = 16'h0089; B = 16'h0034; #100;
A = 16'h0089; B = 16'h0035; #100;
A = 16'h0089; B = 16'h0036; #100;
A = 16'h0089; B = 16'h0037; #100;
A = 16'h0089; B = 16'h0038; #100;
A = 16'h0089; B = 16'h0039; #100;
A = 16'h0089; B = 16'h003A; #100;
A = 16'h0089; B = 16'h003B; #100;
A = 16'h0089; B = 16'h003C; #100;
A = 16'h0089; B = 16'h003D; #100;
A = 16'h0089; B = 16'h003E; #100;
A = 16'h0089; B = 16'h003F; #100;
A = 16'h0089; B = 16'h0040; #100;
A = 16'h0089; B = 16'h0041; #100;
A = 16'h0089; B = 16'h0042; #100;
A = 16'h0089; B = 16'h0043; #100;
A = 16'h0089; B = 16'h0044; #100;
A = 16'h0089; B = 16'h0045; #100;
A = 16'h0089; B = 16'h0046; #100;
A = 16'h0089; B = 16'h0047; #100;
A = 16'h0089; B = 16'h0048; #100;
A = 16'h0089; B = 16'h0049; #100;
A = 16'h0089; B = 16'h004A; #100;
A = 16'h0089; B = 16'h004B; #100;
A = 16'h0089; B = 16'h004C; #100;
A = 16'h0089; B = 16'h004D; #100;
A = 16'h0089; B = 16'h004E; #100;
A = 16'h0089; B = 16'h004F; #100;
A = 16'h0089; B = 16'h0050; #100;
A = 16'h0089; B = 16'h0051; #100;
A = 16'h0089; B = 16'h0052; #100;
A = 16'h0089; B = 16'h0053; #100;
A = 16'h0089; B = 16'h0054; #100;
A = 16'h0089; B = 16'h0055; #100;
A = 16'h0089; B = 16'h0056; #100;
A = 16'h0089; B = 16'h0057; #100;
A = 16'h0089; B = 16'h0058; #100;
A = 16'h0089; B = 16'h0059; #100;
A = 16'h0089; B = 16'h005A; #100;
A = 16'h0089; B = 16'h005B; #100;
A = 16'h0089; B = 16'h005C; #100;
A = 16'h0089; B = 16'h005D; #100;
A = 16'h0089; B = 16'h005E; #100;
A = 16'h0089; B = 16'h005F; #100;
A = 16'h0089; B = 16'h0060; #100;
A = 16'h0089; B = 16'h0061; #100;
A = 16'h0089; B = 16'h0062; #100;
A = 16'h0089; B = 16'h0063; #100;
A = 16'h0089; B = 16'h0064; #100;
A = 16'h0089; B = 16'h0065; #100;
A = 16'h0089; B = 16'h0066; #100;
A = 16'h0089; B = 16'h0067; #100;
A = 16'h0089; B = 16'h0068; #100;
A = 16'h0089; B = 16'h0069; #100;
A = 16'h0089; B = 16'h006A; #100;
A = 16'h0089; B = 16'h006B; #100;
A = 16'h0089; B = 16'h006C; #100;
A = 16'h0089; B = 16'h006D; #100;
A = 16'h0089; B = 16'h006E; #100;
A = 16'h0089; B = 16'h006F; #100;
A = 16'h0089; B = 16'h0070; #100;
A = 16'h0089; B = 16'h0071; #100;
A = 16'h0089; B = 16'h0072; #100;
A = 16'h0089; B = 16'h0073; #100;
A = 16'h0089; B = 16'h0074; #100;
A = 16'h0089; B = 16'h0075; #100;
A = 16'h0089; B = 16'h0076; #100;
A = 16'h0089; B = 16'h0077; #100;
A = 16'h0089; B = 16'h0078; #100;
A = 16'h0089; B = 16'h0079; #100;
A = 16'h0089; B = 16'h007A; #100;
A = 16'h0089; B = 16'h007B; #100;
A = 16'h0089; B = 16'h007C; #100;
A = 16'h0089; B = 16'h007D; #100;
A = 16'h0089; B = 16'h007E; #100;
A = 16'h0089; B = 16'h007F; #100;
A = 16'h0089; B = 16'h0080; #100;
A = 16'h0089; B = 16'h0081; #100;
A = 16'h0089; B = 16'h0082; #100;
A = 16'h0089; B = 16'h0083; #100;
A = 16'h0089; B = 16'h0084; #100;
A = 16'h0089; B = 16'h0085; #100;
A = 16'h0089; B = 16'h0086; #100;
A = 16'h0089; B = 16'h0087; #100;
A = 16'h0089; B = 16'h0088; #100;
A = 16'h0089; B = 16'h0089; #100;
A = 16'h0089; B = 16'h008A; #100;
A = 16'h0089; B = 16'h008B; #100;
A = 16'h0089; B = 16'h008C; #100;
A = 16'h0089; B = 16'h008D; #100;
A = 16'h0089; B = 16'h008E; #100;
A = 16'h0089; B = 16'h008F; #100;
A = 16'h0089; B = 16'h0090; #100;
A = 16'h0089; B = 16'h0091; #100;
A = 16'h0089; B = 16'h0092; #100;
A = 16'h0089; B = 16'h0093; #100;
A = 16'h0089; B = 16'h0094; #100;
A = 16'h0089; B = 16'h0095; #100;
A = 16'h0089; B = 16'h0096; #100;
A = 16'h0089; B = 16'h0097; #100;
A = 16'h0089; B = 16'h0098; #100;
A = 16'h0089; B = 16'h0099; #100;
A = 16'h0089; B = 16'h009A; #100;
A = 16'h0089; B = 16'h009B; #100;
A = 16'h0089; B = 16'h009C; #100;
A = 16'h0089; B = 16'h009D; #100;
A = 16'h0089; B = 16'h009E; #100;
A = 16'h0089; B = 16'h009F; #100;
A = 16'h0089; B = 16'h00A0; #100;
A = 16'h0089; B = 16'h00A1; #100;
A = 16'h0089; B = 16'h00A2; #100;
A = 16'h0089; B = 16'h00A3; #100;
A = 16'h0089; B = 16'h00A4; #100;
A = 16'h0089; B = 16'h00A5; #100;
A = 16'h0089; B = 16'h00A6; #100;
A = 16'h0089; B = 16'h00A7; #100;
A = 16'h0089; B = 16'h00A8; #100;
A = 16'h0089; B = 16'h00A9; #100;
A = 16'h0089; B = 16'h00AA; #100;
A = 16'h0089; B = 16'h00AB; #100;
A = 16'h0089; B = 16'h00AC; #100;
A = 16'h0089; B = 16'h00AD; #100;
A = 16'h0089; B = 16'h00AE; #100;
A = 16'h0089; B = 16'h00AF; #100;
A = 16'h0089; B = 16'h00B0; #100;
A = 16'h0089; B = 16'h00B1; #100;
A = 16'h0089; B = 16'h00B2; #100;
A = 16'h0089; B = 16'h00B3; #100;
A = 16'h0089; B = 16'h00B4; #100;
A = 16'h0089; B = 16'h00B5; #100;
A = 16'h0089; B = 16'h00B6; #100;
A = 16'h0089; B = 16'h00B7; #100;
A = 16'h0089; B = 16'h00B8; #100;
A = 16'h0089; B = 16'h00B9; #100;
A = 16'h0089; B = 16'h00BA; #100;
A = 16'h0089; B = 16'h00BB; #100;
A = 16'h0089; B = 16'h00BC; #100;
A = 16'h0089; B = 16'h00BD; #100;
A = 16'h0089; B = 16'h00BE; #100;
A = 16'h0089; B = 16'h00BF; #100;
A = 16'h0089; B = 16'h00C0; #100;
A = 16'h0089; B = 16'h00C1; #100;
A = 16'h0089; B = 16'h00C2; #100;
A = 16'h0089; B = 16'h00C3; #100;
A = 16'h0089; B = 16'h00C4; #100;
A = 16'h0089; B = 16'h00C5; #100;
A = 16'h0089; B = 16'h00C6; #100;
A = 16'h0089; B = 16'h00C7; #100;
A = 16'h0089; B = 16'h00C8; #100;
A = 16'h0089; B = 16'h00C9; #100;
A = 16'h0089; B = 16'h00CA; #100;
A = 16'h0089; B = 16'h00CB; #100;
A = 16'h0089; B = 16'h00CC; #100;
A = 16'h0089; B = 16'h00CD; #100;
A = 16'h0089; B = 16'h00CE; #100;
A = 16'h0089; B = 16'h00CF; #100;
A = 16'h0089; B = 16'h00D0; #100;
A = 16'h0089; B = 16'h00D1; #100;
A = 16'h0089; B = 16'h00D2; #100;
A = 16'h0089; B = 16'h00D3; #100;
A = 16'h0089; B = 16'h00D4; #100;
A = 16'h0089; B = 16'h00D5; #100;
A = 16'h0089; B = 16'h00D6; #100;
A = 16'h0089; B = 16'h00D7; #100;
A = 16'h0089; B = 16'h00D8; #100;
A = 16'h0089; B = 16'h00D9; #100;
A = 16'h0089; B = 16'h00DA; #100;
A = 16'h0089; B = 16'h00DB; #100;
A = 16'h0089; B = 16'h00DC; #100;
A = 16'h0089; B = 16'h00DD; #100;
A = 16'h0089; B = 16'h00DE; #100;
A = 16'h0089; B = 16'h00DF; #100;
A = 16'h0089; B = 16'h00E0; #100;
A = 16'h0089; B = 16'h00E1; #100;
A = 16'h0089; B = 16'h00E2; #100;
A = 16'h0089; B = 16'h00E3; #100;
A = 16'h0089; B = 16'h00E4; #100;
A = 16'h0089; B = 16'h00E5; #100;
A = 16'h0089; B = 16'h00E6; #100;
A = 16'h0089; B = 16'h00E7; #100;
A = 16'h0089; B = 16'h00E8; #100;
A = 16'h0089; B = 16'h00E9; #100;
A = 16'h0089; B = 16'h00EA; #100;
A = 16'h0089; B = 16'h00EB; #100;
A = 16'h0089; B = 16'h00EC; #100;
A = 16'h0089; B = 16'h00ED; #100;
A = 16'h0089; B = 16'h00EE; #100;
A = 16'h0089; B = 16'h00EF; #100;
A = 16'h0089; B = 16'h00F0; #100;
A = 16'h0089; B = 16'h00F1; #100;
A = 16'h0089; B = 16'h00F2; #100;
A = 16'h0089; B = 16'h00F3; #100;
A = 16'h0089; B = 16'h00F4; #100;
A = 16'h0089; B = 16'h00F5; #100;
A = 16'h0089; B = 16'h00F6; #100;
A = 16'h0089; B = 16'h00F7; #100;
A = 16'h0089; B = 16'h00F8; #100;
A = 16'h0089; B = 16'h00F9; #100;
A = 16'h0089; B = 16'h00FA; #100;
A = 16'h0089; B = 16'h00FB; #100;
A = 16'h0089; B = 16'h00FC; #100;
A = 16'h0089; B = 16'h00FD; #100;
A = 16'h0089; B = 16'h00FE; #100;
A = 16'h0089; B = 16'h00FF; #100;
A = 16'h008A; B = 16'h000; #100;
A = 16'h008A; B = 16'h001; #100;
A = 16'h008A; B = 16'h002; #100;
A = 16'h008A; B = 16'h003; #100;
A = 16'h008A; B = 16'h004; #100;
A = 16'h008A; B = 16'h005; #100;
A = 16'h008A; B = 16'h006; #100;
A = 16'h008A; B = 16'h007; #100;
A = 16'h008A; B = 16'h008; #100;
A = 16'h008A; B = 16'h009; #100;
A = 16'h008A; B = 16'h00A; #100;
A = 16'h008A; B = 16'h00B; #100;
A = 16'h008A; B = 16'h00C; #100;
A = 16'h008A; B = 16'h00D; #100;
A = 16'h008A; B = 16'h00E; #100;
A = 16'h008A; B = 16'h00F; #100;
A = 16'h008A; B = 16'h0010; #100;
A = 16'h008A; B = 16'h0011; #100;
A = 16'h008A; B = 16'h0012; #100;
A = 16'h008A; B = 16'h0013; #100;
A = 16'h008A; B = 16'h0014; #100;
A = 16'h008A; B = 16'h0015; #100;
A = 16'h008A; B = 16'h0016; #100;
A = 16'h008A; B = 16'h0017; #100;
A = 16'h008A; B = 16'h0018; #100;
A = 16'h008A; B = 16'h0019; #100;
A = 16'h008A; B = 16'h001A; #100;
A = 16'h008A; B = 16'h001B; #100;
A = 16'h008A; B = 16'h001C; #100;
A = 16'h008A; B = 16'h001D; #100;
A = 16'h008A; B = 16'h001E; #100;
A = 16'h008A; B = 16'h001F; #100;
A = 16'h008A; B = 16'h0020; #100;
A = 16'h008A; B = 16'h0021; #100;
A = 16'h008A; B = 16'h0022; #100;
A = 16'h008A; B = 16'h0023; #100;
A = 16'h008A; B = 16'h0024; #100;
A = 16'h008A; B = 16'h0025; #100;
A = 16'h008A; B = 16'h0026; #100;
A = 16'h008A; B = 16'h0027; #100;
A = 16'h008A; B = 16'h0028; #100;
A = 16'h008A; B = 16'h0029; #100;
A = 16'h008A; B = 16'h002A; #100;
A = 16'h008A; B = 16'h002B; #100;
A = 16'h008A; B = 16'h002C; #100;
A = 16'h008A; B = 16'h002D; #100;
A = 16'h008A; B = 16'h002E; #100;
A = 16'h008A; B = 16'h002F; #100;
A = 16'h008A; B = 16'h0030; #100;
A = 16'h008A; B = 16'h0031; #100;
A = 16'h008A; B = 16'h0032; #100;
A = 16'h008A; B = 16'h0033; #100;
A = 16'h008A; B = 16'h0034; #100;
A = 16'h008A; B = 16'h0035; #100;
A = 16'h008A; B = 16'h0036; #100;
A = 16'h008A; B = 16'h0037; #100;
A = 16'h008A; B = 16'h0038; #100;
A = 16'h008A; B = 16'h0039; #100;
A = 16'h008A; B = 16'h003A; #100;
A = 16'h008A; B = 16'h003B; #100;
A = 16'h008A; B = 16'h003C; #100;
A = 16'h008A; B = 16'h003D; #100;
A = 16'h008A; B = 16'h003E; #100;
A = 16'h008A; B = 16'h003F; #100;
A = 16'h008A; B = 16'h0040; #100;
A = 16'h008A; B = 16'h0041; #100;
A = 16'h008A; B = 16'h0042; #100;
A = 16'h008A; B = 16'h0043; #100;
A = 16'h008A; B = 16'h0044; #100;
A = 16'h008A; B = 16'h0045; #100;
A = 16'h008A; B = 16'h0046; #100;
A = 16'h008A; B = 16'h0047; #100;
A = 16'h008A; B = 16'h0048; #100;
A = 16'h008A; B = 16'h0049; #100;
A = 16'h008A; B = 16'h004A; #100;
A = 16'h008A; B = 16'h004B; #100;
A = 16'h008A; B = 16'h004C; #100;
A = 16'h008A; B = 16'h004D; #100;
A = 16'h008A; B = 16'h004E; #100;
A = 16'h008A; B = 16'h004F; #100;
A = 16'h008A; B = 16'h0050; #100;
A = 16'h008A; B = 16'h0051; #100;
A = 16'h008A; B = 16'h0052; #100;
A = 16'h008A; B = 16'h0053; #100;
A = 16'h008A; B = 16'h0054; #100;
A = 16'h008A; B = 16'h0055; #100;
A = 16'h008A; B = 16'h0056; #100;
A = 16'h008A; B = 16'h0057; #100;
A = 16'h008A; B = 16'h0058; #100;
A = 16'h008A; B = 16'h0059; #100;
A = 16'h008A; B = 16'h005A; #100;
A = 16'h008A; B = 16'h005B; #100;
A = 16'h008A; B = 16'h005C; #100;
A = 16'h008A; B = 16'h005D; #100;
A = 16'h008A; B = 16'h005E; #100;
A = 16'h008A; B = 16'h005F; #100;
A = 16'h008A; B = 16'h0060; #100;
A = 16'h008A; B = 16'h0061; #100;
A = 16'h008A; B = 16'h0062; #100;
A = 16'h008A; B = 16'h0063; #100;
A = 16'h008A; B = 16'h0064; #100;
A = 16'h008A; B = 16'h0065; #100;
A = 16'h008A; B = 16'h0066; #100;
A = 16'h008A; B = 16'h0067; #100;
A = 16'h008A; B = 16'h0068; #100;
A = 16'h008A; B = 16'h0069; #100;
A = 16'h008A; B = 16'h006A; #100;
A = 16'h008A; B = 16'h006B; #100;
A = 16'h008A; B = 16'h006C; #100;
A = 16'h008A; B = 16'h006D; #100;
A = 16'h008A; B = 16'h006E; #100;
A = 16'h008A; B = 16'h006F; #100;
A = 16'h008A; B = 16'h0070; #100;
A = 16'h008A; B = 16'h0071; #100;
A = 16'h008A; B = 16'h0072; #100;
A = 16'h008A; B = 16'h0073; #100;
A = 16'h008A; B = 16'h0074; #100;
A = 16'h008A; B = 16'h0075; #100;
A = 16'h008A; B = 16'h0076; #100;
A = 16'h008A; B = 16'h0077; #100;
A = 16'h008A; B = 16'h0078; #100;
A = 16'h008A; B = 16'h0079; #100;
A = 16'h008A; B = 16'h007A; #100;
A = 16'h008A; B = 16'h007B; #100;
A = 16'h008A; B = 16'h007C; #100;
A = 16'h008A; B = 16'h007D; #100;
A = 16'h008A; B = 16'h007E; #100;
A = 16'h008A; B = 16'h007F; #100;
A = 16'h008A; B = 16'h0080; #100;
A = 16'h008A; B = 16'h0081; #100;
A = 16'h008A; B = 16'h0082; #100;
A = 16'h008A; B = 16'h0083; #100;
A = 16'h008A; B = 16'h0084; #100;
A = 16'h008A; B = 16'h0085; #100;
A = 16'h008A; B = 16'h0086; #100;
A = 16'h008A; B = 16'h0087; #100;
A = 16'h008A; B = 16'h0088; #100;
A = 16'h008A; B = 16'h0089; #100;
A = 16'h008A; B = 16'h008A; #100;
A = 16'h008A; B = 16'h008B; #100;
A = 16'h008A; B = 16'h008C; #100;
A = 16'h008A; B = 16'h008D; #100;
A = 16'h008A; B = 16'h008E; #100;
A = 16'h008A; B = 16'h008F; #100;
A = 16'h008A; B = 16'h0090; #100;
A = 16'h008A; B = 16'h0091; #100;
A = 16'h008A; B = 16'h0092; #100;
A = 16'h008A; B = 16'h0093; #100;
A = 16'h008A; B = 16'h0094; #100;
A = 16'h008A; B = 16'h0095; #100;
A = 16'h008A; B = 16'h0096; #100;
A = 16'h008A; B = 16'h0097; #100;
A = 16'h008A; B = 16'h0098; #100;
A = 16'h008A; B = 16'h0099; #100;
A = 16'h008A; B = 16'h009A; #100;
A = 16'h008A; B = 16'h009B; #100;
A = 16'h008A; B = 16'h009C; #100;
A = 16'h008A; B = 16'h009D; #100;
A = 16'h008A; B = 16'h009E; #100;
A = 16'h008A; B = 16'h009F; #100;
A = 16'h008A; B = 16'h00A0; #100;
A = 16'h008A; B = 16'h00A1; #100;
A = 16'h008A; B = 16'h00A2; #100;
A = 16'h008A; B = 16'h00A3; #100;
A = 16'h008A; B = 16'h00A4; #100;
A = 16'h008A; B = 16'h00A5; #100;
A = 16'h008A; B = 16'h00A6; #100;
A = 16'h008A; B = 16'h00A7; #100;
A = 16'h008A; B = 16'h00A8; #100;
A = 16'h008A; B = 16'h00A9; #100;
A = 16'h008A; B = 16'h00AA; #100;
A = 16'h008A; B = 16'h00AB; #100;
A = 16'h008A; B = 16'h00AC; #100;
A = 16'h008A; B = 16'h00AD; #100;
A = 16'h008A; B = 16'h00AE; #100;
A = 16'h008A; B = 16'h00AF; #100;
A = 16'h008A; B = 16'h00B0; #100;
A = 16'h008A; B = 16'h00B1; #100;
A = 16'h008A; B = 16'h00B2; #100;
A = 16'h008A; B = 16'h00B3; #100;
A = 16'h008A; B = 16'h00B4; #100;
A = 16'h008A; B = 16'h00B5; #100;
A = 16'h008A; B = 16'h00B6; #100;
A = 16'h008A; B = 16'h00B7; #100;
A = 16'h008A; B = 16'h00B8; #100;
A = 16'h008A; B = 16'h00B9; #100;
A = 16'h008A; B = 16'h00BA; #100;
A = 16'h008A; B = 16'h00BB; #100;
A = 16'h008A; B = 16'h00BC; #100;
A = 16'h008A; B = 16'h00BD; #100;
A = 16'h008A; B = 16'h00BE; #100;
A = 16'h008A; B = 16'h00BF; #100;
A = 16'h008A; B = 16'h00C0; #100;
A = 16'h008A; B = 16'h00C1; #100;
A = 16'h008A; B = 16'h00C2; #100;
A = 16'h008A; B = 16'h00C3; #100;
A = 16'h008A; B = 16'h00C4; #100;
A = 16'h008A; B = 16'h00C5; #100;
A = 16'h008A; B = 16'h00C6; #100;
A = 16'h008A; B = 16'h00C7; #100;
A = 16'h008A; B = 16'h00C8; #100;
A = 16'h008A; B = 16'h00C9; #100;
A = 16'h008A; B = 16'h00CA; #100;
A = 16'h008A; B = 16'h00CB; #100;
A = 16'h008A; B = 16'h00CC; #100;
A = 16'h008A; B = 16'h00CD; #100;
A = 16'h008A; B = 16'h00CE; #100;
A = 16'h008A; B = 16'h00CF; #100;
A = 16'h008A; B = 16'h00D0; #100;
A = 16'h008A; B = 16'h00D1; #100;
A = 16'h008A; B = 16'h00D2; #100;
A = 16'h008A; B = 16'h00D3; #100;
A = 16'h008A; B = 16'h00D4; #100;
A = 16'h008A; B = 16'h00D5; #100;
A = 16'h008A; B = 16'h00D6; #100;
A = 16'h008A; B = 16'h00D7; #100;
A = 16'h008A; B = 16'h00D8; #100;
A = 16'h008A; B = 16'h00D9; #100;
A = 16'h008A; B = 16'h00DA; #100;
A = 16'h008A; B = 16'h00DB; #100;
A = 16'h008A; B = 16'h00DC; #100;
A = 16'h008A; B = 16'h00DD; #100;
A = 16'h008A; B = 16'h00DE; #100;
A = 16'h008A; B = 16'h00DF; #100;
A = 16'h008A; B = 16'h00E0; #100;
A = 16'h008A; B = 16'h00E1; #100;
A = 16'h008A; B = 16'h00E2; #100;
A = 16'h008A; B = 16'h00E3; #100;
A = 16'h008A; B = 16'h00E4; #100;
A = 16'h008A; B = 16'h00E5; #100;
A = 16'h008A; B = 16'h00E6; #100;
A = 16'h008A; B = 16'h00E7; #100;
A = 16'h008A; B = 16'h00E8; #100;
A = 16'h008A; B = 16'h00E9; #100;
A = 16'h008A; B = 16'h00EA; #100;
A = 16'h008A; B = 16'h00EB; #100;
A = 16'h008A; B = 16'h00EC; #100;
A = 16'h008A; B = 16'h00ED; #100;
A = 16'h008A; B = 16'h00EE; #100;
A = 16'h008A; B = 16'h00EF; #100;
A = 16'h008A; B = 16'h00F0; #100;
A = 16'h008A; B = 16'h00F1; #100;
A = 16'h008A; B = 16'h00F2; #100;
A = 16'h008A; B = 16'h00F3; #100;
A = 16'h008A; B = 16'h00F4; #100;
A = 16'h008A; B = 16'h00F5; #100;
A = 16'h008A; B = 16'h00F6; #100;
A = 16'h008A; B = 16'h00F7; #100;
A = 16'h008A; B = 16'h00F8; #100;
A = 16'h008A; B = 16'h00F9; #100;
A = 16'h008A; B = 16'h00FA; #100;
A = 16'h008A; B = 16'h00FB; #100;
A = 16'h008A; B = 16'h00FC; #100;
A = 16'h008A; B = 16'h00FD; #100;
A = 16'h008A; B = 16'h00FE; #100;
A = 16'h008A; B = 16'h00FF; #100;
A = 16'h008B; B = 16'h000; #100;
A = 16'h008B; B = 16'h001; #100;
A = 16'h008B; B = 16'h002; #100;
A = 16'h008B; B = 16'h003; #100;
A = 16'h008B; B = 16'h004; #100;
A = 16'h008B; B = 16'h005; #100;
A = 16'h008B; B = 16'h006; #100;
A = 16'h008B; B = 16'h007; #100;
A = 16'h008B; B = 16'h008; #100;
A = 16'h008B; B = 16'h009; #100;
A = 16'h008B; B = 16'h00A; #100;
A = 16'h008B; B = 16'h00B; #100;
A = 16'h008B; B = 16'h00C; #100;
A = 16'h008B; B = 16'h00D; #100;
A = 16'h008B; B = 16'h00E; #100;
A = 16'h008B; B = 16'h00F; #100;
A = 16'h008B; B = 16'h0010; #100;
A = 16'h008B; B = 16'h0011; #100;
A = 16'h008B; B = 16'h0012; #100;
A = 16'h008B; B = 16'h0013; #100;
A = 16'h008B; B = 16'h0014; #100;
A = 16'h008B; B = 16'h0015; #100;
A = 16'h008B; B = 16'h0016; #100;
A = 16'h008B; B = 16'h0017; #100;
A = 16'h008B; B = 16'h0018; #100;
A = 16'h008B; B = 16'h0019; #100;
A = 16'h008B; B = 16'h001A; #100;
A = 16'h008B; B = 16'h001B; #100;
A = 16'h008B; B = 16'h001C; #100;
A = 16'h008B; B = 16'h001D; #100;
A = 16'h008B; B = 16'h001E; #100;
A = 16'h008B; B = 16'h001F; #100;
A = 16'h008B; B = 16'h0020; #100;
A = 16'h008B; B = 16'h0021; #100;
A = 16'h008B; B = 16'h0022; #100;
A = 16'h008B; B = 16'h0023; #100;
A = 16'h008B; B = 16'h0024; #100;
A = 16'h008B; B = 16'h0025; #100;
A = 16'h008B; B = 16'h0026; #100;
A = 16'h008B; B = 16'h0027; #100;
A = 16'h008B; B = 16'h0028; #100;
A = 16'h008B; B = 16'h0029; #100;
A = 16'h008B; B = 16'h002A; #100;
A = 16'h008B; B = 16'h002B; #100;
A = 16'h008B; B = 16'h002C; #100;
A = 16'h008B; B = 16'h002D; #100;
A = 16'h008B; B = 16'h002E; #100;
A = 16'h008B; B = 16'h002F; #100;
A = 16'h008B; B = 16'h0030; #100;
A = 16'h008B; B = 16'h0031; #100;
A = 16'h008B; B = 16'h0032; #100;
A = 16'h008B; B = 16'h0033; #100;
A = 16'h008B; B = 16'h0034; #100;
A = 16'h008B; B = 16'h0035; #100;
A = 16'h008B; B = 16'h0036; #100;
A = 16'h008B; B = 16'h0037; #100;
A = 16'h008B; B = 16'h0038; #100;
A = 16'h008B; B = 16'h0039; #100;
A = 16'h008B; B = 16'h003A; #100;
A = 16'h008B; B = 16'h003B; #100;
A = 16'h008B; B = 16'h003C; #100;
A = 16'h008B; B = 16'h003D; #100;
A = 16'h008B; B = 16'h003E; #100;
A = 16'h008B; B = 16'h003F; #100;
A = 16'h008B; B = 16'h0040; #100;
A = 16'h008B; B = 16'h0041; #100;
A = 16'h008B; B = 16'h0042; #100;
A = 16'h008B; B = 16'h0043; #100;
A = 16'h008B; B = 16'h0044; #100;
A = 16'h008B; B = 16'h0045; #100;
A = 16'h008B; B = 16'h0046; #100;
A = 16'h008B; B = 16'h0047; #100;
A = 16'h008B; B = 16'h0048; #100;
A = 16'h008B; B = 16'h0049; #100;
A = 16'h008B; B = 16'h004A; #100;
A = 16'h008B; B = 16'h004B; #100;
A = 16'h008B; B = 16'h004C; #100;
A = 16'h008B; B = 16'h004D; #100;
A = 16'h008B; B = 16'h004E; #100;
A = 16'h008B; B = 16'h004F; #100;
A = 16'h008B; B = 16'h0050; #100;
A = 16'h008B; B = 16'h0051; #100;
A = 16'h008B; B = 16'h0052; #100;
A = 16'h008B; B = 16'h0053; #100;
A = 16'h008B; B = 16'h0054; #100;
A = 16'h008B; B = 16'h0055; #100;
A = 16'h008B; B = 16'h0056; #100;
A = 16'h008B; B = 16'h0057; #100;
A = 16'h008B; B = 16'h0058; #100;
A = 16'h008B; B = 16'h0059; #100;
A = 16'h008B; B = 16'h005A; #100;
A = 16'h008B; B = 16'h005B; #100;
A = 16'h008B; B = 16'h005C; #100;
A = 16'h008B; B = 16'h005D; #100;
A = 16'h008B; B = 16'h005E; #100;
A = 16'h008B; B = 16'h005F; #100;
A = 16'h008B; B = 16'h0060; #100;
A = 16'h008B; B = 16'h0061; #100;
A = 16'h008B; B = 16'h0062; #100;
A = 16'h008B; B = 16'h0063; #100;
A = 16'h008B; B = 16'h0064; #100;
A = 16'h008B; B = 16'h0065; #100;
A = 16'h008B; B = 16'h0066; #100;
A = 16'h008B; B = 16'h0067; #100;
A = 16'h008B; B = 16'h0068; #100;
A = 16'h008B; B = 16'h0069; #100;
A = 16'h008B; B = 16'h006A; #100;
A = 16'h008B; B = 16'h006B; #100;
A = 16'h008B; B = 16'h006C; #100;
A = 16'h008B; B = 16'h006D; #100;
A = 16'h008B; B = 16'h006E; #100;
A = 16'h008B; B = 16'h006F; #100;
A = 16'h008B; B = 16'h0070; #100;
A = 16'h008B; B = 16'h0071; #100;
A = 16'h008B; B = 16'h0072; #100;
A = 16'h008B; B = 16'h0073; #100;
A = 16'h008B; B = 16'h0074; #100;
A = 16'h008B; B = 16'h0075; #100;
A = 16'h008B; B = 16'h0076; #100;
A = 16'h008B; B = 16'h0077; #100;
A = 16'h008B; B = 16'h0078; #100;
A = 16'h008B; B = 16'h0079; #100;
A = 16'h008B; B = 16'h007A; #100;
A = 16'h008B; B = 16'h007B; #100;
A = 16'h008B; B = 16'h007C; #100;
A = 16'h008B; B = 16'h007D; #100;
A = 16'h008B; B = 16'h007E; #100;
A = 16'h008B; B = 16'h007F; #100;
A = 16'h008B; B = 16'h0080; #100;
A = 16'h008B; B = 16'h0081; #100;
A = 16'h008B; B = 16'h0082; #100;
A = 16'h008B; B = 16'h0083; #100;
A = 16'h008B; B = 16'h0084; #100;
A = 16'h008B; B = 16'h0085; #100;
A = 16'h008B; B = 16'h0086; #100;
A = 16'h008B; B = 16'h0087; #100;
A = 16'h008B; B = 16'h0088; #100;
A = 16'h008B; B = 16'h0089; #100;
A = 16'h008B; B = 16'h008A; #100;
A = 16'h008B; B = 16'h008B; #100;
A = 16'h008B; B = 16'h008C; #100;
A = 16'h008B; B = 16'h008D; #100;
A = 16'h008B; B = 16'h008E; #100;
A = 16'h008B; B = 16'h008F; #100;
A = 16'h008B; B = 16'h0090; #100;
A = 16'h008B; B = 16'h0091; #100;
A = 16'h008B; B = 16'h0092; #100;
A = 16'h008B; B = 16'h0093; #100;
A = 16'h008B; B = 16'h0094; #100;
A = 16'h008B; B = 16'h0095; #100;
A = 16'h008B; B = 16'h0096; #100;
A = 16'h008B; B = 16'h0097; #100;
A = 16'h008B; B = 16'h0098; #100;
A = 16'h008B; B = 16'h0099; #100;
A = 16'h008B; B = 16'h009A; #100;
A = 16'h008B; B = 16'h009B; #100;
A = 16'h008B; B = 16'h009C; #100;
A = 16'h008B; B = 16'h009D; #100;
A = 16'h008B; B = 16'h009E; #100;
A = 16'h008B; B = 16'h009F; #100;
A = 16'h008B; B = 16'h00A0; #100;
A = 16'h008B; B = 16'h00A1; #100;
A = 16'h008B; B = 16'h00A2; #100;
A = 16'h008B; B = 16'h00A3; #100;
A = 16'h008B; B = 16'h00A4; #100;
A = 16'h008B; B = 16'h00A5; #100;
A = 16'h008B; B = 16'h00A6; #100;
A = 16'h008B; B = 16'h00A7; #100;
A = 16'h008B; B = 16'h00A8; #100;
A = 16'h008B; B = 16'h00A9; #100;
A = 16'h008B; B = 16'h00AA; #100;
A = 16'h008B; B = 16'h00AB; #100;
A = 16'h008B; B = 16'h00AC; #100;
A = 16'h008B; B = 16'h00AD; #100;
A = 16'h008B; B = 16'h00AE; #100;
A = 16'h008B; B = 16'h00AF; #100;
A = 16'h008B; B = 16'h00B0; #100;
A = 16'h008B; B = 16'h00B1; #100;
A = 16'h008B; B = 16'h00B2; #100;
A = 16'h008B; B = 16'h00B3; #100;
A = 16'h008B; B = 16'h00B4; #100;
A = 16'h008B; B = 16'h00B5; #100;
A = 16'h008B; B = 16'h00B6; #100;
A = 16'h008B; B = 16'h00B7; #100;
A = 16'h008B; B = 16'h00B8; #100;
A = 16'h008B; B = 16'h00B9; #100;
A = 16'h008B; B = 16'h00BA; #100;
A = 16'h008B; B = 16'h00BB; #100;
A = 16'h008B; B = 16'h00BC; #100;
A = 16'h008B; B = 16'h00BD; #100;
A = 16'h008B; B = 16'h00BE; #100;
A = 16'h008B; B = 16'h00BF; #100;
A = 16'h008B; B = 16'h00C0; #100;
A = 16'h008B; B = 16'h00C1; #100;
A = 16'h008B; B = 16'h00C2; #100;
A = 16'h008B; B = 16'h00C3; #100;
A = 16'h008B; B = 16'h00C4; #100;
A = 16'h008B; B = 16'h00C5; #100;
A = 16'h008B; B = 16'h00C6; #100;
A = 16'h008B; B = 16'h00C7; #100;
A = 16'h008B; B = 16'h00C8; #100;
A = 16'h008B; B = 16'h00C9; #100;
A = 16'h008B; B = 16'h00CA; #100;
A = 16'h008B; B = 16'h00CB; #100;
A = 16'h008B; B = 16'h00CC; #100;
A = 16'h008B; B = 16'h00CD; #100;
A = 16'h008B; B = 16'h00CE; #100;
A = 16'h008B; B = 16'h00CF; #100;
A = 16'h008B; B = 16'h00D0; #100;
A = 16'h008B; B = 16'h00D1; #100;
A = 16'h008B; B = 16'h00D2; #100;
A = 16'h008B; B = 16'h00D3; #100;
A = 16'h008B; B = 16'h00D4; #100;
A = 16'h008B; B = 16'h00D5; #100;
A = 16'h008B; B = 16'h00D6; #100;
A = 16'h008B; B = 16'h00D7; #100;
A = 16'h008B; B = 16'h00D8; #100;
A = 16'h008B; B = 16'h00D9; #100;
A = 16'h008B; B = 16'h00DA; #100;
A = 16'h008B; B = 16'h00DB; #100;
A = 16'h008B; B = 16'h00DC; #100;
A = 16'h008B; B = 16'h00DD; #100;
A = 16'h008B; B = 16'h00DE; #100;
A = 16'h008B; B = 16'h00DF; #100;
A = 16'h008B; B = 16'h00E0; #100;
A = 16'h008B; B = 16'h00E1; #100;
A = 16'h008B; B = 16'h00E2; #100;
A = 16'h008B; B = 16'h00E3; #100;
A = 16'h008B; B = 16'h00E4; #100;
A = 16'h008B; B = 16'h00E5; #100;
A = 16'h008B; B = 16'h00E6; #100;
A = 16'h008B; B = 16'h00E7; #100;
A = 16'h008B; B = 16'h00E8; #100;
A = 16'h008B; B = 16'h00E9; #100;
A = 16'h008B; B = 16'h00EA; #100;
A = 16'h008B; B = 16'h00EB; #100;
A = 16'h008B; B = 16'h00EC; #100;
A = 16'h008B; B = 16'h00ED; #100;
A = 16'h008B; B = 16'h00EE; #100;
A = 16'h008B; B = 16'h00EF; #100;
A = 16'h008B; B = 16'h00F0; #100;
A = 16'h008B; B = 16'h00F1; #100;
A = 16'h008B; B = 16'h00F2; #100;
A = 16'h008B; B = 16'h00F3; #100;
A = 16'h008B; B = 16'h00F4; #100;
A = 16'h008B; B = 16'h00F5; #100;
A = 16'h008B; B = 16'h00F6; #100;
A = 16'h008B; B = 16'h00F7; #100;
A = 16'h008B; B = 16'h00F8; #100;
A = 16'h008B; B = 16'h00F9; #100;
A = 16'h008B; B = 16'h00FA; #100;
A = 16'h008B; B = 16'h00FB; #100;
A = 16'h008B; B = 16'h00FC; #100;
A = 16'h008B; B = 16'h00FD; #100;
A = 16'h008B; B = 16'h00FE; #100;
A = 16'h008B; B = 16'h00FF; #100;
A = 16'h008C; B = 16'h000; #100;
A = 16'h008C; B = 16'h001; #100;
A = 16'h008C; B = 16'h002; #100;
A = 16'h008C; B = 16'h003; #100;
A = 16'h008C; B = 16'h004; #100;
A = 16'h008C; B = 16'h005; #100;
A = 16'h008C; B = 16'h006; #100;
A = 16'h008C; B = 16'h007; #100;
A = 16'h008C; B = 16'h008; #100;
A = 16'h008C; B = 16'h009; #100;
A = 16'h008C; B = 16'h00A; #100;
A = 16'h008C; B = 16'h00B; #100;
A = 16'h008C; B = 16'h00C; #100;
A = 16'h008C; B = 16'h00D; #100;
A = 16'h008C; B = 16'h00E; #100;
A = 16'h008C; B = 16'h00F; #100;
A = 16'h008C; B = 16'h0010; #100;
A = 16'h008C; B = 16'h0011; #100;
A = 16'h008C; B = 16'h0012; #100;
A = 16'h008C; B = 16'h0013; #100;
A = 16'h008C; B = 16'h0014; #100;
A = 16'h008C; B = 16'h0015; #100;
A = 16'h008C; B = 16'h0016; #100;
A = 16'h008C; B = 16'h0017; #100;
A = 16'h008C; B = 16'h0018; #100;
A = 16'h008C; B = 16'h0019; #100;
A = 16'h008C; B = 16'h001A; #100;
A = 16'h008C; B = 16'h001B; #100;
A = 16'h008C; B = 16'h001C; #100;
A = 16'h008C; B = 16'h001D; #100;
A = 16'h008C; B = 16'h001E; #100;
A = 16'h008C; B = 16'h001F; #100;
A = 16'h008C; B = 16'h0020; #100;
A = 16'h008C; B = 16'h0021; #100;
A = 16'h008C; B = 16'h0022; #100;
A = 16'h008C; B = 16'h0023; #100;
A = 16'h008C; B = 16'h0024; #100;
A = 16'h008C; B = 16'h0025; #100;
A = 16'h008C; B = 16'h0026; #100;
A = 16'h008C; B = 16'h0027; #100;
A = 16'h008C; B = 16'h0028; #100;
A = 16'h008C; B = 16'h0029; #100;
A = 16'h008C; B = 16'h002A; #100;
A = 16'h008C; B = 16'h002B; #100;
A = 16'h008C; B = 16'h002C; #100;
A = 16'h008C; B = 16'h002D; #100;
A = 16'h008C; B = 16'h002E; #100;
A = 16'h008C; B = 16'h002F; #100;
A = 16'h008C; B = 16'h0030; #100;
A = 16'h008C; B = 16'h0031; #100;
A = 16'h008C; B = 16'h0032; #100;
A = 16'h008C; B = 16'h0033; #100;
A = 16'h008C; B = 16'h0034; #100;
A = 16'h008C; B = 16'h0035; #100;
A = 16'h008C; B = 16'h0036; #100;
A = 16'h008C; B = 16'h0037; #100;
A = 16'h008C; B = 16'h0038; #100;
A = 16'h008C; B = 16'h0039; #100;
A = 16'h008C; B = 16'h003A; #100;
A = 16'h008C; B = 16'h003B; #100;
A = 16'h008C; B = 16'h003C; #100;
A = 16'h008C; B = 16'h003D; #100;
A = 16'h008C; B = 16'h003E; #100;
A = 16'h008C; B = 16'h003F; #100;
A = 16'h008C; B = 16'h0040; #100;
A = 16'h008C; B = 16'h0041; #100;
A = 16'h008C; B = 16'h0042; #100;
A = 16'h008C; B = 16'h0043; #100;
A = 16'h008C; B = 16'h0044; #100;
A = 16'h008C; B = 16'h0045; #100;
A = 16'h008C; B = 16'h0046; #100;
A = 16'h008C; B = 16'h0047; #100;
A = 16'h008C; B = 16'h0048; #100;
A = 16'h008C; B = 16'h0049; #100;
A = 16'h008C; B = 16'h004A; #100;
A = 16'h008C; B = 16'h004B; #100;
A = 16'h008C; B = 16'h004C; #100;
A = 16'h008C; B = 16'h004D; #100;
A = 16'h008C; B = 16'h004E; #100;
A = 16'h008C; B = 16'h004F; #100;
A = 16'h008C; B = 16'h0050; #100;
A = 16'h008C; B = 16'h0051; #100;
A = 16'h008C; B = 16'h0052; #100;
A = 16'h008C; B = 16'h0053; #100;
A = 16'h008C; B = 16'h0054; #100;
A = 16'h008C; B = 16'h0055; #100;
A = 16'h008C; B = 16'h0056; #100;
A = 16'h008C; B = 16'h0057; #100;
A = 16'h008C; B = 16'h0058; #100;
A = 16'h008C; B = 16'h0059; #100;
A = 16'h008C; B = 16'h005A; #100;
A = 16'h008C; B = 16'h005B; #100;
A = 16'h008C; B = 16'h005C; #100;
A = 16'h008C; B = 16'h005D; #100;
A = 16'h008C; B = 16'h005E; #100;
A = 16'h008C; B = 16'h005F; #100;
A = 16'h008C; B = 16'h0060; #100;
A = 16'h008C; B = 16'h0061; #100;
A = 16'h008C; B = 16'h0062; #100;
A = 16'h008C; B = 16'h0063; #100;
A = 16'h008C; B = 16'h0064; #100;
A = 16'h008C; B = 16'h0065; #100;
A = 16'h008C; B = 16'h0066; #100;
A = 16'h008C; B = 16'h0067; #100;
A = 16'h008C; B = 16'h0068; #100;
A = 16'h008C; B = 16'h0069; #100;
A = 16'h008C; B = 16'h006A; #100;
A = 16'h008C; B = 16'h006B; #100;
A = 16'h008C; B = 16'h006C; #100;
A = 16'h008C; B = 16'h006D; #100;
A = 16'h008C; B = 16'h006E; #100;
A = 16'h008C; B = 16'h006F; #100;
A = 16'h008C; B = 16'h0070; #100;
A = 16'h008C; B = 16'h0071; #100;
A = 16'h008C; B = 16'h0072; #100;
A = 16'h008C; B = 16'h0073; #100;
A = 16'h008C; B = 16'h0074; #100;
A = 16'h008C; B = 16'h0075; #100;
A = 16'h008C; B = 16'h0076; #100;
A = 16'h008C; B = 16'h0077; #100;
A = 16'h008C; B = 16'h0078; #100;
A = 16'h008C; B = 16'h0079; #100;
A = 16'h008C; B = 16'h007A; #100;
A = 16'h008C; B = 16'h007B; #100;
A = 16'h008C; B = 16'h007C; #100;
A = 16'h008C; B = 16'h007D; #100;
A = 16'h008C; B = 16'h007E; #100;
A = 16'h008C; B = 16'h007F; #100;
A = 16'h008C; B = 16'h0080; #100;
A = 16'h008C; B = 16'h0081; #100;
A = 16'h008C; B = 16'h0082; #100;
A = 16'h008C; B = 16'h0083; #100;
A = 16'h008C; B = 16'h0084; #100;
A = 16'h008C; B = 16'h0085; #100;
A = 16'h008C; B = 16'h0086; #100;
A = 16'h008C; B = 16'h0087; #100;
A = 16'h008C; B = 16'h0088; #100;
A = 16'h008C; B = 16'h0089; #100;
A = 16'h008C; B = 16'h008A; #100;
A = 16'h008C; B = 16'h008B; #100;
A = 16'h008C; B = 16'h008C; #100;
A = 16'h008C; B = 16'h008D; #100;
A = 16'h008C; B = 16'h008E; #100;
A = 16'h008C; B = 16'h008F; #100;
A = 16'h008C; B = 16'h0090; #100;
A = 16'h008C; B = 16'h0091; #100;
A = 16'h008C; B = 16'h0092; #100;
A = 16'h008C; B = 16'h0093; #100;
A = 16'h008C; B = 16'h0094; #100;
A = 16'h008C; B = 16'h0095; #100;
A = 16'h008C; B = 16'h0096; #100;
A = 16'h008C; B = 16'h0097; #100;
A = 16'h008C; B = 16'h0098; #100;
A = 16'h008C; B = 16'h0099; #100;
A = 16'h008C; B = 16'h009A; #100;
A = 16'h008C; B = 16'h009B; #100;
A = 16'h008C; B = 16'h009C; #100;
A = 16'h008C; B = 16'h009D; #100;
A = 16'h008C; B = 16'h009E; #100;
A = 16'h008C; B = 16'h009F; #100;
A = 16'h008C; B = 16'h00A0; #100;
A = 16'h008C; B = 16'h00A1; #100;
A = 16'h008C; B = 16'h00A2; #100;
A = 16'h008C; B = 16'h00A3; #100;
A = 16'h008C; B = 16'h00A4; #100;
A = 16'h008C; B = 16'h00A5; #100;
A = 16'h008C; B = 16'h00A6; #100;
A = 16'h008C; B = 16'h00A7; #100;
A = 16'h008C; B = 16'h00A8; #100;
A = 16'h008C; B = 16'h00A9; #100;
A = 16'h008C; B = 16'h00AA; #100;
A = 16'h008C; B = 16'h00AB; #100;
A = 16'h008C; B = 16'h00AC; #100;
A = 16'h008C; B = 16'h00AD; #100;
A = 16'h008C; B = 16'h00AE; #100;
A = 16'h008C; B = 16'h00AF; #100;
A = 16'h008C; B = 16'h00B0; #100;
A = 16'h008C; B = 16'h00B1; #100;
A = 16'h008C; B = 16'h00B2; #100;
A = 16'h008C; B = 16'h00B3; #100;
A = 16'h008C; B = 16'h00B4; #100;
A = 16'h008C; B = 16'h00B5; #100;
A = 16'h008C; B = 16'h00B6; #100;
A = 16'h008C; B = 16'h00B7; #100;
A = 16'h008C; B = 16'h00B8; #100;
A = 16'h008C; B = 16'h00B9; #100;
A = 16'h008C; B = 16'h00BA; #100;
A = 16'h008C; B = 16'h00BB; #100;
A = 16'h008C; B = 16'h00BC; #100;
A = 16'h008C; B = 16'h00BD; #100;
A = 16'h008C; B = 16'h00BE; #100;
A = 16'h008C; B = 16'h00BF; #100;
A = 16'h008C; B = 16'h00C0; #100;
A = 16'h008C; B = 16'h00C1; #100;
A = 16'h008C; B = 16'h00C2; #100;
A = 16'h008C; B = 16'h00C3; #100;
A = 16'h008C; B = 16'h00C4; #100;
A = 16'h008C; B = 16'h00C5; #100;
A = 16'h008C; B = 16'h00C6; #100;
A = 16'h008C; B = 16'h00C7; #100;
A = 16'h008C; B = 16'h00C8; #100;
A = 16'h008C; B = 16'h00C9; #100;
A = 16'h008C; B = 16'h00CA; #100;
A = 16'h008C; B = 16'h00CB; #100;
A = 16'h008C; B = 16'h00CC; #100;
A = 16'h008C; B = 16'h00CD; #100;
A = 16'h008C; B = 16'h00CE; #100;
A = 16'h008C; B = 16'h00CF; #100;
A = 16'h008C; B = 16'h00D0; #100;
A = 16'h008C; B = 16'h00D1; #100;
A = 16'h008C; B = 16'h00D2; #100;
A = 16'h008C; B = 16'h00D3; #100;
A = 16'h008C; B = 16'h00D4; #100;
A = 16'h008C; B = 16'h00D5; #100;
A = 16'h008C; B = 16'h00D6; #100;
A = 16'h008C; B = 16'h00D7; #100;
A = 16'h008C; B = 16'h00D8; #100;
A = 16'h008C; B = 16'h00D9; #100;
A = 16'h008C; B = 16'h00DA; #100;
A = 16'h008C; B = 16'h00DB; #100;
A = 16'h008C; B = 16'h00DC; #100;
A = 16'h008C; B = 16'h00DD; #100;
A = 16'h008C; B = 16'h00DE; #100;
A = 16'h008C; B = 16'h00DF; #100;
A = 16'h008C; B = 16'h00E0; #100;
A = 16'h008C; B = 16'h00E1; #100;
A = 16'h008C; B = 16'h00E2; #100;
A = 16'h008C; B = 16'h00E3; #100;
A = 16'h008C; B = 16'h00E4; #100;
A = 16'h008C; B = 16'h00E5; #100;
A = 16'h008C; B = 16'h00E6; #100;
A = 16'h008C; B = 16'h00E7; #100;
A = 16'h008C; B = 16'h00E8; #100;
A = 16'h008C; B = 16'h00E9; #100;
A = 16'h008C; B = 16'h00EA; #100;
A = 16'h008C; B = 16'h00EB; #100;
A = 16'h008C; B = 16'h00EC; #100;
A = 16'h008C; B = 16'h00ED; #100;
A = 16'h008C; B = 16'h00EE; #100;
A = 16'h008C; B = 16'h00EF; #100;
A = 16'h008C; B = 16'h00F0; #100;
A = 16'h008C; B = 16'h00F1; #100;
A = 16'h008C; B = 16'h00F2; #100;
A = 16'h008C; B = 16'h00F3; #100;
A = 16'h008C; B = 16'h00F4; #100;
A = 16'h008C; B = 16'h00F5; #100;
A = 16'h008C; B = 16'h00F6; #100;
A = 16'h008C; B = 16'h00F7; #100;
A = 16'h008C; B = 16'h00F8; #100;
A = 16'h008C; B = 16'h00F9; #100;
A = 16'h008C; B = 16'h00FA; #100;
A = 16'h008C; B = 16'h00FB; #100;
A = 16'h008C; B = 16'h00FC; #100;
A = 16'h008C; B = 16'h00FD; #100;
A = 16'h008C; B = 16'h00FE; #100;
A = 16'h008C; B = 16'h00FF; #100;
A = 16'h008D; B = 16'h000; #100;
A = 16'h008D; B = 16'h001; #100;
A = 16'h008D; B = 16'h002; #100;
A = 16'h008D; B = 16'h003; #100;
A = 16'h008D; B = 16'h004; #100;
A = 16'h008D; B = 16'h005; #100;
A = 16'h008D; B = 16'h006; #100;
A = 16'h008D; B = 16'h007; #100;
A = 16'h008D; B = 16'h008; #100;
A = 16'h008D; B = 16'h009; #100;
A = 16'h008D; B = 16'h00A; #100;
A = 16'h008D; B = 16'h00B; #100;
A = 16'h008D; B = 16'h00C; #100;
A = 16'h008D; B = 16'h00D; #100;
A = 16'h008D; B = 16'h00E; #100;
A = 16'h008D; B = 16'h00F; #100;
A = 16'h008D; B = 16'h0010; #100;
A = 16'h008D; B = 16'h0011; #100;
A = 16'h008D; B = 16'h0012; #100;
A = 16'h008D; B = 16'h0013; #100;
A = 16'h008D; B = 16'h0014; #100;
A = 16'h008D; B = 16'h0015; #100;
A = 16'h008D; B = 16'h0016; #100;
A = 16'h008D; B = 16'h0017; #100;
A = 16'h008D; B = 16'h0018; #100;
A = 16'h008D; B = 16'h0019; #100;
A = 16'h008D; B = 16'h001A; #100;
A = 16'h008D; B = 16'h001B; #100;
A = 16'h008D; B = 16'h001C; #100;
A = 16'h008D; B = 16'h001D; #100;
A = 16'h008D; B = 16'h001E; #100;
A = 16'h008D; B = 16'h001F; #100;
A = 16'h008D; B = 16'h0020; #100;
A = 16'h008D; B = 16'h0021; #100;
A = 16'h008D; B = 16'h0022; #100;
A = 16'h008D; B = 16'h0023; #100;
A = 16'h008D; B = 16'h0024; #100;
A = 16'h008D; B = 16'h0025; #100;
A = 16'h008D; B = 16'h0026; #100;
A = 16'h008D; B = 16'h0027; #100;
A = 16'h008D; B = 16'h0028; #100;
A = 16'h008D; B = 16'h0029; #100;
A = 16'h008D; B = 16'h002A; #100;
A = 16'h008D; B = 16'h002B; #100;
A = 16'h008D; B = 16'h002C; #100;
A = 16'h008D; B = 16'h002D; #100;
A = 16'h008D; B = 16'h002E; #100;
A = 16'h008D; B = 16'h002F; #100;
A = 16'h008D; B = 16'h0030; #100;
A = 16'h008D; B = 16'h0031; #100;
A = 16'h008D; B = 16'h0032; #100;
A = 16'h008D; B = 16'h0033; #100;
A = 16'h008D; B = 16'h0034; #100;
A = 16'h008D; B = 16'h0035; #100;
A = 16'h008D; B = 16'h0036; #100;
A = 16'h008D; B = 16'h0037; #100;
A = 16'h008D; B = 16'h0038; #100;
A = 16'h008D; B = 16'h0039; #100;
A = 16'h008D; B = 16'h003A; #100;
A = 16'h008D; B = 16'h003B; #100;
A = 16'h008D; B = 16'h003C; #100;
A = 16'h008D; B = 16'h003D; #100;
A = 16'h008D; B = 16'h003E; #100;
A = 16'h008D; B = 16'h003F; #100;
A = 16'h008D; B = 16'h0040; #100;
A = 16'h008D; B = 16'h0041; #100;
A = 16'h008D; B = 16'h0042; #100;
A = 16'h008D; B = 16'h0043; #100;
A = 16'h008D; B = 16'h0044; #100;
A = 16'h008D; B = 16'h0045; #100;
A = 16'h008D; B = 16'h0046; #100;
A = 16'h008D; B = 16'h0047; #100;
A = 16'h008D; B = 16'h0048; #100;
A = 16'h008D; B = 16'h0049; #100;
A = 16'h008D; B = 16'h004A; #100;
A = 16'h008D; B = 16'h004B; #100;
A = 16'h008D; B = 16'h004C; #100;
A = 16'h008D; B = 16'h004D; #100;
A = 16'h008D; B = 16'h004E; #100;
A = 16'h008D; B = 16'h004F; #100;
A = 16'h008D; B = 16'h0050; #100;
A = 16'h008D; B = 16'h0051; #100;
A = 16'h008D; B = 16'h0052; #100;
A = 16'h008D; B = 16'h0053; #100;
A = 16'h008D; B = 16'h0054; #100;
A = 16'h008D; B = 16'h0055; #100;
A = 16'h008D; B = 16'h0056; #100;
A = 16'h008D; B = 16'h0057; #100;
A = 16'h008D; B = 16'h0058; #100;
A = 16'h008D; B = 16'h0059; #100;
A = 16'h008D; B = 16'h005A; #100;
A = 16'h008D; B = 16'h005B; #100;
A = 16'h008D; B = 16'h005C; #100;
A = 16'h008D; B = 16'h005D; #100;
A = 16'h008D; B = 16'h005E; #100;
A = 16'h008D; B = 16'h005F; #100;
A = 16'h008D; B = 16'h0060; #100;
A = 16'h008D; B = 16'h0061; #100;
A = 16'h008D; B = 16'h0062; #100;
A = 16'h008D; B = 16'h0063; #100;
A = 16'h008D; B = 16'h0064; #100;
A = 16'h008D; B = 16'h0065; #100;
A = 16'h008D; B = 16'h0066; #100;
A = 16'h008D; B = 16'h0067; #100;
A = 16'h008D; B = 16'h0068; #100;
A = 16'h008D; B = 16'h0069; #100;
A = 16'h008D; B = 16'h006A; #100;
A = 16'h008D; B = 16'h006B; #100;
A = 16'h008D; B = 16'h006C; #100;
A = 16'h008D; B = 16'h006D; #100;
A = 16'h008D; B = 16'h006E; #100;
A = 16'h008D; B = 16'h006F; #100;
A = 16'h008D; B = 16'h0070; #100;
A = 16'h008D; B = 16'h0071; #100;
A = 16'h008D; B = 16'h0072; #100;
A = 16'h008D; B = 16'h0073; #100;
A = 16'h008D; B = 16'h0074; #100;
A = 16'h008D; B = 16'h0075; #100;
A = 16'h008D; B = 16'h0076; #100;
A = 16'h008D; B = 16'h0077; #100;
A = 16'h008D; B = 16'h0078; #100;
A = 16'h008D; B = 16'h0079; #100;
A = 16'h008D; B = 16'h007A; #100;
A = 16'h008D; B = 16'h007B; #100;
A = 16'h008D; B = 16'h007C; #100;
A = 16'h008D; B = 16'h007D; #100;
A = 16'h008D; B = 16'h007E; #100;
A = 16'h008D; B = 16'h007F; #100;
A = 16'h008D; B = 16'h0080; #100;
A = 16'h008D; B = 16'h0081; #100;
A = 16'h008D; B = 16'h0082; #100;
A = 16'h008D; B = 16'h0083; #100;
A = 16'h008D; B = 16'h0084; #100;
A = 16'h008D; B = 16'h0085; #100;
A = 16'h008D; B = 16'h0086; #100;
A = 16'h008D; B = 16'h0087; #100;
A = 16'h008D; B = 16'h0088; #100;
A = 16'h008D; B = 16'h0089; #100;
A = 16'h008D; B = 16'h008A; #100;
A = 16'h008D; B = 16'h008B; #100;
A = 16'h008D; B = 16'h008C; #100;
A = 16'h008D; B = 16'h008D; #100;
A = 16'h008D; B = 16'h008E; #100;
A = 16'h008D; B = 16'h008F; #100;
A = 16'h008D; B = 16'h0090; #100;
A = 16'h008D; B = 16'h0091; #100;
A = 16'h008D; B = 16'h0092; #100;
A = 16'h008D; B = 16'h0093; #100;
A = 16'h008D; B = 16'h0094; #100;
A = 16'h008D; B = 16'h0095; #100;
A = 16'h008D; B = 16'h0096; #100;
A = 16'h008D; B = 16'h0097; #100;
A = 16'h008D; B = 16'h0098; #100;
A = 16'h008D; B = 16'h0099; #100;
A = 16'h008D; B = 16'h009A; #100;
A = 16'h008D; B = 16'h009B; #100;
A = 16'h008D; B = 16'h009C; #100;
A = 16'h008D; B = 16'h009D; #100;
A = 16'h008D; B = 16'h009E; #100;
A = 16'h008D; B = 16'h009F; #100;
A = 16'h008D; B = 16'h00A0; #100;
A = 16'h008D; B = 16'h00A1; #100;
A = 16'h008D; B = 16'h00A2; #100;
A = 16'h008D; B = 16'h00A3; #100;
A = 16'h008D; B = 16'h00A4; #100;
A = 16'h008D; B = 16'h00A5; #100;
A = 16'h008D; B = 16'h00A6; #100;
A = 16'h008D; B = 16'h00A7; #100;
A = 16'h008D; B = 16'h00A8; #100;
A = 16'h008D; B = 16'h00A9; #100;
A = 16'h008D; B = 16'h00AA; #100;
A = 16'h008D; B = 16'h00AB; #100;
A = 16'h008D; B = 16'h00AC; #100;
A = 16'h008D; B = 16'h00AD; #100;
A = 16'h008D; B = 16'h00AE; #100;
A = 16'h008D; B = 16'h00AF; #100;
A = 16'h008D; B = 16'h00B0; #100;
A = 16'h008D; B = 16'h00B1; #100;
A = 16'h008D; B = 16'h00B2; #100;
A = 16'h008D; B = 16'h00B3; #100;
A = 16'h008D; B = 16'h00B4; #100;
A = 16'h008D; B = 16'h00B5; #100;
A = 16'h008D; B = 16'h00B6; #100;
A = 16'h008D; B = 16'h00B7; #100;
A = 16'h008D; B = 16'h00B8; #100;
A = 16'h008D; B = 16'h00B9; #100;
A = 16'h008D; B = 16'h00BA; #100;
A = 16'h008D; B = 16'h00BB; #100;
A = 16'h008D; B = 16'h00BC; #100;
A = 16'h008D; B = 16'h00BD; #100;
A = 16'h008D; B = 16'h00BE; #100;
A = 16'h008D; B = 16'h00BF; #100;
A = 16'h008D; B = 16'h00C0; #100;
A = 16'h008D; B = 16'h00C1; #100;
A = 16'h008D; B = 16'h00C2; #100;
A = 16'h008D; B = 16'h00C3; #100;
A = 16'h008D; B = 16'h00C4; #100;
A = 16'h008D; B = 16'h00C5; #100;
A = 16'h008D; B = 16'h00C6; #100;
A = 16'h008D; B = 16'h00C7; #100;
A = 16'h008D; B = 16'h00C8; #100;
A = 16'h008D; B = 16'h00C9; #100;
A = 16'h008D; B = 16'h00CA; #100;
A = 16'h008D; B = 16'h00CB; #100;
A = 16'h008D; B = 16'h00CC; #100;
A = 16'h008D; B = 16'h00CD; #100;
A = 16'h008D; B = 16'h00CE; #100;
A = 16'h008D; B = 16'h00CF; #100;
A = 16'h008D; B = 16'h00D0; #100;
A = 16'h008D; B = 16'h00D1; #100;
A = 16'h008D; B = 16'h00D2; #100;
A = 16'h008D; B = 16'h00D3; #100;
A = 16'h008D; B = 16'h00D4; #100;
A = 16'h008D; B = 16'h00D5; #100;
A = 16'h008D; B = 16'h00D6; #100;
A = 16'h008D; B = 16'h00D7; #100;
A = 16'h008D; B = 16'h00D8; #100;
A = 16'h008D; B = 16'h00D9; #100;
A = 16'h008D; B = 16'h00DA; #100;
A = 16'h008D; B = 16'h00DB; #100;
A = 16'h008D; B = 16'h00DC; #100;
A = 16'h008D; B = 16'h00DD; #100;
A = 16'h008D; B = 16'h00DE; #100;
A = 16'h008D; B = 16'h00DF; #100;
A = 16'h008D; B = 16'h00E0; #100;
A = 16'h008D; B = 16'h00E1; #100;
A = 16'h008D; B = 16'h00E2; #100;
A = 16'h008D; B = 16'h00E3; #100;
A = 16'h008D; B = 16'h00E4; #100;
A = 16'h008D; B = 16'h00E5; #100;
A = 16'h008D; B = 16'h00E6; #100;
A = 16'h008D; B = 16'h00E7; #100;
A = 16'h008D; B = 16'h00E8; #100;
A = 16'h008D; B = 16'h00E9; #100;
A = 16'h008D; B = 16'h00EA; #100;
A = 16'h008D; B = 16'h00EB; #100;
A = 16'h008D; B = 16'h00EC; #100;
A = 16'h008D; B = 16'h00ED; #100;
A = 16'h008D; B = 16'h00EE; #100;
A = 16'h008D; B = 16'h00EF; #100;
A = 16'h008D; B = 16'h00F0; #100;
A = 16'h008D; B = 16'h00F1; #100;
A = 16'h008D; B = 16'h00F2; #100;
A = 16'h008D; B = 16'h00F3; #100;
A = 16'h008D; B = 16'h00F4; #100;
A = 16'h008D; B = 16'h00F5; #100;
A = 16'h008D; B = 16'h00F6; #100;
A = 16'h008D; B = 16'h00F7; #100;
A = 16'h008D; B = 16'h00F8; #100;
A = 16'h008D; B = 16'h00F9; #100;
A = 16'h008D; B = 16'h00FA; #100;
A = 16'h008D; B = 16'h00FB; #100;
A = 16'h008D; B = 16'h00FC; #100;
A = 16'h008D; B = 16'h00FD; #100;
A = 16'h008D; B = 16'h00FE; #100;
A = 16'h008D; B = 16'h00FF; #100;
A = 16'h008E; B = 16'h000; #100;
A = 16'h008E; B = 16'h001; #100;
A = 16'h008E; B = 16'h002; #100;
A = 16'h008E; B = 16'h003; #100;
A = 16'h008E; B = 16'h004; #100;
A = 16'h008E; B = 16'h005; #100;
A = 16'h008E; B = 16'h006; #100;
A = 16'h008E; B = 16'h007; #100;
A = 16'h008E; B = 16'h008; #100;
A = 16'h008E; B = 16'h009; #100;
A = 16'h008E; B = 16'h00A; #100;
A = 16'h008E; B = 16'h00B; #100;
A = 16'h008E; B = 16'h00C; #100;
A = 16'h008E; B = 16'h00D; #100;
A = 16'h008E; B = 16'h00E; #100;
A = 16'h008E; B = 16'h00F; #100;
A = 16'h008E; B = 16'h0010; #100;
A = 16'h008E; B = 16'h0011; #100;
A = 16'h008E; B = 16'h0012; #100;
A = 16'h008E; B = 16'h0013; #100;
A = 16'h008E; B = 16'h0014; #100;
A = 16'h008E; B = 16'h0015; #100;
A = 16'h008E; B = 16'h0016; #100;
A = 16'h008E; B = 16'h0017; #100;
A = 16'h008E; B = 16'h0018; #100;
A = 16'h008E; B = 16'h0019; #100;
A = 16'h008E; B = 16'h001A; #100;
A = 16'h008E; B = 16'h001B; #100;
A = 16'h008E; B = 16'h001C; #100;
A = 16'h008E; B = 16'h001D; #100;
A = 16'h008E; B = 16'h001E; #100;
A = 16'h008E; B = 16'h001F; #100;
A = 16'h008E; B = 16'h0020; #100;
A = 16'h008E; B = 16'h0021; #100;
A = 16'h008E; B = 16'h0022; #100;
A = 16'h008E; B = 16'h0023; #100;
A = 16'h008E; B = 16'h0024; #100;
A = 16'h008E; B = 16'h0025; #100;
A = 16'h008E; B = 16'h0026; #100;
A = 16'h008E; B = 16'h0027; #100;
A = 16'h008E; B = 16'h0028; #100;
A = 16'h008E; B = 16'h0029; #100;
A = 16'h008E; B = 16'h002A; #100;
A = 16'h008E; B = 16'h002B; #100;
A = 16'h008E; B = 16'h002C; #100;
A = 16'h008E; B = 16'h002D; #100;
A = 16'h008E; B = 16'h002E; #100;
A = 16'h008E; B = 16'h002F; #100;
A = 16'h008E; B = 16'h0030; #100;
A = 16'h008E; B = 16'h0031; #100;
A = 16'h008E; B = 16'h0032; #100;
A = 16'h008E; B = 16'h0033; #100;
A = 16'h008E; B = 16'h0034; #100;
A = 16'h008E; B = 16'h0035; #100;
A = 16'h008E; B = 16'h0036; #100;
A = 16'h008E; B = 16'h0037; #100;
A = 16'h008E; B = 16'h0038; #100;
A = 16'h008E; B = 16'h0039; #100;
A = 16'h008E; B = 16'h003A; #100;
A = 16'h008E; B = 16'h003B; #100;
A = 16'h008E; B = 16'h003C; #100;
A = 16'h008E; B = 16'h003D; #100;
A = 16'h008E; B = 16'h003E; #100;
A = 16'h008E; B = 16'h003F; #100;
A = 16'h008E; B = 16'h0040; #100;
A = 16'h008E; B = 16'h0041; #100;
A = 16'h008E; B = 16'h0042; #100;
A = 16'h008E; B = 16'h0043; #100;
A = 16'h008E; B = 16'h0044; #100;
A = 16'h008E; B = 16'h0045; #100;
A = 16'h008E; B = 16'h0046; #100;
A = 16'h008E; B = 16'h0047; #100;
A = 16'h008E; B = 16'h0048; #100;
A = 16'h008E; B = 16'h0049; #100;
A = 16'h008E; B = 16'h004A; #100;
A = 16'h008E; B = 16'h004B; #100;
A = 16'h008E; B = 16'h004C; #100;
A = 16'h008E; B = 16'h004D; #100;
A = 16'h008E; B = 16'h004E; #100;
A = 16'h008E; B = 16'h004F; #100;
A = 16'h008E; B = 16'h0050; #100;
A = 16'h008E; B = 16'h0051; #100;
A = 16'h008E; B = 16'h0052; #100;
A = 16'h008E; B = 16'h0053; #100;
A = 16'h008E; B = 16'h0054; #100;
A = 16'h008E; B = 16'h0055; #100;
A = 16'h008E; B = 16'h0056; #100;
A = 16'h008E; B = 16'h0057; #100;
A = 16'h008E; B = 16'h0058; #100;
A = 16'h008E; B = 16'h0059; #100;
A = 16'h008E; B = 16'h005A; #100;
A = 16'h008E; B = 16'h005B; #100;
A = 16'h008E; B = 16'h005C; #100;
A = 16'h008E; B = 16'h005D; #100;
A = 16'h008E; B = 16'h005E; #100;
A = 16'h008E; B = 16'h005F; #100;
A = 16'h008E; B = 16'h0060; #100;
A = 16'h008E; B = 16'h0061; #100;
A = 16'h008E; B = 16'h0062; #100;
A = 16'h008E; B = 16'h0063; #100;
A = 16'h008E; B = 16'h0064; #100;
A = 16'h008E; B = 16'h0065; #100;
A = 16'h008E; B = 16'h0066; #100;
A = 16'h008E; B = 16'h0067; #100;
A = 16'h008E; B = 16'h0068; #100;
A = 16'h008E; B = 16'h0069; #100;
A = 16'h008E; B = 16'h006A; #100;
A = 16'h008E; B = 16'h006B; #100;
A = 16'h008E; B = 16'h006C; #100;
A = 16'h008E; B = 16'h006D; #100;
A = 16'h008E; B = 16'h006E; #100;
A = 16'h008E; B = 16'h006F; #100;
A = 16'h008E; B = 16'h0070; #100;
A = 16'h008E; B = 16'h0071; #100;
A = 16'h008E; B = 16'h0072; #100;
A = 16'h008E; B = 16'h0073; #100;
A = 16'h008E; B = 16'h0074; #100;
A = 16'h008E; B = 16'h0075; #100;
A = 16'h008E; B = 16'h0076; #100;
A = 16'h008E; B = 16'h0077; #100;
A = 16'h008E; B = 16'h0078; #100;
A = 16'h008E; B = 16'h0079; #100;
A = 16'h008E; B = 16'h007A; #100;
A = 16'h008E; B = 16'h007B; #100;
A = 16'h008E; B = 16'h007C; #100;
A = 16'h008E; B = 16'h007D; #100;
A = 16'h008E; B = 16'h007E; #100;
A = 16'h008E; B = 16'h007F; #100;
A = 16'h008E; B = 16'h0080; #100;
A = 16'h008E; B = 16'h0081; #100;
A = 16'h008E; B = 16'h0082; #100;
A = 16'h008E; B = 16'h0083; #100;
A = 16'h008E; B = 16'h0084; #100;
A = 16'h008E; B = 16'h0085; #100;
A = 16'h008E; B = 16'h0086; #100;
A = 16'h008E; B = 16'h0087; #100;
A = 16'h008E; B = 16'h0088; #100;
A = 16'h008E; B = 16'h0089; #100;
A = 16'h008E; B = 16'h008A; #100;
A = 16'h008E; B = 16'h008B; #100;
A = 16'h008E; B = 16'h008C; #100;
A = 16'h008E; B = 16'h008D; #100;
A = 16'h008E; B = 16'h008E; #100;
A = 16'h008E; B = 16'h008F; #100;
A = 16'h008E; B = 16'h0090; #100;
A = 16'h008E; B = 16'h0091; #100;
A = 16'h008E; B = 16'h0092; #100;
A = 16'h008E; B = 16'h0093; #100;
A = 16'h008E; B = 16'h0094; #100;
A = 16'h008E; B = 16'h0095; #100;
A = 16'h008E; B = 16'h0096; #100;
A = 16'h008E; B = 16'h0097; #100;
A = 16'h008E; B = 16'h0098; #100;
A = 16'h008E; B = 16'h0099; #100;
A = 16'h008E; B = 16'h009A; #100;
A = 16'h008E; B = 16'h009B; #100;
A = 16'h008E; B = 16'h009C; #100;
A = 16'h008E; B = 16'h009D; #100;
A = 16'h008E; B = 16'h009E; #100;
A = 16'h008E; B = 16'h009F; #100;
A = 16'h008E; B = 16'h00A0; #100;
A = 16'h008E; B = 16'h00A1; #100;
A = 16'h008E; B = 16'h00A2; #100;
A = 16'h008E; B = 16'h00A3; #100;
A = 16'h008E; B = 16'h00A4; #100;
A = 16'h008E; B = 16'h00A5; #100;
A = 16'h008E; B = 16'h00A6; #100;
A = 16'h008E; B = 16'h00A7; #100;
A = 16'h008E; B = 16'h00A8; #100;
A = 16'h008E; B = 16'h00A9; #100;
A = 16'h008E; B = 16'h00AA; #100;
A = 16'h008E; B = 16'h00AB; #100;
A = 16'h008E; B = 16'h00AC; #100;
A = 16'h008E; B = 16'h00AD; #100;
A = 16'h008E; B = 16'h00AE; #100;
A = 16'h008E; B = 16'h00AF; #100;
A = 16'h008E; B = 16'h00B0; #100;
A = 16'h008E; B = 16'h00B1; #100;
A = 16'h008E; B = 16'h00B2; #100;
A = 16'h008E; B = 16'h00B3; #100;
A = 16'h008E; B = 16'h00B4; #100;
A = 16'h008E; B = 16'h00B5; #100;
A = 16'h008E; B = 16'h00B6; #100;
A = 16'h008E; B = 16'h00B7; #100;
A = 16'h008E; B = 16'h00B8; #100;
A = 16'h008E; B = 16'h00B9; #100;
A = 16'h008E; B = 16'h00BA; #100;
A = 16'h008E; B = 16'h00BB; #100;
A = 16'h008E; B = 16'h00BC; #100;
A = 16'h008E; B = 16'h00BD; #100;
A = 16'h008E; B = 16'h00BE; #100;
A = 16'h008E; B = 16'h00BF; #100;
A = 16'h008E; B = 16'h00C0; #100;
A = 16'h008E; B = 16'h00C1; #100;
A = 16'h008E; B = 16'h00C2; #100;
A = 16'h008E; B = 16'h00C3; #100;
A = 16'h008E; B = 16'h00C4; #100;
A = 16'h008E; B = 16'h00C5; #100;
A = 16'h008E; B = 16'h00C6; #100;
A = 16'h008E; B = 16'h00C7; #100;
A = 16'h008E; B = 16'h00C8; #100;
A = 16'h008E; B = 16'h00C9; #100;
A = 16'h008E; B = 16'h00CA; #100;
A = 16'h008E; B = 16'h00CB; #100;
A = 16'h008E; B = 16'h00CC; #100;
A = 16'h008E; B = 16'h00CD; #100;
A = 16'h008E; B = 16'h00CE; #100;
A = 16'h008E; B = 16'h00CF; #100;
A = 16'h008E; B = 16'h00D0; #100;
A = 16'h008E; B = 16'h00D1; #100;
A = 16'h008E; B = 16'h00D2; #100;
A = 16'h008E; B = 16'h00D3; #100;
A = 16'h008E; B = 16'h00D4; #100;
A = 16'h008E; B = 16'h00D5; #100;
A = 16'h008E; B = 16'h00D6; #100;
A = 16'h008E; B = 16'h00D7; #100;
A = 16'h008E; B = 16'h00D8; #100;
A = 16'h008E; B = 16'h00D9; #100;
A = 16'h008E; B = 16'h00DA; #100;
A = 16'h008E; B = 16'h00DB; #100;
A = 16'h008E; B = 16'h00DC; #100;
A = 16'h008E; B = 16'h00DD; #100;
A = 16'h008E; B = 16'h00DE; #100;
A = 16'h008E; B = 16'h00DF; #100;
A = 16'h008E; B = 16'h00E0; #100;
A = 16'h008E; B = 16'h00E1; #100;
A = 16'h008E; B = 16'h00E2; #100;
A = 16'h008E; B = 16'h00E3; #100;
A = 16'h008E; B = 16'h00E4; #100;
A = 16'h008E; B = 16'h00E5; #100;
A = 16'h008E; B = 16'h00E6; #100;
A = 16'h008E; B = 16'h00E7; #100;
A = 16'h008E; B = 16'h00E8; #100;
A = 16'h008E; B = 16'h00E9; #100;
A = 16'h008E; B = 16'h00EA; #100;
A = 16'h008E; B = 16'h00EB; #100;
A = 16'h008E; B = 16'h00EC; #100;
A = 16'h008E; B = 16'h00ED; #100;
A = 16'h008E; B = 16'h00EE; #100;
A = 16'h008E; B = 16'h00EF; #100;
A = 16'h008E; B = 16'h00F0; #100;
A = 16'h008E; B = 16'h00F1; #100;
A = 16'h008E; B = 16'h00F2; #100;
A = 16'h008E; B = 16'h00F3; #100;
A = 16'h008E; B = 16'h00F4; #100;
A = 16'h008E; B = 16'h00F5; #100;
A = 16'h008E; B = 16'h00F6; #100;
A = 16'h008E; B = 16'h00F7; #100;
A = 16'h008E; B = 16'h00F8; #100;
A = 16'h008E; B = 16'h00F9; #100;
A = 16'h008E; B = 16'h00FA; #100;
A = 16'h008E; B = 16'h00FB; #100;
A = 16'h008E; B = 16'h00FC; #100;
A = 16'h008E; B = 16'h00FD; #100;
A = 16'h008E; B = 16'h00FE; #100;
A = 16'h008E; B = 16'h00FF; #100;
A = 16'h008F; B = 16'h000; #100;
A = 16'h008F; B = 16'h001; #100;
A = 16'h008F; B = 16'h002; #100;
A = 16'h008F; B = 16'h003; #100;
A = 16'h008F; B = 16'h004; #100;
A = 16'h008F; B = 16'h005; #100;
A = 16'h008F; B = 16'h006; #100;
A = 16'h008F; B = 16'h007; #100;
A = 16'h008F; B = 16'h008; #100;
A = 16'h008F; B = 16'h009; #100;
A = 16'h008F; B = 16'h00A; #100;
A = 16'h008F; B = 16'h00B; #100;
A = 16'h008F; B = 16'h00C; #100;
A = 16'h008F; B = 16'h00D; #100;
A = 16'h008F; B = 16'h00E; #100;
A = 16'h008F; B = 16'h00F; #100;
A = 16'h008F; B = 16'h0010; #100;
A = 16'h008F; B = 16'h0011; #100;
A = 16'h008F; B = 16'h0012; #100;
A = 16'h008F; B = 16'h0013; #100;
A = 16'h008F; B = 16'h0014; #100;
A = 16'h008F; B = 16'h0015; #100;
A = 16'h008F; B = 16'h0016; #100;
A = 16'h008F; B = 16'h0017; #100;
A = 16'h008F; B = 16'h0018; #100;
A = 16'h008F; B = 16'h0019; #100;
A = 16'h008F; B = 16'h001A; #100;
A = 16'h008F; B = 16'h001B; #100;
A = 16'h008F; B = 16'h001C; #100;
A = 16'h008F; B = 16'h001D; #100;
A = 16'h008F; B = 16'h001E; #100;
A = 16'h008F; B = 16'h001F; #100;
A = 16'h008F; B = 16'h0020; #100;
A = 16'h008F; B = 16'h0021; #100;
A = 16'h008F; B = 16'h0022; #100;
A = 16'h008F; B = 16'h0023; #100;
A = 16'h008F; B = 16'h0024; #100;
A = 16'h008F; B = 16'h0025; #100;
A = 16'h008F; B = 16'h0026; #100;
A = 16'h008F; B = 16'h0027; #100;
A = 16'h008F; B = 16'h0028; #100;
A = 16'h008F; B = 16'h0029; #100;
A = 16'h008F; B = 16'h002A; #100;
A = 16'h008F; B = 16'h002B; #100;
A = 16'h008F; B = 16'h002C; #100;
A = 16'h008F; B = 16'h002D; #100;
A = 16'h008F; B = 16'h002E; #100;
A = 16'h008F; B = 16'h002F; #100;
A = 16'h008F; B = 16'h0030; #100;
A = 16'h008F; B = 16'h0031; #100;
A = 16'h008F; B = 16'h0032; #100;
A = 16'h008F; B = 16'h0033; #100;
A = 16'h008F; B = 16'h0034; #100;
A = 16'h008F; B = 16'h0035; #100;
A = 16'h008F; B = 16'h0036; #100;
A = 16'h008F; B = 16'h0037; #100;
A = 16'h008F; B = 16'h0038; #100;
A = 16'h008F; B = 16'h0039; #100;
A = 16'h008F; B = 16'h003A; #100;
A = 16'h008F; B = 16'h003B; #100;
A = 16'h008F; B = 16'h003C; #100;
A = 16'h008F; B = 16'h003D; #100;
A = 16'h008F; B = 16'h003E; #100;
A = 16'h008F; B = 16'h003F; #100;
A = 16'h008F; B = 16'h0040; #100;
A = 16'h008F; B = 16'h0041; #100;
A = 16'h008F; B = 16'h0042; #100;
A = 16'h008F; B = 16'h0043; #100;
A = 16'h008F; B = 16'h0044; #100;
A = 16'h008F; B = 16'h0045; #100;
A = 16'h008F; B = 16'h0046; #100;
A = 16'h008F; B = 16'h0047; #100;
A = 16'h008F; B = 16'h0048; #100;
A = 16'h008F; B = 16'h0049; #100;
A = 16'h008F; B = 16'h004A; #100;
A = 16'h008F; B = 16'h004B; #100;
A = 16'h008F; B = 16'h004C; #100;
A = 16'h008F; B = 16'h004D; #100;
A = 16'h008F; B = 16'h004E; #100;
A = 16'h008F; B = 16'h004F; #100;
A = 16'h008F; B = 16'h0050; #100;
A = 16'h008F; B = 16'h0051; #100;
A = 16'h008F; B = 16'h0052; #100;
A = 16'h008F; B = 16'h0053; #100;
A = 16'h008F; B = 16'h0054; #100;
A = 16'h008F; B = 16'h0055; #100;
A = 16'h008F; B = 16'h0056; #100;
A = 16'h008F; B = 16'h0057; #100;
A = 16'h008F; B = 16'h0058; #100;
A = 16'h008F; B = 16'h0059; #100;
A = 16'h008F; B = 16'h005A; #100;
A = 16'h008F; B = 16'h005B; #100;
A = 16'h008F; B = 16'h005C; #100;
A = 16'h008F; B = 16'h005D; #100;
A = 16'h008F; B = 16'h005E; #100;
A = 16'h008F; B = 16'h005F; #100;
A = 16'h008F; B = 16'h0060; #100;
A = 16'h008F; B = 16'h0061; #100;
A = 16'h008F; B = 16'h0062; #100;
A = 16'h008F; B = 16'h0063; #100;
A = 16'h008F; B = 16'h0064; #100;
A = 16'h008F; B = 16'h0065; #100;
A = 16'h008F; B = 16'h0066; #100;
A = 16'h008F; B = 16'h0067; #100;
A = 16'h008F; B = 16'h0068; #100;
A = 16'h008F; B = 16'h0069; #100;
A = 16'h008F; B = 16'h006A; #100;
A = 16'h008F; B = 16'h006B; #100;
A = 16'h008F; B = 16'h006C; #100;
A = 16'h008F; B = 16'h006D; #100;
A = 16'h008F; B = 16'h006E; #100;
A = 16'h008F; B = 16'h006F; #100;
A = 16'h008F; B = 16'h0070; #100;
A = 16'h008F; B = 16'h0071; #100;
A = 16'h008F; B = 16'h0072; #100;
A = 16'h008F; B = 16'h0073; #100;
A = 16'h008F; B = 16'h0074; #100;
A = 16'h008F; B = 16'h0075; #100;
A = 16'h008F; B = 16'h0076; #100;
A = 16'h008F; B = 16'h0077; #100;
A = 16'h008F; B = 16'h0078; #100;
A = 16'h008F; B = 16'h0079; #100;
A = 16'h008F; B = 16'h007A; #100;
A = 16'h008F; B = 16'h007B; #100;
A = 16'h008F; B = 16'h007C; #100;
A = 16'h008F; B = 16'h007D; #100;
A = 16'h008F; B = 16'h007E; #100;
A = 16'h008F; B = 16'h007F; #100;
A = 16'h008F; B = 16'h0080; #100;
A = 16'h008F; B = 16'h0081; #100;
A = 16'h008F; B = 16'h0082; #100;
A = 16'h008F; B = 16'h0083; #100;
A = 16'h008F; B = 16'h0084; #100;
A = 16'h008F; B = 16'h0085; #100;
A = 16'h008F; B = 16'h0086; #100;
A = 16'h008F; B = 16'h0087; #100;
A = 16'h008F; B = 16'h0088; #100;
A = 16'h008F; B = 16'h0089; #100;
A = 16'h008F; B = 16'h008A; #100;
A = 16'h008F; B = 16'h008B; #100;
A = 16'h008F; B = 16'h008C; #100;
A = 16'h008F; B = 16'h008D; #100;
A = 16'h008F; B = 16'h008E; #100;
A = 16'h008F; B = 16'h008F; #100;
A = 16'h008F; B = 16'h0090; #100;
A = 16'h008F; B = 16'h0091; #100;
A = 16'h008F; B = 16'h0092; #100;
A = 16'h008F; B = 16'h0093; #100;
A = 16'h008F; B = 16'h0094; #100;
A = 16'h008F; B = 16'h0095; #100;
A = 16'h008F; B = 16'h0096; #100;
A = 16'h008F; B = 16'h0097; #100;
A = 16'h008F; B = 16'h0098; #100;
A = 16'h008F; B = 16'h0099; #100;
A = 16'h008F; B = 16'h009A; #100;
A = 16'h008F; B = 16'h009B; #100;
A = 16'h008F; B = 16'h009C; #100;
A = 16'h008F; B = 16'h009D; #100;
A = 16'h008F; B = 16'h009E; #100;
A = 16'h008F; B = 16'h009F; #100;
A = 16'h008F; B = 16'h00A0; #100;
A = 16'h008F; B = 16'h00A1; #100;
A = 16'h008F; B = 16'h00A2; #100;
A = 16'h008F; B = 16'h00A3; #100;
A = 16'h008F; B = 16'h00A4; #100;
A = 16'h008F; B = 16'h00A5; #100;
A = 16'h008F; B = 16'h00A6; #100;
A = 16'h008F; B = 16'h00A7; #100;
A = 16'h008F; B = 16'h00A8; #100;
A = 16'h008F; B = 16'h00A9; #100;
A = 16'h008F; B = 16'h00AA; #100;
A = 16'h008F; B = 16'h00AB; #100;
A = 16'h008F; B = 16'h00AC; #100;
A = 16'h008F; B = 16'h00AD; #100;
A = 16'h008F; B = 16'h00AE; #100;
A = 16'h008F; B = 16'h00AF; #100;
A = 16'h008F; B = 16'h00B0; #100;
A = 16'h008F; B = 16'h00B1; #100;
A = 16'h008F; B = 16'h00B2; #100;
A = 16'h008F; B = 16'h00B3; #100;
A = 16'h008F; B = 16'h00B4; #100;
A = 16'h008F; B = 16'h00B5; #100;
A = 16'h008F; B = 16'h00B6; #100;
A = 16'h008F; B = 16'h00B7; #100;
A = 16'h008F; B = 16'h00B8; #100;
A = 16'h008F; B = 16'h00B9; #100;
A = 16'h008F; B = 16'h00BA; #100;
A = 16'h008F; B = 16'h00BB; #100;
A = 16'h008F; B = 16'h00BC; #100;
A = 16'h008F; B = 16'h00BD; #100;
A = 16'h008F; B = 16'h00BE; #100;
A = 16'h008F; B = 16'h00BF; #100;
A = 16'h008F; B = 16'h00C0; #100;
A = 16'h008F; B = 16'h00C1; #100;
A = 16'h008F; B = 16'h00C2; #100;
A = 16'h008F; B = 16'h00C3; #100;
A = 16'h008F; B = 16'h00C4; #100;
A = 16'h008F; B = 16'h00C5; #100;
A = 16'h008F; B = 16'h00C6; #100;
A = 16'h008F; B = 16'h00C7; #100;
A = 16'h008F; B = 16'h00C8; #100;
A = 16'h008F; B = 16'h00C9; #100;
A = 16'h008F; B = 16'h00CA; #100;
A = 16'h008F; B = 16'h00CB; #100;
A = 16'h008F; B = 16'h00CC; #100;
A = 16'h008F; B = 16'h00CD; #100;
A = 16'h008F; B = 16'h00CE; #100;
A = 16'h008F; B = 16'h00CF; #100;
A = 16'h008F; B = 16'h00D0; #100;
A = 16'h008F; B = 16'h00D1; #100;
A = 16'h008F; B = 16'h00D2; #100;
A = 16'h008F; B = 16'h00D3; #100;
A = 16'h008F; B = 16'h00D4; #100;
A = 16'h008F; B = 16'h00D5; #100;
A = 16'h008F; B = 16'h00D6; #100;
A = 16'h008F; B = 16'h00D7; #100;
A = 16'h008F; B = 16'h00D8; #100;
A = 16'h008F; B = 16'h00D9; #100;
A = 16'h008F; B = 16'h00DA; #100;
A = 16'h008F; B = 16'h00DB; #100;
A = 16'h008F; B = 16'h00DC; #100;
A = 16'h008F; B = 16'h00DD; #100;
A = 16'h008F; B = 16'h00DE; #100;
A = 16'h008F; B = 16'h00DF; #100;
A = 16'h008F; B = 16'h00E0; #100;
A = 16'h008F; B = 16'h00E1; #100;
A = 16'h008F; B = 16'h00E2; #100;
A = 16'h008F; B = 16'h00E3; #100;
A = 16'h008F; B = 16'h00E4; #100;
A = 16'h008F; B = 16'h00E5; #100;
A = 16'h008F; B = 16'h00E6; #100;
A = 16'h008F; B = 16'h00E7; #100;
A = 16'h008F; B = 16'h00E8; #100;
A = 16'h008F; B = 16'h00E9; #100;
A = 16'h008F; B = 16'h00EA; #100;
A = 16'h008F; B = 16'h00EB; #100;
A = 16'h008F; B = 16'h00EC; #100;
A = 16'h008F; B = 16'h00ED; #100;
A = 16'h008F; B = 16'h00EE; #100;
A = 16'h008F; B = 16'h00EF; #100;
A = 16'h008F; B = 16'h00F0; #100;
A = 16'h008F; B = 16'h00F1; #100;
A = 16'h008F; B = 16'h00F2; #100;
A = 16'h008F; B = 16'h00F3; #100;
A = 16'h008F; B = 16'h00F4; #100;
A = 16'h008F; B = 16'h00F5; #100;
A = 16'h008F; B = 16'h00F6; #100;
A = 16'h008F; B = 16'h00F7; #100;
A = 16'h008F; B = 16'h00F8; #100;
A = 16'h008F; B = 16'h00F9; #100;
A = 16'h008F; B = 16'h00FA; #100;
A = 16'h008F; B = 16'h00FB; #100;
A = 16'h008F; B = 16'h00FC; #100;
A = 16'h008F; B = 16'h00FD; #100;
A = 16'h008F; B = 16'h00FE; #100;
A = 16'h008F; B = 16'h00FF; #100;
A = 16'h0090; B = 16'h000; #100;
A = 16'h0090; B = 16'h001; #100;
A = 16'h0090; B = 16'h002; #100;
A = 16'h0090; B = 16'h003; #100;
A = 16'h0090; B = 16'h004; #100;
A = 16'h0090; B = 16'h005; #100;
A = 16'h0090; B = 16'h006; #100;
A = 16'h0090; B = 16'h007; #100;
A = 16'h0090; B = 16'h008; #100;
A = 16'h0090; B = 16'h009; #100;
A = 16'h0090; B = 16'h00A; #100;
A = 16'h0090; B = 16'h00B; #100;
A = 16'h0090; B = 16'h00C; #100;
A = 16'h0090; B = 16'h00D; #100;
A = 16'h0090; B = 16'h00E; #100;
A = 16'h0090; B = 16'h00F; #100;
A = 16'h0090; B = 16'h0010; #100;
A = 16'h0090; B = 16'h0011; #100;
A = 16'h0090; B = 16'h0012; #100;
A = 16'h0090; B = 16'h0013; #100;
A = 16'h0090; B = 16'h0014; #100;
A = 16'h0090; B = 16'h0015; #100;
A = 16'h0090; B = 16'h0016; #100;
A = 16'h0090; B = 16'h0017; #100;
A = 16'h0090; B = 16'h0018; #100;
A = 16'h0090; B = 16'h0019; #100;
A = 16'h0090; B = 16'h001A; #100;
A = 16'h0090; B = 16'h001B; #100;
A = 16'h0090; B = 16'h001C; #100;
A = 16'h0090; B = 16'h001D; #100;
A = 16'h0090; B = 16'h001E; #100;
A = 16'h0090; B = 16'h001F; #100;
A = 16'h0090; B = 16'h0020; #100;
A = 16'h0090; B = 16'h0021; #100;
A = 16'h0090; B = 16'h0022; #100;
A = 16'h0090; B = 16'h0023; #100;
A = 16'h0090; B = 16'h0024; #100;
A = 16'h0090; B = 16'h0025; #100;
A = 16'h0090; B = 16'h0026; #100;
A = 16'h0090; B = 16'h0027; #100;
A = 16'h0090; B = 16'h0028; #100;
A = 16'h0090; B = 16'h0029; #100;
A = 16'h0090; B = 16'h002A; #100;
A = 16'h0090; B = 16'h002B; #100;
A = 16'h0090; B = 16'h002C; #100;
A = 16'h0090; B = 16'h002D; #100;
A = 16'h0090; B = 16'h002E; #100;
A = 16'h0090; B = 16'h002F; #100;
A = 16'h0090; B = 16'h0030; #100;
A = 16'h0090; B = 16'h0031; #100;
A = 16'h0090; B = 16'h0032; #100;
A = 16'h0090; B = 16'h0033; #100;
A = 16'h0090; B = 16'h0034; #100;
A = 16'h0090; B = 16'h0035; #100;
A = 16'h0090; B = 16'h0036; #100;
A = 16'h0090; B = 16'h0037; #100;
A = 16'h0090; B = 16'h0038; #100;
A = 16'h0090; B = 16'h0039; #100;
A = 16'h0090; B = 16'h003A; #100;
A = 16'h0090; B = 16'h003B; #100;
A = 16'h0090; B = 16'h003C; #100;
A = 16'h0090; B = 16'h003D; #100;
A = 16'h0090; B = 16'h003E; #100;
A = 16'h0090; B = 16'h003F; #100;
A = 16'h0090; B = 16'h0040; #100;
A = 16'h0090; B = 16'h0041; #100;
A = 16'h0090; B = 16'h0042; #100;
A = 16'h0090; B = 16'h0043; #100;
A = 16'h0090; B = 16'h0044; #100;
A = 16'h0090; B = 16'h0045; #100;
A = 16'h0090; B = 16'h0046; #100;
A = 16'h0090; B = 16'h0047; #100;
A = 16'h0090; B = 16'h0048; #100;
A = 16'h0090; B = 16'h0049; #100;
A = 16'h0090; B = 16'h004A; #100;
A = 16'h0090; B = 16'h004B; #100;
A = 16'h0090; B = 16'h004C; #100;
A = 16'h0090; B = 16'h004D; #100;
A = 16'h0090; B = 16'h004E; #100;
A = 16'h0090; B = 16'h004F; #100;
A = 16'h0090; B = 16'h0050; #100;
A = 16'h0090; B = 16'h0051; #100;
A = 16'h0090; B = 16'h0052; #100;
A = 16'h0090; B = 16'h0053; #100;
A = 16'h0090; B = 16'h0054; #100;
A = 16'h0090; B = 16'h0055; #100;
A = 16'h0090; B = 16'h0056; #100;
A = 16'h0090; B = 16'h0057; #100;
A = 16'h0090; B = 16'h0058; #100;
A = 16'h0090; B = 16'h0059; #100;
A = 16'h0090; B = 16'h005A; #100;
A = 16'h0090; B = 16'h005B; #100;
A = 16'h0090; B = 16'h005C; #100;
A = 16'h0090; B = 16'h005D; #100;
A = 16'h0090; B = 16'h005E; #100;
A = 16'h0090; B = 16'h005F; #100;
A = 16'h0090; B = 16'h0060; #100;
A = 16'h0090; B = 16'h0061; #100;
A = 16'h0090; B = 16'h0062; #100;
A = 16'h0090; B = 16'h0063; #100;
A = 16'h0090; B = 16'h0064; #100;
A = 16'h0090; B = 16'h0065; #100;
A = 16'h0090; B = 16'h0066; #100;
A = 16'h0090; B = 16'h0067; #100;
A = 16'h0090; B = 16'h0068; #100;
A = 16'h0090; B = 16'h0069; #100;
A = 16'h0090; B = 16'h006A; #100;
A = 16'h0090; B = 16'h006B; #100;
A = 16'h0090; B = 16'h006C; #100;
A = 16'h0090; B = 16'h006D; #100;
A = 16'h0090; B = 16'h006E; #100;
A = 16'h0090; B = 16'h006F; #100;
A = 16'h0090; B = 16'h0070; #100;
A = 16'h0090; B = 16'h0071; #100;
A = 16'h0090; B = 16'h0072; #100;
A = 16'h0090; B = 16'h0073; #100;
A = 16'h0090; B = 16'h0074; #100;
A = 16'h0090; B = 16'h0075; #100;
A = 16'h0090; B = 16'h0076; #100;
A = 16'h0090; B = 16'h0077; #100;
A = 16'h0090; B = 16'h0078; #100;
A = 16'h0090; B = 16'h0079; #100;
A = 16'h0090; B = 16'h007A; #100;
A = 16'h0090; B = 16'h007B; #100;
A = 16'h0090; B = 16'h007C; #100;
A = 16'h0090; B = 16'h007D; #100;
A = 16'h0090; B = 16'h007E; #100;
A = 16'h0090; B = 16'h007F; #100;
A = 16'h0090; B = 16'h0080; #100;
A = 16'h0090; B = 16'h0081; #100;
A = 16'h0090; B = 16'h0082; #100;
A = 16'h0090; B = 16'h0083; #100;
A = 16'h0090; B = 16'h0084; #100;
A = 16'h0090; B = 16'h0085; #100;
A = 16'h0090; B = 16'h0086; #100;
A = 16'h0090; B = 16'h0087; #100;
A = 16'h0090; B = 16'h0088; #100;
A = 16'h0090; B = 16'h0089; #100;
A = 16'h0090; B = 16'h008A; #100;
A = 16'h0090; B = 16'h008B; #100;
A = 16'h0090; B = 16'h008C; #100;
A = 16'h0090; B = 16'h008D; #100;
A = 16'h0090; B = 16'h008E; #100;
A = 16'h0090; B = 16'h008F; #100;
A = 16'h0090; B = 16'h0090; #100;
A = 16'h0090; B = 16'h0091; #100;
A = 16'h0090; B = 16'h0092; #100;
A = 16'h0090; B = 16'h0093; #100;
A = 16'h0090; B = 16'h0094; #100;
A = 16'h0090; B = 16'h0095; #100;
A = 16'h0090; B = 16'h0096; #100;
A = 16'h0090; B = 16'h0097; #100;
A = 16'h0090; B = 16'h0098; #100;
A = 16'h0090; B = 16'h0099; #100;
A = 16'h0090; B = 16'h009A; #100;
A = 16'h0090; B = 16'h009B; #100;
A = 16'h0090; B = 16'h009C; #100;
A = 16'h0090; B = 16'h009D; #100;
A = 16'h0090; B = 16'h009E; #100;
A = 16'h0090; B = 16'h009F; #100;
A = 16'h0090; B = 16'h00A0; #100;
A = 16'h0090; B = 16'h00A1; #100;
A = 16'h0090; B = 16'h00A2; #100;
A = 16'h0090; B = 16'h00A3; #100;
A = 16'h0090; B = 16'h00A4; #100;
A = 16'h0090; B = 16'h00A5; #100;
A = 16'h0090; B = 16'h00A6; #100;
A = 16'h0090; B = 16'h00A7; #100;
A = 16'h0090; B = 16'h00A8; #100;
A = 16'h0090; B = 16'h00A9; #100;
A = 16'h0090; B = 16'h00AA; #100;
A = 16'h0090; B = 16'h00AB; #100;
A = 16'h0090; B = 16'h00AC; #100;
A = 16'h0090; B = 16'h00AD; #100;
A = 16'h0090; B = 16'h00AE; #100;
A = 16'h0090; B = 16'h00AF; #100;
A = 16'h0090; B = 16'h00B0; #100;
A = 16'h0090; B = 16'h00B1; #100;
A = 16'h0090; B = 16'h00B2; #100;
A = 16'h0090; B = 16'h00B3; #100;
A = 16'h0090; B = 16'h00B4; #100;
A = 16'h0090; B = 16'h00B5; #100;
A = 16'h0090; B = 16'h00B6; #100;
A = 16'h0090; B = 16'h00B7; #100;
A = 16'h0090; B = 16'h00B8; #100;
A = 16'h0090; B = 16'h00B9; #100;
A = 16'h0090; B = 16'h00BA; #100;
A = 16'h0090; B = 16'h00BB; #100;
A = 16'h0090; B = 16'h00BC; #100;
A = 16'h0090; B = 16'h00BD; #100;
A = 16'h0090; B = 16'h00BE; #100;
A = 16'h0090; B = 16'h00BF; #100;
A = 16'h0090; B = 16'h00C0; #100;
A = 16'h0090; B = 16'h00C1; #100;
A = 16'h0090; B = 16'h00C2; #100;
A = 16'h0090; B = 16'h00C3; #100;
A = 16'h0090; B = 16'h00C4; #100;
A = 16'h0090; B = 16'h00C5; #100;
A = 16'h0090; B = 16'h00C6; #100;
A = 16'h0090; B = 16'h00C7; #100;
A = 16'h0090; B = 16'h00C8; #100;
A = 16'h0090; B = 16'h00C9; #100;
A = 16'h0090; B = 16'h00CA; #100;
A = 16'h0090; B = 16'h00CB; #100;
A = 16'h0090; B = 16'h00CC; #100;
A = 16'h0090; B = 16'h00CD; #100;
A = 16'h0090; B = 16'h00CE; #100;
A = 16'h0090; B = 16'h00CF; #100;
A = 16'h0090; B = 16'h00D0; #100;
A = 16'h0090; B = 16'h00D1; #100;
A = 16'h0090; B = 16'h00D2; #100;
A = 16'h0090; B = 16'h00D3; #100;
A = 16'h0090; B = 16'h00D4; #100;
A = 16'h0090; B = 16'h00D5; #100;
A = 16'h0090; B = 16'h00D6; #100;
A = 16'h0090; B = 16'h00D7; #100;
A = 16'h0090; B = 16'h00D8; #100;
A = 16'h0090; B = 16'h00D9; #100;
A = 16'h0090; B = 16'h00DA; #100;
A = 16'h0090; B = 16'h00DB; #100;
A = 16'h0090; B = 16'h00DC; #100;
A = 16'h0090; B = 16'h00DD; #100;
A = 16'h0090; B = 16'h00DE; #100;
A = 16'h0090; B = 16'h00DF; #100;
A = 16'h0090; B = 16'h00E0; #100;
A = 16'h0090; B = 16'h00E1; #100;
A = 16'h0090; B = 16'h00E2; #100;
A = 16'h0090; B = 16'h00E3; #100;
A = 16'h0090; B = 16'h00E4; #100;
A = 16'h0090; B = 16'h00E5; #100;
A = 16'h0090; B = 16'h00E6; #100;
A = 16'h0090; B = 16'h00E7; #100;
A = 16'h0090; B = 16'h00E8; #100;
A = 16'h0090; B = 16'h00E9; #100;
A = 16'h0090; B = 16'h00EA; #100;
A = 16'h0090; B = 16'h00EB; #100;
A = 16'h0090; B = 16'h00EC; #100;
A = 16'h0090; B = 16'h00ED; #100;
A = 16'h0090; B = 16'h00EE; #100;
A = 16'h0090; B = 16'h00EF; #100;
A = 16'h0090; B = 16'h00F0; #100;
A = 16'h0090; B = 16'h00F1; #100;
A = 16'h0090; B = 16'h00F2; #100;
A = 16'h0090; B = 16'h00F3; #100;
A = 16'h0090; B = 16'h00F4; #100;
A = 16'h0090; B = 16'h00F5; #100;
A = 16'h0090; B = 16'h00F6; #100;
A = 16'h0090; B = 16'h00F7; #100;
A = 16'h0090; B = 16'h00F8; #100;
A = 16'h0090; B = 16'h00F9; #100;
A = 16'h0090; B = 16'h00FA; #100;
A = 16'h0090; B = 16'h00FB; #100;
A = 16'h0090; B = 16'h00FC; #100;
A = 16'h0090; B = 16'h00FD; #100;
A = 16'h0090; B = 16'h00FE; #100;
A = 16'h0090; B = 16'h00FF; #100;
A = 16'h0091; B = 16'h000; #100;
A = 16'h0091; B = 16'h001; #100;
A = 16'h0091; B = 16'h002; #100;
A = 16'h0091; B = 16'h003; #100;
A = 16'h0091; B = 16'h004; #100;
A = 16'h0091; B = 16'h005; #100;
A = 16'h0091; B = 16'h006; #100;
A = 16'h0091; B = 16'h007; #100;
A = 16'h0091; B = 16'h008; #100;
A = 16'h0091; B = 16'h009; #100;
A = 16'h0091; B = 16'h00A; #100;
A = 16'h0091; B = 16'h00B; #100;
A = 16'h0091; B = 16'h00C; #100;
A = 16'h0091; B = 16'h00D; #100;
A = 16'h0091; B = 16'h00E; #100;
A = 16'h0091; B = 16'h00F; #100;
A = 16'h0091; B = 16'h0010; #100;
A = 16'h0091; B = 16'h0011; #100;
A = 16'h0091; B = 16'h0012; #100;
A = 16'h0091; B = 16'h0013; #100;
A = 16'h0091; B = 16'h0014; #100;
A = 16'h0091; B = 16'h0015; #100;
A = 16'h0091; B = 16'h0016; #100;
A = 16'h0091; B = 16'h0017; #100;
A = 16'h0091; B = 16'h0018; #100;
A = 16'h0091; B = 16'h0019; #100;
A = 16'h0091; B = 16'h001A; #100;
A = 16'h0091; B = 16'h001B; #100;
A = 16'h0091; B = 16'h001C; #100;
A = 16'h0091; B = 16'h001D; #100;
A = 16'h0091; B = 16'h001E; #100;
A = 16'h0091; B = 16'h001F; #100;
A = 16'h0091; B = 16'h0020; #100;
A = 16'h0091; B = 16'h0021; #100;
A = 16'h0091; B = 16'h0022; #100;
A = 16'h0091; B = 16'h0023; #100;
A = 16'h0091; B = 16'h0024; #100;
A = 16'h0091; B = 16'h0025; #100;
A = 16'h0091; B = 16'h0026; #100;
A = 16'h0091; B = 16'h0027; #100;
A = 16'h0091; B = 16'h0028; #100;
A = 16'h0091; B = 16'h0029; #100;
A = 16'h0091; B = 16'h002A; #100;
A = 16'h0091; B = 16'h002B; #100;
A = 16'h0091; B = 16'h002C; #100;
A = 16'h0091; B = 16'h002D; #100;
A = 16'h0091; B = 16'h002E; #100;
A = 16'h0091; B = 16'h002F; #100;
A = 16'h0091; B = 16'h0030; #100;
A = 16'h0091; B = 16'h0031; #100;
A = 16'h0091; B = 16'h0032; #100;
A = 16'h0091; B = 16'h0033; #100;
A = 16'h0091; B = 16'h0034; #100;
A = 16'h0091; B = 16'h0035; #100;
A = 16'h0091; B = 16'h0036; #100;
A = 16'h0091; B = 16'h0037; #100;
A = 16'h0091; B = 16'h0038; #100;
A = 16'h0091; B = 16'h0039; #100;
A = 16'h0091; B = 16'h003A; #100;
A = 16'h0091; B = 16'h003B; #100;
A = 16'h0091; B = 16'h003C; #100;
A = 16'h0091; B = 16'h003D; #100;
A = 16'h0091; B = 16'h003E; #100;
A = 16'h0091; B = 16'h003F; #100;
A = 16'h0091; B = 16'h0040; #100;
A = 16'h0091; B = 16'h0041; #100;
A = 16'h0091; B = 16'h0042; #100;
A = 16'h0091; B = 16'h0043; #100;
A = 16'h0091; B = 16'h0044; #100;
A = 16'h0091; B = 16'h0045; #100;
A = 16'h0091; B = 16'h0046; #100;
A = 16'h0091; B = 16'h0047; #100;
A = 16'h0091; B = 16'h0048; #100;
A = 16'h0091; B = 16'h0049; #100;
A = 16'h0091; B = 16'h004A; #100;
A = 16'h0091; B = 16'h004B; #100;
A = 16'h0091; B = 16'h004C; #100;
A = 16'h0091; B = 16'h004D; #100;
A = 16'h0091; B = 16'h004E; #100;
A = 16'h0091; B = 16'h004F; #100;
A = 16'h0091; B = 16'h0050; #100;
A = 16'h0091; B = 16'h0051; #100;
A = 16'h0091; B = 16'h0052; #100;
A = 16'h0091; B = 16'h0053; #100;
A = 16'h0091; B = 16'h0054; #100;
A = 16'h0091; B = 16'h0055; #100;
A = 16'h0091; B = 16'h0056; #100;
A = 16'h0091; B = 16'h0057; #100;
A = 16'h0091; B = 16'h0058; #100;
A = 16'h0091; B = 16'h0059; #100;
A = 16'h0091; B = 16'h005A; #100;
A = 16'h0091; B = 16'h005B; #100;
A = 16'h0091; B = 16'h005C; #100;
A = 16'h0091; B = 16'h005D; #100;
A = 16'h0091; B = 16'h005E; #100;
A = 16'h0091; B = 16'h005F; #100;
A = 16'h0091; B = 16'h0060; #100;
A = 16'h0091; B = 16'h0061; #100;
A = 16'h0091; B = 16'h0062; #100;
A = 16'h0091; B = 16'h0063; #100;
A = 16'h0091; B = 16'h0064; #100;
A = 16'h0091; B = 16'h0065; #100;
A = 16'h0091; B = 16'h0066; #100;
A = 16'h0091; B = 16'h0067; #100;
A = 16'h0091; B = 16'h0068; #100;
A = 16'h0091; B = 16'h0069; #100;
A = 16'h0091; B = 16'h006A; #100;
A = 16'h0091; B = 16'h006B; #100;
A = 16'h0091; B = 16'h006C; #100;
A = 16'h0091; B = 16'h006D; #100;
A = 16'h0091; B = 16'h006E; #100;
A = 16'h0091; B = 16'h006F; #100;
A = 16'h0091; B = 16'h0070; #100;
A = 16'h0091; B = 16'h0071; #100;
A = 16'h0091; B = 16'h0072; #100;
A = 16'h0091; B = 16'h0073; #100;
A = 16'h0091; B = 16'h0074; #100;
A = 16'h0091; B = 16'h0075; #100;
A = 16'h0091; B = 16'h0076; #100;
A = 16'h0091; B = 16'h0077; #100;
A = 16'h0091; B = 16'h0078; #100;
A = 16'h0091; B = 16'h0079; #100;
A = 16'h0091; B = 16'h007A; #100;
A = 16'h0091; B = 16'h007B; #100;
A = 16'h0091; B = 16'h007C; #100;
A = 16'h0091; B = 16'h007D; #100;
A = 16'h0091; B = 16'h007E; #100;
A = 16'h0091; B = 16'h007F; #100;
A = 16'h0091; B = 16'h0080; #100;
A = 16'h0091; B = 16'h0081; #100;
A = 16'h0091; B = 16'h0082; #100;
A = 16'h0091; B = 16'h0083; #100;
A = 16'h0091; B = 16'h0084; #100;
A = 16'h0091; B = 16'h0085; #100;
A = 16'h0091; B = 16'h0086; #100;
A = 16'h0091; B = 16'h0087; #100;
A = 16'h0091; B = 16'h0088; #100;
A = 16'h0091; B = 16'h0089; #100;
A = 16'h0091; B = 16'h008A; #100;
A = 16'h0091; B = 16'h008B; #100;
A = 16'h0091; B = 16'h008C; #100;
A = 16'h0091; B = 16'h008D; #100;
A = 16'h0091; B = 16'h008E; #100;
A = 16'h0091; B = 16'h008F; #100;
A = 16'h0091; B = 16'h0090; #100;
A = 16'h0091; B = 16'h0091; #100;
A = 16'h0091; B = 16'h0092; #100;
A = 16'h0091; B = 16'h0093; #100;
A = 16'h0091; B = 16'h0094; #100;
A = 16'h0091; B = 16'h0095; #100;
A = 16'h0091; B = 16'h0096; #100;
A = 16'h0091; B = 16'h0097; #100;
A = 16'h0091; B = 16'h0098; #100;
A = 16'h0091; B = 16'h0099; #100;
A = 16'h0091; B = 16'h009A; #100;
A = 16'h0091; B = 16'h009B; #100;
A = 16'h0091; B = 16'h009C; #100;
A = 16'h0091; B = 16'h009D; #100;
A = 16'h0091; B = 16'h009E; #100;
A = 16'h0091; B = 16'h009F; #100;
A = 16'h0091; B = 16'h00A0; #100;
A = 16'h0091; B = 16'h00A1; #100;
A = 16'h0091; B = 16'h00A2; #100;
A = 16'h0091; B = 16'h00A3; #100;
A = 16'h0091; B = 16'h00A4; #100;
A = 16'h0091; B = 16'h00A5; #100;
A = 16'h0091; B = 16'h00A6; #100;
A = 16'h0091; B = 16'h00A7; #100;
A = 16'h0091; B = 16'h00A8; #100;
A = 16'h0091; B = 16'h00A9; #100;
A = 16'h0091; B = 16'h00AA; #100;
A = 16'h0091; B = 16'h00AB; #100;
A = 16'h0091; B = 16'h00AC; #100;
A = 16'h0091; B = 16'h00AD; #100;
A = 16'h0091; B = 16'h00AE; #100;
A = 16'h0091; B = 16'h00AF; #100;
A = 16'h0091; B = 16'h00B0; #100;
A = 16'h0091; B = 16'h00B1; #100;
A = 16'h0091; B = 16'h00B2; #100;
A = 16'h0091; B = 16'h00B3; #100;
A = 16'h0091; B = 16'h00B4; #100;
A = 16'h0091; B = 16'h00B5; #100;
A = 16'h0091; B = 16'h00B6; #100;
A = 16'h0091; B = 16'h00B7; #100;
A = 16'h0091; B = 16'h00B8; #100;
A = 16'h0091; B = 16'h00B9; #100;
A = 16'h0091; B = 16'h00BA; #100;
A = 16'h0091; B = 16'h00BB; #100;
A = 16'h0091; B = 16'h00BC; #100;
A = 16'h0091; B = 16'h00BD; #100;
A = 16'h0091; B = 16'h00BE; #100;
A = 16'h0091; B = 16'h00BF; #100;
A = 16'h0091; B = 16'h00C0; #100;
A = 16'h0091; B = 16'h00C1; #100;
A = 16'h0091; B = 16'h00C2; #100;
A = 16'h0091; B = 16'h00C3; #100;
A = 16'h0091; B = 16'h00C4; #100;
A = 16'h0091; B = 16'h00C5; #100;
A = 16'h0091; B = 16'h00C6; #100;
A = 16'h0091; B = 16'h00C7; #100;
A = 16'h0091; B = 16'h00C8; #100;
A = 16'h0091; B = 16'h00C9; #100;
A = 16'h0091; B = 16'h00CA; #100;
A = 16'h0091; B = 16'h00CB; #100;
A = 16'h0091; B = 16'h00CC; #100;
A = 16'h0091; B = 16'h00CD; #100;
A = 16'h0091; B = 16'h00CE; #100;
A = 16'h0091; B = 16'h00CF; #100;
A = 16'h0091; B = 16'h00D0; #100;
A = 16'h0091; B = 16'h00D1; #100;
A = 16'h0091; B = 16'h00D2; #100;
A = 16'h0091; B = 16'h00D3; #100;
A = 16'h0091; B = 16'h00D4; #100;
A = 16'h0091; B = 16'h00D5; #100;
A = 16'h0091; B = 16'h00D6; #100;
A = 16'h0091; B = 16'h00D7; #100;
A = 16'h0091; B = 16'h00D8; #100;
A = 16'h0091; B = 16'h00D9; #100;
A = 16'h0091; B = 16'h00DA; #100;
A = 16'h0091; B = 16'h00DB; #100;
A = 16'h0091; B = 16'h00DC; #100;
A = 16'h0091; B = 16'h00DD; #100;
A = 16'h0091; B = 16'h00DE; #100;
A = 16'h0091; B = 16'h00DF; #100;
A = 16'h0091; B = 16'h00E0; #100;
A = 16'h0091; B = 16'h00E1; #100;
A = 16'h0091; B = 16'h00E2; #100;
A = 16'h0091; B = 16'h00E3; #100;
A = 16'h0091; B = 16'h00E4; #100;
A = 16'h0091; B = 16'h00E5; #100;
A = 16'h0091; B = 16'h00E6; #100;
A = 16'h0091; B = 16'h00E7; #100;
A = 16'h0091; B = 16'h00E8; #100;
A = 16'h0091; B = 16'h00E9; #100;
A = 16'h0091; B = 16'h00EA; #100;
A = 16'h0091; B = 16'h00EB; #100;
A = 16'h0091; B = 16'h00EC; #100;
A = 16'h0091; B = 16'h00ED; #100;
A = 16'h0091; B = 16'h00EE; #100;
A = 16'h0091; B = 16'h00EF; #100;
A = 16'h0091; B = 16'h00F0; #100;
A = 16'h0091; B = 16'h00F1; #100;
A = 16'h0091; B = 16'h00F2; #100;
A = 16'h0091; B = 16'h00F3; #100;
A = 16'h0091; B = 16'h00F4; #100;
A = 16'h0091; B = 16'h00F5; #100;
A = 16'h0091; B = 16'h00F6; #100;
A = 16'h0091; B = 16'h00F7; #100;
A = 16'h0091; B = 16'h00F8; #100;
A = 16'h0091; B = 16'h00F9; #100;
A = 16'h0091; B = 16'h00FA; #100;
A = 16'h0091; B = 16'h00FB; #100;
A = 16'h0091; B = 16'h00FC; #100;
A = 16'h0091; B = 16'h00FD; #100;
A = 16'h0091; B = 16'h00FE; #100;
A = 16'h0091; B = 16'h00FF; #100;
A = 16'h0092; B = 16'h000; #100;
A = 16'h0092; B = 16'h001; #100;
A = 16'h0092; B = 16'h002; #100;
A = 16'h0092; B = 16'h003; #100;
A = 16'h0092; B = 16'h004; #100;
A = 16'h0092; B = 16'h005; #100;
A = 16'h0092; B = 16'h006; #100;
A = 16'h0092; B = 16'h007; #100;
A = 16'h0092; B = 16'h008; #100;
A = 16'h0092; B = 16'h009; #100;
A = 16'h0092; B = 16'h00A; #100;
A = 16'h0092; B = 16'h00B; #100;
A = 16'h0092; B = 16'h00C; #100;
A = 16'h0092; B = 16'h00D; #100;
A = 16'h0092; B = 16'h00E; #100;
A = 16'h0092; B = 16'h00F; #100;
A = 16'h0092; B = 16'h0010; #100;
A = 16'h0092; B = 16'h0011; #100;
A = 16'h0092; B = 16'h0012; #100;
A = 16'h0092; B = 16'h0013; #100;
A = 16'h0092; B = 16'h0014; #100;
A = 16'h0092; B = 16'h0015; #100;
A = 16'h0092; B = 16'h0016; #100;
A = 16'h0092; B = 16'h0017; #100;
A = 16'h0092; B = 16'h0018; #100;
A = 16'h0092; B = 16'h0019; #100;
A = 16'h0092; B = 16'h001A; #100;
A = 16'h0092; B = 16'h001B; #100;
A = 16'h0092; B = 16'h001C; #100;
A = 16'h0092; B = 16'h001D; #100;
A = 16'h0092; B = 16'h001E; #100;
A = 16'h0092; B = 16'h001F; #100;
A = 16'h0092; B = 16'h0020; #100;
A = 16'h0092; B = 16'h0021; #100;
A = 16'h0092; B = 16'h0022; #100;
A = 16'h0092; B = 16'h0023; #100;
A = 16'h0092; B = 16'h0024; #100;
A = 16'h0092; B = 16'h0025; #100;
A = 16'h0092; B = 16'h0026; #100;
A = 16'h0092; B = 16'h0027; #100;
A = 16'h0092; B = 16'h0028; #100;
A = 16'h0092; B = 16'h0029; #100;
A = 16'h0092; B = 16'h002A; #100;
A = 16'h0092; B = 16'h002B; #100;
A = 16'h0092; B = 16'h002C; #100;
A = 16'h0092; B = 16'h002D; #100;
A = 16'h0092; B = 16'h002E; #100;
A = 16'h0092; B = 16'h002F; #100;
A = 16'h0092; B = 16'h0030; #100;
A = 16'h0092; B = 16'h0031; #100;
A = 16'h0092; B = 16'h0032; #100;
A = 16'h0092; B = 16'h0033; #100;
A = 16'h0092; B = 16'h0034; #100;
A = 16'h0092; B = 16'h0035; #100;
A = 16'h0092; B = 16'h0036; #100;
A = 16'h0092; B = 16'h0037; #100;
A = 16'h0092; B = 16'h0038; #100;
A = 16'h0092; B = 16'h0039; #100;
A = 16'h0092; B = 16'h003A; #100;
A = 16'h0092; B = 16'h003B; #100;
A = 16'h0092; B = 16'h003C; #100;
A = 16'h0092; B = 16'h003D; #100;
A = 16'h0092; B = 16'h003E; #100;
A = 16'h0092; B = 16'h003F; #100;
A = 16'h0092; B = 16'h0040; #100;
A = 16'h0092; B = 16'h0041; #100;
A = 16'h0092; B = 16'h0042; #100;
A = 16'h0092; B = 16'h0043; #100;
A = 16'h0092; B = 16'h0044; #100;
A = 16'h0092; B = 16'h0045; #100;
A = 16'h0092; B = 16'h0046; #100;
A = 16'h0092; B = 16'h0047; #100;
A = 16'h0092; B = 16'h0048; #100;
A = 16'h0092; B = 16'h0049; #100;
A = 16'h0092; B = 16'h004A; #100;
A = 16'h0092; B = 16'h004B; #100;
A = 16'h0092; B = 16'h004C; #100;
A = 16'h0092; B = 16'h004D; #100;
A = 16'h0092; B = 16'h004E; #100;
A = 16'h0092; B = 16'h004F; #100;
A = 16'h0092; B = 16'h0050; #100;
A = 16'h0092; B = 16'h0051; #100;
A = 16'h0092; B = 16'h0052; #100;
A = 16'h0092; B = 16'h0053; #100;
A = 16'h0092; B = 16'h0054; #100;
A = 16'h0092; B = 16'h0055; #100;
A = 16'h0092; B = 16'h0056; #100;
A = 16'h0092; B = 16'h0057; #100;
A = 16'h0092; B = 16'h0058; #100;
A = 16'h0092; B = 16'h0059; #100;
A = 16'h0092; B = 16'h005A; #100;
A = 16'h0092; B = 16'h005B; #100;
A = 16'h0092; B = 16'h005C; #100;
A = 16'h0092; B = 16'h005D; #100;
A = 16'h0092; B = 16'h005E; #100;
A = 16'h0092; B = 16'h005F; #100;
A = 16'h0092; B = 16'h0060; #100;
A = 16'h0092; B = 16'h0061; #100;
A = 16'h0092; B = 16'h0062; #100;
A = 16'h0092; B = 16'h0063; #100;
A = 16'h0092; B = 16'h0064; #100;
A = 16'h0092; B = 16'h0065; #100;
A = 16'h0092; B = 16'h0066; #100;
A = 16'h0092; B = 16'h0067; #100;
A = 16'h0092; B = 16'h0068; #100;
A = 16'h0092; B = 16'h0069; #100;
A = 16'h0092; B = 16'h006A; #100;
A = 16'h0092; B = 16'h006B; #100;
A = 16'h0092; B = 16'h006C; #100;
A = 16'h0092; B = 16'h006D; #100;
A = 16'h0092; B = 16'h006E; #100;
A = 16'h0092; B = 16'h006F; #100;
A = 16'h0092; B = 16'h0070; #100;
A = 16'h0092; B = 16'h0071; #100;
A = 16'h0092; B = 16'h0072; #100;
A = 16'h0092; B = 16'h0073; #100;
A = 16'h0092; B = 16'h0074; #100;
A = 16'h0092; B = 16'h0075; #100;
A = 16'h0092; B = 16'h0076; #100;
A = 16'h0092; B = 16'h0077; #100;
A = 16'h0092; B = 16'h0078; #100;
A = 16'h0092; B = 16'h0079; #100;
A = 16'h0092; B = 16'h007A; #100;
A = 16'h0092; B = 16'h007B; #100;
A = 16'h0092; B = 16'h007C; #100;
A = 16'h0092; B = 16'h007D; #100;
A = 16'h0092; B = 16'h007E; #100;
A = 16'h0092; B = 16'h007F; #100;
A = 16'h0092; B = 16'h0080; #100;
A = 16'h0092; B = 16'h0081; #100;
A = 16'h0092; B = 16'h0082; #100;
A = 16'h0092; B = 16'h0083; #100;
A = 16'h0092; B = 16'h0084; #100;
A = 16'h0092; B = 16'h0085; #100;
A = 16'h0092; B = 16'h0086; #100;
A = 16'h0092; B = 16'h0087; #100;
A = 16'h0092; B = 16'h0088; #100;
A = 16'h0092; B = 16'h0089; #100;
A = 16'h0092; B = 16'h008A; #100;
A = 16'h0092; B = 16'h008B; #100;
A = 16'h0092; B = 16'h008C; #100;
A = 16'h0092; B = 16'h008D; #100;
A = 16'h0092; B = 16'h008E; #100;
A = 16'h0092; B = 16'h008F; #100;
A = 16'h0092; B = 16'h0090; #100;
A = 16'h0092; B = 16'h0091; #100;
A = 16'h0092; B = 16'h0092; #100;
A = 16'h0092; B = 16'h0093; #100;
A = 16'h0092; B = 16'h0094; #100;
A = 16'h0092; B = 16'h0095; #100;
A = 16'h0092; B = 16'h0096; #100;
A = 16'h0092; B = 16'h0097; #100;
A = 16'h0092; B = 16'h0098; #100;
A = 16'h0092; B = 16'h0099; #100;
A = 16'h0092; B = 16'h009A; #100;
A = 16'h0092; B = 16'h009B; #100;
A = 16'h0092; B = 16'h009C; #100;
A = 16'h0092; B = 16'h009D; #100;
A = 16'h0092; B = 16'h009E; #100;
A = 16'h0092; B = 16'h009F; #100;
A = 16'h0092; B = 16'h00A0; #100;
A = 16'h0092; B = 16'h00A1; #100;
A = 16'h0092; B = 16'h00A2; #100;
A = 16'h0092; B = 16'h00A3; #100;
A = 16'h0092; B = 16'h00A4; #100;
A = 16'h0092; B = 16'h00A5; #100;
A = 16'h0092; B = 16'h00A6; #100;
A = 16'h0092; B = 16'h00A7; #100;
A = 16'h0092; B = 16'h00A8; #100;
A = 16'h0092; B = 16'h00A9; #100;
A = 16'h0092; B = 16'h00AA; #100;
A = 16'h0092; B = 16'h00AB; #100;
A = 16'h0092; B = 16'h00AC; #100;
A = 16'h0092; B = 16'h00AD; #100;
A = 16'h0092; B = 16'h00AE; #100;
A = 16'h0092; B = 16'h00AF; #100;
A = 16'h0092; B = 16'h00B0; #100;
A = 16'h0092; B = 16'h00B1; #100;
A = 16'h0092; B = 16'h00B2; #100;
A = 16'h0092; B = 16'h00B3; #100;
A = 16'h0092; B = 16'h00B4; #100;
A = 16'h0092; B = 16'h00B5; #100;
A = 16'h0092; B = 16'h00B6; #100;
A = 16'h0092; B = 16'h00B7; #100;
A = 16'h0092; B = 16'h00B8; #100;
A = 16'h0092; B = 16'h00B9; #100;
A = 16'h0092; B = 16'h00BA; #100;
A = 16'h0092; B = 16'h00BB; #100;
A = 16'h0092; B = 16'h00BC; #100;
A = 16'h0092; B = 16'h00BD; #100;
A = 16'h0092; B = 16'h00BE; #100;
A = 16'h0092; B = 16'h00BF; #100;
A = 16'h0092; B = 16'h00C0; #100;
A = 16'h0092; B = 16'h00C1; #100;
A = 16'h0092; B = 16'h00C2; #100;
A = 16'h0092; B = 16'h00C3; #100;
A = 16'h0092; B = 16'h00C4; #100;
A = 16'h0092; B = 16'h00C5; #100;
A = 16'h0092; B = 16'h00C6; #100;
A = 16'h0092; B = 16'h00C7; #100;
A = 16'h0092; B = 16'h00C8; #100;
A = 16'h0092; B = 16'h00C9; #100;
A = 16'h0092; B = 16'h00CA; #100;
A = 16'h0092; B = 16'h00CB; #100;
A = 16'h0092; B = 16'h00CC; #100;
A = 16'h0092; B = 16'h00CD; #100;
A = 16'h0092; B = 16'h00CE; #100;
A = 16'h0092; B = 16'h00CF; #100;
A = 16'h0092; B = 16'h00D0; #100;
A = 16'h0092; B = 16'h00D1; #100;
A = 16'h0092; B = 16'h00D2; #100;
A = 16'h0092; B = 16'h00D3; #100;
A = 16'h0092; B = 16'h00D4; #100;
A = 16'h0092; B = 16'h00D5; #100;
A = 16'h0092; B = 16'h00D6; #100;
A = 16'h0092; B = 16'h00D7; #100;
A = 16'h0092; B = 16'h00D8; #100;
A = 16'h0092; B = 16'h00D9; #100;
A = 16'h0092; B = 16'h00DA; #100;
A = 16'h0092; B = 16'h00DB; #100;
A = 16'h0092; B = 16'h00DC; #100;
A = 16'h0092; B = 16'h00DD; #100;
A = 16'h0092; B = 16'h00DE; #100;
A = 16'h0092; B = 16'h00DF; #100;
A = 16'h0092; B = 16'h00E0; #100;
A = 16'h0092; B = 16'h00E1; #100;
A = 16'h0092; B = 16'h00E2; #100;
A = 16'h0092; B = 16'h00E3; #100;
A = 16'h0092; B = 16'h00E4; #100;
A = 16'h0092; B = 16'h00E5; #100;
A = 16'h0092; B = 16'h00E6; #100;
A = 16'h0092; B = 16'h00E7; #100;
A = 16'h0092; B = 16'h00E8; #100;
A = 16'h0092; B = 16'h00E9; #100;
A = 16'h0092; B = 16'h00EA; #100;
A = 16'h0092; B = 16'h00EB; #100;
A = 16'h0092; B = 16'h00EC; #100;
A = 16'h0092; B = 16'h00ED; #100;
A = 16'h0092; B = 16'h00EE; #100;
A = 16'h0092; B = 16'h00EF; #100;
A = 16'h0092; B = 16'h00F0; #100;
A = 16'h0092; B = 16'h00F1; #100;
A = 16'h0092; B = 16'h00F2; #100;
A = 16'h0092; B = 16'h00F3; #100;
A = 16'h0092; B = 16'h00F4; #100;
A = 16'h0092; B = 16'h00F5; #100;
A = 16'h0092; B = 16'h00F6; #100;
A = 16'h0092; B = 16'h00F7; #100;
A = 16'h0092; B = 16'h00F8; #100;
A = 16'h0092; B = 16'h00F9; #100;
A = 16'h0092; B = 16'h00FA; #100;
A = 16'h0092; B = 16'h00FB; #100;
A = 16'h0092; B = 16'h00FC; #100;
A = 16'h0092; B = 16'h00FD; #100;
A = 16'h0092; B = 16'h00FE; #100;
A = 16'h0092; B = 16'h00FF; #100;
A = 16'h0093; B = 16'h000; #100;
A = 16'h0093; B = 16'h001; #100;
A = 16'h0093; B = 16'h002; #100;
A = 16'h0093; B = 16'h003; #100;
A = 16'h0093; B = 16'h004; #100;
A = 16'h0093; B = 16'h005; #100;
A = 16'h0093; B = 16'h006; #100;
A = 16'h0093; B = 16'h007; #100;
A = 16'h0093; B = 16'h008; #100;
A = 16'h0093; B = 16'h009; #100;
A = 16'h0093; B = 16'h00A; #100;
A = 16'h0093; B = 16'h00B; #100;
A = 16'h0093; B = 16'h00C; #100;
A = 16'h0093; B = 16'h00D; #100;
A = 16'h0093; B = 16'h00E; #100;
A = 16'h0093; B = 16'h00F; #100;
A = 16'h0093; B = 16'h0010; #100;
A = 16'h0093; B = 16'h0011; #100;
A = 16'h0093; B = 16'h0012; #100;
A = 16'h0093; B = 16'h0013; #100;
A = 16'h0093; B = 16'h0014; #100;
A = 16'h0093; B = 16'h0015; #100;
A = 16'h0093; B = 16'h0016; #100;
A = 16'h0093; B = 16'h0017; #100;
A = 16'h0093; B = 16'h0018; #100;
A = 16'h0093; B = 16'h0019; #100;
A = 16'h0093; B = 16'h001A; #100;
A = 16'h0093; B = 16'h001B; #100;
A = 16'h0093; B = 16'h001C; #100;
A = 16'h0093; B = 16'h001D; #100;
A = 16'h0093; B = 16'h001E; #100;
A = 16'h0093; B = 16'h001F; #100;
A = 16'h0093; B = 16'h0020; #100;
A = 16'h0093; B = 16'h0021; #100;
A = 16'h0093; B = 16'h0022; #100;
A = 16'h0093; B = 16'h0023; #100;
A = 16'h0093; B = 16'h0024; #100;
A = 16'h0093; B = 16'h0025; #100;
A = 16'h0093; B = 16'h0026; #100;
A = 16'h0093; B = 16'h0027; #100;
A = 16'h0093; B = 16'h0028; #100;
A = 16'h0093; B = 16'h0029; #100;
A = 16'h0093; B = 16'h002A; #100;
A = 16'h0093; B = 16'h002B; #100;
A = 16'h0093; B = 16'h002C; #100;
A = 16'h0093; B = 16'h002D; #100;
A = 16'h0093; B = 16'h002E; #100;
A = 16'h0093; B = 16'h002F; #100;
A = 16'h0093; B = 16'h0030; #100;
A = 16'h0093; B = 16'h0031; #100;
A = 16'h0093; B = 16'h0032; #100;
A = 16'h0093; B = 16'h0033; #100;
A = 16'h0093; B = 16'h0034; #100;
A = 16'h0093; B = 16'h0035; #100;
A = 16'h0093; B = 16'h0036; #100;
A = 16'h0093; B = 16'h0037; #100;
A = 16'h0093; B = 16'h0038; #100;
A = 16'h0093; B = 16'h0039; #100;
A = 16'h0093; B = 16'h003A; #100;
A = 16'h0093; B = 16'h003B; #100;
A = 16'h0093; B = 16'h003C; #100;
A = 16'h0093; B = 16'h003D; #100;
A = 16'h0093; B = 16'h003E; #100;
A = 16'h0093; B = 16'h003F; #100;
A = 16'h0093; B = 16'h0040; #100;
A = 16'h0093; B = 16'h0041; #100;
A = 16'h0093; B = 16'h0042; #100;
A = 16'h0093; B = 16'h0043; #100;
A = 16'h0093; B = 16'h0044; #100;
A = 16'h0093; B = 16'h0045; #100;
A = 16'h0093; B = 16'h0046; #100;
A = 16'h0093; B = 16'h0047; #100;
A = 16'h0093; B = 16'h0048; #100;
A = 16'h0093; B = 16'h0049; #100;
A = 16'h0093; B = 16'h004A; #100;
A = 16'h0093; B = 16'h004B; #100;
A = 16'h0093; B = 16'h004C; #100;
A = 16'h0093; B = 16'h004D; #100;
A = 16'h0093; B = 16'h004E; #100;
A = 16'h0093; B = 16'h004F; #100;
A = 16'h0093; B = 16'h0050; #100;
A = 16'h0093; B = 16'h0051; #100;
A = 16'h0093; B = 16'h0052; #100;
A = 16'h0093; B = 16'h0053; #100;
A = 16'h0093; B = 16'h0054; #100;
A = 16'h0093; B = 16'h0055; #100;
A = 16'h0093; B = 16'h0056; #100;
A = 16'h0093; B = 16'h0057; #100;
A = 16'h0093; B = 16'h0058; #100;
A = 16'h0093; B = 16'h0059; #100;
A = 16'h0093; B = 16'h005A; #100;
A = 16'h0093; B = 16'h005B; #100;
A = 16'h0093; B = 16'h005C; #100;
A = 16'h0093; B = 16'h005D; #100;
A = 16'h0093; B = 16'h005E; #100;
A = 16'h0093; B = 16'h005F; #100;
A = 16'h0093; B = 16'h0060; #100;
A = 16'h0093; B = 16'h0061; #100;
A = 16'h0093; B = 16'h0062; #100;
A = 16'h0093; B = 16'h0063; #100;
A = 16'h0093; B = 16'h0064; #100;
A = 16'h0093; B = 16'h0065; #100;
A = 16'h0093; B = 16'h0066; #100;
A = 16'h0093; B = 16'h0067; #100;
A = 16'h0093; B = 16'h0068; #100;
A = 16'h0093; B = 16'h0069; #100;
A = 16'h0093; B = 16'h006A; #100;
A = 16'h0093; B = 16'h006B; #100;
A = 16'h0093; B = 16'h006C; #100;
A = 16'h0093; B = 16'h006D; #100;
A = 16'h0093; B = 16'h006E; #100;
A = 16'h0093; B = 16'h006F; #100;
A = 16'h0093; B = 16'h0070; #100;
A = 16'h0093; B = 16'h0071; #100;
A = 16'h0093; B = 16'h0072; #100;
A = 16'h0093; B = 16'h0073; #100;
A = 16'h0093; B = 16'h0074; #100;
A = 16'h0093; B = 16'h0075; #100;
A = 16'h0093; B = 16'h0076; #100;
A = 16'h0093; B = 16'h0077; #100;
A = 16'h0093; B = 16'h0078; #100;
A = 16'h0093; B = 16'h0079; #100;
A = 16'h0093; B = 16'h007A; #100;
A = 16'h0093; B = 16'h007B; #100;
A = 16'h0093; B = 16'h007C; #100;
A = 16'h0093; B = 16'h007D; #100;
A = 16'h0093; B = 16'h007E; #100;
A = 16'h0093; B = 16'h007F; #100;
A = 16'h0093; B = 16'h0080; #100;
A = 16'h0093; B = 16'h0081; #100;
A = 16'h0093; B = 16'h0082; #100;
A = 16'h0093; B = 16'h0083; #100;
A = 16'h0093; B = 16'h0084; #100;
A = 16'h0093; B = 16'h0085; #100;
A = 16'h0093; B = 16'h0086; #100;
A = 16'h0093; B = 16'h0087; #100;
A = 16'h0093; B = 16'h0088; #100;
A = 16'h0093; B = 16'h0089; #100;
A = 16'h0093; B = 16'h008A; #100;
A = 16'h0093; B = 16'h008B; #100;
A = 16'h0093; B = 16'h008C; #100;
A = 16'h0093; B = 16'h008D; #100;
A = 16'h0093; B = 16'h008E; #100;
A = 16'h0093; B = 16'h008F; #100;
A = 16'h0093; B = 16'h0090; #100;
A = 16'h0093; B = 16'h0091; #100;
A = 16'h0093; B = 16'h0092; #100;
A = 16'h0093; B = 16'h0093; #100;
A = 16'h0093; B = 16'h0094; #100;
A = 16'h0093; B = 16'h0095; #100;
A = 16'h0093; B = 16'h0096; #100;
A = 16'h0093; B = 16'h0097; #100;
A = 16'h0093; B = 16'h0098; #100;
A = 16'h0093; B = 16'h0099; #100;
A = 16'h0093; B = 16'h009A; #100;
A = 16'h0093; B = 16'h009B; #100;
A = 16'h0093; B = 16'h009C; #100;
A = 16'h0093; B = 16'h009D; #100;
A = 16'h0093; B = 16'h009E; #100;
A = 16'h0093; B = 16'h009F; #100;
A = 16'h0093; B = 16'h00A0; #100;
A = 16'h0093; B = 16'h00A1; #100;
A = 16'h0093; B = 16'h00A2; #100;
A = 16'h0093; B = 16'h00A3; #100;
A = 16'h0093; B = 16'h00A4; #100;
A = 16'h0093; B = 16'h00A5; #100;
A = 16'h0093; B = 16'h00A6; #100;
A = 16'h0093; B = 16'h00A7; #100;
A = 16'h0093; B = 16'h00A8; #100;
A = 16'h0093; B = 16'h00A9; #100;
A = 16'h0093; B = 16'h00AA; #100;
A = 16'h0093; B = 16'h00AB; #100;
A = 16'h0093; B = 16'h00AC; #100;
A = 16'h0093; B = 16'h00AD; #100;
A = 16'h0093; B = 16'h00AE; #100;
A = 16'h0093; B = 16'h00AF; #100;
A = 16'h0093; B = 16'h00B0; #100;
A = 16'h0093; B = 16'h00B1; #100;
A = 16'h0093; B = 16'h00B2; #100;
A = 16'h0093; B = 16'h00B3; #100;
A = 16'h0093; B = 16'h00B4; #100;
A = 16'h0093; B = 16'h00B5; #100;
A = 16'h0093; B = 16'h00B6; #100;
A = 16'h0093; B = 16'h00B7; #100;
A = 16'h0093; B = 16'h00B8; #100;
A = 16'h0093; B = 16'h00B9; #100;
A = 16'h0093; B = 16'h00BA; #100;
A = 16'h0093; B = 16'h00BB; #100;
A = 16'h0093; B = 16'h00BC; #100;
A = 16'h0093; B = 16'h00BD; #100;
A = 16'h0093; B = 16'h00BE; #100;
A = 16'h0093; B = 16'h00BF; #100;
A = 16'h0093; B = 16'h00C0; #100;
A = 16'h0093; B = 16'h00C1; #100;
A = 16'h0093; B = 16'h00C2; #100;
A = 16'h0093; B = 16'h00C3; #100;
A = 16'h0093; B = 16'h00C4; #100;
A = 16'h0093; B = 16'h00C5; #100;
A = 16'h0093; B = 16'h00C6; #100;
A = 16'h0093; B = 16'h00C7; #100;
A = 16'h0093; B = 16'h00C8; #100;
A = 16'h0093; B = 16'h00C9; #100;
A = 16'h0093; B = 16'h00CA; #100;
A = 16'h0093; B = 16'h00CB; #100;
A = 16'h0093; B = 16'h00CC; #100;
A = 16'h0093; B = 16'h00CD; #100;
A = 16'h0093; B = 16'h00CE; #100;
A = 16'h0093; B = 16'h00CF; #100;
A = 16'h0093; B = 16'h00D0; #100;
A = 16'h0093; B = 16'h00D1; #100;
A = 16'h0093; B = 16'h00D2; #100;
A = 16'h0093; B = 16'h00D3; #100;
A = 16'h0093; B = 16'h00D4; #100;
A = 16'h0093; B = 16'h00D5; #100;
A = 16'h0093; B = 16'h00D6; #100;
A = 16'h0093; B = 16'h00D7; #100;
A = 16'h0093; B = 16'h00D8; #100;
A = 16'h0093; B = 16'h00D9; #100;
A = 16'h0093; B = 16'h00DA; #100;
A = 16'h0093; B = 16'h00DB; #100;
A = 16'h0093; B = 16'h00DC; #100;
A = 16'h0093; B = 16'h00DD; #100;
A = 16'h0093; B = 16'h00DE; #100;
A = 16'h0093; B = 16'h00DF; #100;
A = 16'h0093; B = 16'h00E0; #100;
A = 16'h0093; B = 16'h00E1; #100;
A = 16'h0093; B = 16'h00E2; #100;
A = 16'h0093; B = 16'h00E3; #100;
A = 16'h0093; B = 16'h00E4; #100;
A = 16'h0093; B = 16'h00E5; #100;
A = 16'h0093; B = 16'h00E6; #100;
A = 16'h0093; B = 16'h00E7; #100;
A = 16'h0093; B = 16'h00E8; #100;
A = 16'h0093; B = 16'h00E9; #100;
A = 16'h0093; B = 16'h00EA; #100;
A = 16'h0093; B = 16'h00EB; #100;
A = 16'h0093; B = 16'h00EC; #100;
A = 16'h0093; B = 16'h00ED; #100;
A = 16'h0093; B = 16'h00EE; #100;
A = 16'h0093; B = 16'h00EF; #100;
A = 16'h0093; B = 16'h00F0; #100;
A = 16'h0093; B = 16'h00F1; #100;
A = 16'h0093; B = 16'h00F2; #100;
A = 16'h0093; B = 16'h00F3; #100;
A = 16'h0093; B = 16'h00F4; #100;
A = 16'h0093; B = 16'h00F5; #100;
A = 16'h0093; B = 16'h00F6; #100;
A = 16'h0093; B = 16'h00F7; #100;
A = 16'h0093; B = 16'h00F8; #100;
A = 16'h0093; B = 16'h00F9; #100;
A = 16'h0093; B = 16'h00FA; #100;
A = 16'h0093; B = 16'h00FB; #100;
A = 16'h0093; B = 16'h00FC; #100;
A = 16'h0093; B = 16'h00FD; #100;
A = 16'h0093; B = 16'h00FE; #100;
A = 16'h0093; B = 16'h00FF; #100;
A = 16'h0094; B = 16'h000; #100;
A = 16'h0094; B = 16'h001; #100;
A = 16'h0094; B = 16'h002; #100;
A = 16'h0094; B = 16'h003; #100;
A = 16'h0094; B = 16'h004; #100;
A = 16'h0094; B = 16'h005; #100;
A = 16'h0094; B = 16'h006; #100;
A = 16'h0094; B = 16'h007; #100;
A = 16'h0094; B = 16'h008; #100;
A = 16'h0094; B = 16'h009; #100;
A = 16'h0094; B = 16'h00A; #100;
A = 16'h0094; B = 16'h00B; #100;
A = 16'h0094; B = 16'h00C; #100;
A = 16'h0094; B = 16'h00D; #100;
A = 16'h0094; B = 16'h00E; #100;
A = 16'h0094; B = 16'h00F; #100;
A = 16'h0094; B = 16'h0010; #100;
A = 16'h0094; B = 16'h0011; #100;
A = 16'h0094; B = 16'h0012; #100;
A = 16'h0094; B = 16'h0013; #100;
A = 16'h0094; B = 16'h0014; #100;
A = 16'h0094; B = 16'h0015; #100;
A = 16'h0094; B = 16'h0016; #100;
A = 16'h0094; B = 16'h0017; #100;
A = 16'h0094; B = 16'h0018; #100;
A = 16'h0094; B = 16'h0019; #100;
A = 16'h0094; B = 16'h001A; #100;
A = 16'h0094; B = 16'h001B; #100;
A = 16'h0094; B = 16'h001C; #100;
A = 16'h0094; B = 16'h001D; #100;
A = 16'h0094; B = 16'h001E; #100;
A = 16'h0094; B = 16'h001F; #100;
A = 16'h0094; B = 16'h0020; #100;
A = 16'h0094; B = 16'h0021; #100;
A = 16'h0094; B = 16'h0022; #100;
A = 16'h0094; B = 16'h0023; #100;
A = 16'h0094; B = 16'h0024; #100;
A = 16'h0094; B = 16'h0025; #100;
A = 16'h0094; B = 16'h0026; #100;
A = 16'h0094; B = 16'h0027; #100;
A = 16'h0094; B = 16'h0028; #100;
A = 16'h0094; B = 16'h0029; #100;
A = 16'h0094; B = 16'h002A; #100;
A = 16'h0094; B = 16'h002B; #100;
A = 16'h0094; B = 16'h002C; #100;
A = 16'h0094; B = 16'h002D; #100;
A = 16'h0094; B = 16'h002E; #100;
A = 16'h0094; B = 16'h002F; #100;
A = 16'h0094; B = 16'h0030; #100;
A = 16'h0094; B = 16'h0031; #100;
A = 16'h0094; B = 16'h0032; #100;
A = 16'h0094; B = 16'h0033; #100;
A = 16'h0094; B = 16'h0034; #100;
A = 16'h0094; B = 16'h0035; #100;
A = 16'h0094; B = 16'h0036; #100;
A = 16'h0094; B = 16'h0037; #100;
A = 16'h0094; B = 16'h0038; #100;
A = 16'h0094; B = 16'h0039; #100;
A = 16'h0094; B = 16'h003A; #100;
A = 16'h0094; B = 16'h003B; #100;
A = 16'h0094; B = 16'h003C; #100;
A = 16'h0094; B = 16'h003D; #100;
A = 16'h0094; B = 16'h003E; #100;
A = 16'h0094; B = 16'h003F; #100;
A = 16'h0094; B = 16'h0040; #100;
A = 16'h0094; B = 16'h0041; #100;
A = 16'h0094; B = 16'h0042; #100;
A = 16'h0094; B = 16'h0043; #100;
A = 16'h0094; B = 16'h0044; #100;
A = 16'h0094; B = 16'h0045; #100;
A = 16'h0094; B = 16'h0046; #100;
A = 16'h0094; B = 16'h0047; #100;
A = 16'h0094; B = 16'h0048; #100;
A = 16'h0094; B = 16'h0049; #100;
A = 16'h0094; B = 16'h004A; #100;
A = 16'h0094; B = 16'h004B; #100;
A = 16'h0094; B = 16'h004C; #100;
A = 16'h0094; B = 16'h004D; #100;
A = 16'h0094; B = 16'h004E; #100;
A = 16'h0094; B = 16'h004F; #100;
A = 16'h0094; B = 16'h0050; #100;
A = 16'h0094; B = 16'h0051; #100;
A = 16'h0094; B = 16'h0052; #100;
A = 16'h0094; B = 16'h0053; #100;
A = 16'h0094; B = 16'h0054; #100;
A = 16'h0094; B = 16'h0055; #100;
A = 16'h0094; B = 16'h0056; #100;
A = 16'h0094; B = 16'h0057; #100;
A = 16'h0094; B = 16'h0058; #100;
A = 16'h0094; B = 16'h0059; #100;
A = 16'h0094; B = 16'h005A; #100;
A = 16'h0094; B = 16'h005B; #100;
A = 16'h0094; B = 16'h005C; #100;
A = 16'h0094; B = 16'h005D; #100;
A = 16'h0094; B = 16'h005E; #100;
A = 16'h0094; B = 16'h005F; #100;
A = 16'h0094; B = 16'h0060; #100;
A = 16'h0094; B = 16'h0061; #100;
A = 16'h0094; B = 16'h0062; #100;
A = 16'h0094; B = 16'h0063; #100;
A = 16'h0094; B = 16'h0064; #100;
A = 16'h0094; B = 16'h0065; #100;
A = 16'h0094; B = 16'h0066; #100;
A = 16'h0094; B = 16'h0067; #100;
A = 16'h0094; B = 16'h0068; #100;
A = 16'h0094; B = 16'h0069; #100;
A = 16'h0094; B = 16'h006A; #100;
A = 16'h0094; B = 16'h006B; #100;
A = 16'h0094; B = 16'h006C; #100;
A = 16'h0094; B = 16'h006D; #100;
A = 16'h0094; B = 16'h006E; #100;
A = 16'h0094; B = 16'h006F; #100;
A = 16'h0094; B = 16'h0070; #100;
A = 16'h0094; B = 16'h0071; #100;
A = 16'h0094; B = 16'h0072; #100;
A = 16'h0094; B = 16'h0073; #100;
A = 16'h0094; B = 16'h0074; #100;
A = 16'h0094; B = 16'h0075; #100;
A = 16'h0094; B = 16'h0076; #100;
A = 16'h0094; B = 16'h0077; #100;
A = 16'h0094; B = 16'h0078; #100;
A = 16'h0094; B = 16'h0079; #100;
A = 16'h0094; B = 16'h007A; #100;
A = 16'h0094; B = 16'h007B; #100;
A = 16'h0094; B = 16'h007C; #100;
A = 16'h0094; B = 16'h007D; #100;
A = 16'h0094; B = 16'h007E; #100;
A = 16'h0094; B = 16'h007F; #100;
A = 16'h0094; B = 16'h0080; #100;
A = 16'h0094; B = 16'h0081; #100;
A = 16'h0094; B = 16'h0082; #100;
A = 16'h0094; B = 16'h0083; #100;
A = 16'h0094; B = 16'h0084; #100;
A = 16'h0094; B = 16'h0085; #100;
A = 16'h0094; B = 16'h0086; #100;
A = 16'h0094; B = 16'h0087; #100;
A = 16'h0094; B = 16'h0088; #100;
A = 16'h0094; B = 16'h0089; #100;
A = 16'h0094; B = 16'h008A; #100;
A = 16'h0094; B = 16'h008B; #100;
A = 16'h0094; B = 16'h008C; #100;
A = 16'h0094; B = 16'h008D; #100;
A = 16'h0094; B = 16'h008E; #100;
A = 16'h0094; B = 16'h008F; #100;
A = 16'h0094; B = 16'h0090; #100;
A = 16'h0094; B = 16'h0091; #100;
A = 16'h0094; B = 16'h0092; #100;
A = 16'h0094; B = 16'h0093; #100;
A = 16'h0094; B = 16'h0094; #100;
A = 16'h0094; B = 16'h0095; #100;
A = 16'h0094; B = 16'h0096; #100;
A = 16'h0094; B = 16'h0097; #100;
A = 16'h0094; B = 16'h0098; #100;
A = 16'h0094; B = 16'h0099; #100;
A = 16'h0094; B = 16'h009A; #100;
A = 16'h0094; B = 16'h009B; #100;
A = 16'h0094; B = 16'h009C; #100;
A = 16'h0094; B = 16'h009D; #100;
A = 16'h0094; B = 16'h009E; #100;
A = 16'h0094; B = 16'h009F; #100;
A = 16'h0094; B = 16'h00A0; #100;
A = 16'h0094; B = 16'h00A1; #100;
A = 16'h0094; B = 16'h00A2; #100;
A = 16'h0094; B = 16'h00A3; #100;
A = 16'h0094; B = 16'h00A4; #100;
A = 16'h0094; B = 16'h00A5; #100;
A = 16'h0094; B = 16'h00A6; #100;
A = 16'h0094; B = 16'h00A7; #100;
A = 16'h0094; B = 16'h00A8; #100;
A = 16'h0094; B = 16'h00A9; #100;
A = 16'h0094; B = 16'h00AA; #100;
A = 16'h0094; B = 16'h00AB; #100;
A = 16'h0094; B = 16'h00AC; #100;
A = 16'h0094; B = 16'h00AD; #100;
A = 16'h0094; B = 16'h00AE; #100;
A = 16'h0094; B = 16'h00AF; #100;
A = 16'h0094; B = 16'h00B0; #100;
A = 16'h0094; B = 16'h00B1; #100;
A = 16'h0094; B = 16'h00B2; #100;
A = 16'h0094; B = 16'h00B3; #100;
A = 16'h0094; B = 16'h00B4; #100;
A = 16'h0094; B = 16'h00B5; #100;
A = 16'h0094; B = 16'h00B6; #100;
A = 16'h0094; B = 16'h00B7; #100;
A = 16'h0094; B = 16'h00B8; #100;
A = 16'h0094; B = 16'h00B9; #100;
A = 16'h0094; B = 16'h00BA; #100;
A = 16'h0094; B = 16'h00BB; #100;
A = 16'h0094; B = 16'h00BC; #100;
A = 16'h0094; B = 16'h00BD; #100;
A = 16'h0094; B = 16'h00BE; #100;
A = 16'h0094; B = 16'h00BF; #100;
A = 16'h0094; B = 16'h00C0; #100;
A = 16'h0094; B = 16'h00C1; #100;
A = 16'h0094; B = 16'h00C2; #100;
A = 16'h0094; B = 16'h00C3; #100;
A = 16'h0094; B = 16'h00C4; #100;
A = 16'h0094; B = 16'h00C5; #100;
A = 16'h0094; B = 16'h00C6; #100;
A = 16'h0094; B = 16'h00C7; #100;
A = 16'h0094; B = 16'h00C8; #100;
A = 16'h0094; B = 16'h00C9; #100;
A = 16'h0094; B = 16'h00CA; #100;
A = 16'h0094; B = 16'h00CB; #100;
A = 16'h0094; B = 16'h00CC; #100;
A = 16'h0094; B = 16'h00CD; #100;
A = 16'h0094; B = 16'h00CE; #100;
A = 16'h0094; B = 16'h00CF; #100;
A = 16'h0094; B = 16'h00D0; #100;
A = 16'h0094; B = 16'h00D1; #100;
A = 16'h0094; B = 16'h00D2; #100;
A = 16'h0094; B = 16'h00D3; #100;
A = 16'h0094; B = 16'h00D4; #100;
A = 16'h0094; B = 16'h00D5; #100;
A = 16'h0094; B = 16'h00D6; #100;
A = 16'h0094; B = 16'h00D7; #100;
A = 16'h0094; B = 16'h00D8; #100;
A = 16'h0094; B = 16'h00D9; #100;
A = 16'h0094; B = 16'h00DA; #100;
A = 16'h0094; B = 16'h00DB; #100;
A = 16'h0094; B = 16'h00DC; #100;
A = 16'h0094; B = 16'h00DD; #100;
A = 16'h0094; B = 16'h00DE; #100;
A = 16'h0094; B = 16'h00DF; #100;
A = 16'h0094; B = 16'h00E0; #100;
A = 16'h0094; B = 16'h00E1; #100;
A = 16'h0094; B = 16'h00E2; #100;
A = 16'h0094; B = 16'h00E3; #100;
A = 16'h0094; B = 16'h00E4; #100;
A = 16'h0094; B = 16'h00E5; #100;
A = 16'h0094; B = 16'h00E6; #100;
A = 16'h0094; B = 16'h00E7; #100;
A = 16'h0094; B = 16'h00E8; #100;
A = 16'h0094; B = 16'h00E9; #100;
A = 16'h0094; B = 16'h00EA; #100;
A = 16'h0094; B = 16'h00EB; #100;
A = 16'h0094; B = 16'h00EC; #100;
A = 16'h0094; B = 16'h00ED; #100;
A = 16'h0094; B = 16'h00EE; #100;
A = 16'h0094; B = 16'h00EF; #100;
A = 16'h0094; B = 16'h00F0; #100;
A = 16'h0094; B = 16'h00F1; #100;
A = 16'h0094; B = 16'h00F2; #100;
A = 16'h0094; B = 16'h00F3; #100;
A = 16'h0094; B = 16'h00F4; #100;
A = 16'h0094; B = 16'h00F5; #100;
A = 16'h0094; B = 16'h00F6; #100;
A = 16'h0094; B = 16'h00F7; #100;
A = 16'h0094; B = 16'h00F8; #100;
A = 16'h0094; B = 16'h00F9; #100;
A = 16'h0094; B = 16'h00FA; #100;
A = 16'h0094; B = 16'h00FB; #100;
A = 16'h0094; B = 16'h00FC; #100;
A = 16'h0094; B = 16'h00FD; #100;
A = 16'h0094; B = 16'h00FE; #100;
A = 16'h0094; B = 16'h00FF; #100;
A = 16'h0095; B = 16'h000; #100;
A = 16'h0095; B = 16'h001; #100;
A = 16'h0095; B = 16'h002; #100;
A = 16'h0095; B = 16'h003; #100;
A = 16'h0095; B = 16'h004; #100;
A = 16'h0095; B = 16'h005; #100;
A = 16'h0095; B = 16'h006; #100;
A = 16'h0095; B = 16'h007; #100;
A = 16'h0095; B = 16'h008; #100;
A = 16'h0095; B = 16'h009; #100;
A = 16'h0095; B = 16'h00A; #100;
A = 16'h0095; B = 16'h00B; #100;
A = 16'h0095; B = 16'h00C; #100;
A = 16'h0095; B = 16'h00D; #100;
A = 16'h0095; B = 16'h00E; #100;
A = 16'h0095; B = 16'h00F; #100;
A = 16'h0095; B = 16'h0010; #100;
A = 16'h0095; B = 16'h0011; #100;
A = 16'h0095; B = 16'h0012; #100;
A = 16'h0095; B = 16'h0013; #100;
A = 16'h0095; B = 16'h0014; #100;
A = 16'h0095; B = 16'h0015; #100;
A = 16'h0095; B = 16'h0016; #100;
A = 16'h0095; B = 16'h0017; #100;
A = 16'h0095; B = 16'h0018; #100;
A = 16'h0095; B = 16'h0019; #100;
A = 16'h0095; B = 16'h001A; #100;
A = 16'h0095; B = 16'h001B; #100;
A = 16'h0095; B = 16'h001C; #100;
A = 16'h0095; B = 16'h001D; #100;
A = 16'h0095; B = 16'h001E; #100;
A = 16'h0095; B = 16'h001F; #100;
A = 16'h0095; B = 16'h0020; #100;
A = 16'h0095; B = 16'h0021; #100;
A = 16'h0095; B = 16'h0022; #100;
A = 16'h0095; B = 16'h0023; #100;
A = 16'h0095; B = 16'h0024; #100;
A = 16'h0095; B = 16'h0025; #100;
A = 16'h0095; B = 16'h0026; #100;
A = 16'h0095; B = 16'h0027; #100;
A = 16'h0095; B = 16'h0028; #100;
A = 16'h0095; B = 16'h0029; #100;
A = 16'h0095; B = 16'h002A; #100;
A = 16'h0095; B = 16'h002B; #100;
A = 16'h0095; B = 16'h002C; #100;
A = 16'h0095; B = 16'h002D; #100;
A = 16'h0095; B = 16'h002E; #100;
A = 16'h0095; B = 16'h002F; #100;
A = 16'h0095; B = 16'h0030; #100;
A = 16'h0095; B = 16'h0031; #100;
A = 16'h0095; B = 16'h0032; #100;
A = 16'h0095; B = 16'h0033; #100;
A = 16'h0095; B = 16'h0034; #100;
A = 16'h0095; B = 16'h0035; #100;
A = 16'h0095; B = 16'h0036; #100;
A = 16'h0095; B = 16'h0037; #100;
A = 16'h0095; B = 16'h0038; #100;
A = 16'h0095; B = 16'h0039; #100;
A = 16'h0095; B = 16'h003A; #100;
A = 16'h0095; B = 16'h003B; #100;
A = 16'h0095; B = 16'h003C; #100;
A = 16'h0095; B = 16'h003D; #100;
A = 16'h0095; B = 16'h003E; #100;
A = 16'h0095; B = 16'h003F; #100;
A = 16'h0095; B = 16'h0040; #100;
A = 16'h0095; B = 16'h0041; #100;
A = 16'h0095; B = 16'h0042; #100;
A = 16'h0095; B = 16'h0043; #100;
A = 16'h0095; B = 16'h0044; #100;
A = 16'h0095; B = 16'h0045; #100;
A = 16'h0095; B = 16'h0046; #100;
A = 16'h0095; B = 16'h0047; #100;
A = 16'h0095; B = 16'h0048; #100;
A = 16'h0095; B = 16'h0049; #100;
A = 16'h0095; B = 16'h004A; #100;
A = 16'h0095; B = 16'h004B; #100;
A = 16'h0095; B = 16'h004C; #100;
A = 16'h0095; B = 16'h004D; #100;
A = 16'h0095; B = 16'h004E; #100;
A = 16'h0095; B = 16'h004F; #100;
A = 16'h0095; B = 16'h0050; #100;
A = 16'h0095; B = 16'h0051; #100;
A = 16'h0095; B = 16'h0052; #100;
A = 16'h0095; B = 16'h0053; #100;
A = 16'h0095; B = 16'h0054; #100;
A = 16'h0095; B = 16'h0055; #100;
A = 16'h0095; B = 16'h0056; #100;
A = 16'h0095; B = 16'h0057; #100;
A = 16'h0095; B = 16'h0058; #100;
A = 16'h0095; B = 16'h0059; #100;
A = 16'h0095; B = 16'h005A; #100;
A = 16'h0095; B = 16'h005B; #100;
A = 16'h0095; B = 16'h005C; #100;
A = 16'h0095; B = 16'h005D; #100;
A = 16'h0095; B = 16'h005E; #100;
A = 16'h0095; B = 16'h005F; #100;
A = 16'h0095; B = 16'h0060; #100;
A = 16'h0095; B = 16'h0061; #100;
A = 16'h0095; B = 16'h0062; #100;
A = 16'h0095; B = 16'h0063; #100;
A = 16'h0095; B = 16'h0064; #100;
A = 16'h0095; B = 16'h0065; #100;
A = 16'h0095; B = 16'h0066; #100;
A = 16'h0095; B = 16'h0067; #100;
A = 16'h0095; B = 16'h0068; #100;
A = 16'h0095; B = 16'h0069; #100;
A = 16'h0095; B = 16'h006A; #100;
A = 16'h0095; B = 16'h006B; #100;
A = 16'h0095; B = 16'h006C; #100;
A = 16'h0095; B = 16'h006D; #100;
A = 16'h0095; B = 16'h006E; #100;
A = 16'h0095; B = 16'h006F; #100;
A = 16'h0095; B = 16'h0070; #100;
A = 16'h0095; B = 16'h0071; #100;
A = 16'h0095; B = 16'h0072; #100;
A = 16'h0095; B = 16'h0073; #100;
A = 16'h0095; B = 16'h0074; #100;
A = 16'h0095; B = 16'h0075; #100;
A = 16'h0095; B = 16'h0076; #100;
A = 16'h0095; B = 16'h0077; #100;
A = 16'h0095; B = 16'h0078; #100;
A = 16'h0095; B = 16'h0079; #100;
A = 16'h0095; B = 16'h007A; #100;
A = 16'h0095; B = 16'h007B; #100;
A = 16'h0095; B = 16'h007C; #100;
A = 16'h0095; B = 16'h007D; #100;
A = 16'h0095; B = 16'h007E; #100;
A = 16'h0095; B = 16'h007F; #100;
A = 16'h0095; B = 16'h0080; #100;
A = 16'h0095; B = 16'h0081; #100;
A = 16'h0095; B = 16'h0082; #100;
A = 16'h0095; B = 16'h0083; #100;
A = 16'h0095; B = 16'h0084; #100;
A = 16'h0095; B = 16'h0085; #100;
A = 16'h0095; B = 16'h0086; #100;
A = 16'h0095; B = 16'h0087; #100;
A = 16'h0095; B = 16'h0088; #100;
A = 16'h0095; B = 16'h0089; #100;
A = 16'h0095; B = 16'h008A; #100;
A = 16'h0095; B = 16'h008B; #100;
A = 16'h0095; B = 16'h008C; #100;
A = 16'h0095; B = 16'h008D; #100;
A = 16'h0095; B = 16'h008E; #100;
A = 16'h0095; B = 16'h008F; #100;
A = 16'h0095; B = 16'h0090; #100;
A = 16'h0095; B = 16'h0091; #100;
A = 16'h0095; B = 16'h0092; #100;
A = 16'h0095; B = 16'h0093; #100;
A = 16'h0095; B = 16'h0094; #100;
A = 16'h0095; B = 16'h0095; #100;
A = 16'h0095; B = 16'h0096; #100;
A = 16'h0095; B = 16'h0097; #100;
A = 16'h0095; B = 16'h0098; #100;
A = 16'h0095; B = 16'h0099; #100;
A = 16'h0095; B = 16'h009A; #100;
A = 16'h0095; B = 16'h009B; #100;
A = 16'h0095; B = 16'h009C; #100;
A = 16'h0095; B = 16'h009D; #100;
A = 16'h0095; B = 16'h009E; #100;
A = 16'h0095; B = 16'h009F; #100;
A = 16'h0095; B = 16'h00A0; #100;
A = 16'h0095; B = 16'h00A1; #100;
A = 16'h0095; B = 16'h00A2; #100;
A = 16'h0095; B = 16'h00A3; #100;
A = 16'h0095; B = 16'h00A4; #100;
A = 16'h0095; B = 16'h00A5; #100;
A = 16'h0095; B = 16'h00A6; #100;
A = 16'h0095; B = 16'h00A7; #100;
A = 16'h0095; B = 16'h00A8; #100;
A = 16'h0095; B = 16'h00A9; #100;
A = 16'h0095; B = 16'h00AA; #100;
A = 16'h0095; B = 16'h00AB; #100;
A = 16'h0095; B = 16'h00AC; #100;
A = 16'h0095; B = 16'h00AD; #100;
A = 16'h0095; B = 16'h00AE; #100;
A = 16'h0095; B = 16'h00AF; #100;
A = 16'h0095; B = 16'h00B0; #100;
A = 16'h0095; B = 16'h00B1; #100;
A = 16'h0095; B = 16'h00B2; #100;
A = 16'h0095; B = 16'h00B3; #100;
A = 16'h0095; B = 16'h00B4; #100;
A = 16'h0095; B = 16'h00B5; #100;
A = 16'h0095; B = 16'h00B6; #100;
A = 16'h0095; B = 16'h00B7; #100;
A = 16'h0095; B = 16'h00B8; #100;
A = 16'h0095; B = 16'h00B9; #100;
A = 16'h0095; B = 16'h00BA; #100;
A = 16'h0095; B = 16'h00BB; #100;
A = 16'h0095; B = 16'h00BC; #100;
A = 16'h0095; B = 16'h00BD; #100;
A = 16'h0095; B = 16'h00BE; #100;
A = 16'h0095; B = 16'h00BF; #100;
A = 16'h0095; B = 16'h00C0; #100;
A = 16'h0095; B = 16'h00C1; #100;
A = 16'h0095; B = 16'h00C2; #100;
A = 16'h0095; B = 16'h00C3; #100;
A = 16'h0095; B = 16'h00C4; #100;
A = 16'h0095; B = 16'h00C5; #100;
A = 16'h0095; B = 16'h00C6; #100;
A = 16'h0095; B = 16'h00C7; #100;
A = 16'h0095; B = 16'h00C8; #100;
A = 16'h0095; B = 16'h00C9; #100;
A = 16'h0095; B = 16'h00CA; #100;
A = 16'h0095; B = 16'h00CB; #100;
A = 16'h0095; B = 16'h00CC; #100;
A = 16'h0095; B = 16'h00CD; #100;
A = 16'h0095; B = 16'h00CE; #100;
A = 16'h0095; B = 16'h00CF; #100;
A = 16'h0095; B = 16'h00D0; #100;
A = 16'h0095; B = 16'h00D1; #100;
A = 16'h0095; B = 16'h00D2; #100;
A = 16'h0095; B = 16'h00D3; #100;
A = 16'h0095; B = 16'h00D4; #100;
A = 16'h0095; B = 16'h00D5; #100;
A = 16'h0095; B = 16'h00D6; #100;
A = 16'h0095; B = 16'h00D7; #100;
A = 16'h0095; B = 16'h00D8; #100;
A = 16'h0095; B = 16'h00D9; #100;
A = 16'h0095; B = 16'h00DA; #100;
A = 16'h0095; B = 16'h00DB; #100;
A = 16'h0095; B = 16'h00DC; #100;
A = 16'h0095; B = 16'h00DD; #100;
A = 16'h0095; B = 16'h00DE; #100;
A = 16'h0095; B = 16'h00DF; #100;
A = 16'h0095; B = 16'h00E0; #100;
A = 16'h0095; B = 16'h00E1; #100;
A = 16'h0095; B = 16'h00E2; #100;
A = 16'h0095; B = 16'h00E3; #100;
A = 16'h0095; B = 16'h00E4; #100;
A = 16'h0095; B = 16'h00E5; #100;
A = 16'h0095; B = 16'h00E6; #100;
A = 16'h0095; B = 16'h00E7; #100;
A = 16'h0095; B = 16'h00E8; #100;
A = 16'h0095; B = 16'h00E9; #100;
A = 16'h0095; B = 16'h00EA; #100;
A = 16'h0095; B = 16'h00EB; #100;
A = 16'h0095; B = 16'h00EC; #100;
A = 16'h0095; B = 16'h00ED; #100;
A = 16'h0095; B = 16'h00EE; #100;
A = 16'h0095; B = 16'h00EF; #100;
A = 16'h0095; B = 16'h00F0; #100;
A = 16'h0095; B = 16'h00F1; #100;
A = 16'h0095; B = 16'h00F2; #100;
A = 16'h0095; B = 16'h00F3; #100;
A = 16'h0095; B = 16'h00F4; #100;
A = 16'h0095; B = 16'h00F5; #100;
A = 16'h0095; B = 16'h00F6; #100;
A = 16'h0095; B = 16'h00F7; #100;
A = 16'h0095; B = 16'h00F8; #100;
A = 16'h0095; B = 16'h00F9; #100;
A = 16'h0095; B = 16'h00FA; #100;
A = 16'h0095; B = 16'h00FB; #100;
A = 16'h0095; B = 16'h00FC; #100;
A = 16'h0095; B = 16'h00FD; #100;
A = 16'h0095; B = 16'h00FE; #100;
A = 16'h0095; B = 16'h00FF; #100;
A = 16'h0096; B = 16'h000; #100;
A = 16'h0096; B = 16'h001; #100;
A = 16'h0096; B = 16'h002; #100;
A = 16'h0096; B = 16'h003; #100;
A = 16'h0096; B = 16'h004; #100;
A = 16'h0096; B = 16'h005; #100;
A = 16'h0096; B = 16'h006; #100;
A = 16'h0096; B = 16'h007; #100;
A = 16'h0096; B = 16'h008; #100;
A = 16'h0096; B = 16'h009; #100;
A = 16'h0096; B = 16'h00A; #100;
A = 16'h0096; B = 16'h00B; #100;
A = 16'h0096; B = 16'h00C; #100;
A = 16'h0096; B = 16'h00D; #100;
A = 16'h0096; B = 16'h00E; #100;
A = 16'h0096; B = 16'h00F; #100;
A = 16'h0096; B = 16'h0010; #100;
A = 16'h0096; B = 16'h0011; #100;
A = 16'h0096; B = 16'h0012; #100;
A = 16'h0096; B = 16'h0013; #100;
A = 16'h0096; B = 16'h0014; #100;
A = 16'h0096; B = 16'h0015; #100;
A = 16'h0096; B = 16'h0016; #100;
A = 16'h0096; B = 16'h0017; #100;
A = 16'h0096; B = 16'h0018; #100;
A = 16'h0096; B = 16'h0019; #100;
A = 16'h0096; B = 16'h001A; #100;
A = 16'h0096; B = 16'h001B; #100;
A = 16'h0096; B = 16'h001C; #100;
A = 16'h0096; B = 16'h001D; #100;
A = 16'h0096; B = 16'h001E; #100;
A = 16'h0096; B = 16'h001F; #100;
A = 16'h0096; B = 16'h0020; #100;
A = 16'h0096; B = 16'h0021; #100;
A = 16'h0096; B = 16'h0022; #100;
A = 16'h0096; B = 16'h0023; #100;
A = 16'h0096; B = 16'h0024; #100;
A = 16'h0096; B = 16'h0025; #100;
A = 16'h0096; B = 16'h0026; #100;
A = 16'h0096; B = 16'h0027; #100;
A = 16'h0096; B = 16'h0028; #100;
A = 16'h0096; B = 16'h0029; #100;
A = 16'h0096; B = 16'h002A; #100;
A = 16'h0096; B = 16'h002B; #100;
A = 16'h0096; B = 16'h002C; #100;
A = 16'h0096; B = 16'h002D; #100;
A = 16'h0096; B = 16'h002E; #100;
A = 16'h0096; B = 16'h002F; #100;
A = 16'h0096; B = 16'h0030; #100;
A = 16'h0096; B = 16'h0031; #100;
A = 16'h0096; B = 16'h0032; #100;
A = 16'h0096; B = 16'h0033; #100;
A = 16'h0096; B = 16'h0034; #100;
A = 16'h0096; B = 16'h0035; #100;
A = 16'h0096; B = 16'h0036; #100;
A = 16'h0096; B = 16'h0037; #100;
A = 16'h0096; B = 16'h0038; #100;
A = 16'h0096; B = 16'h0039; #100;
A = 16'h0096; B = 16'h003A; #100;
A = 16'h0096; B = 16'h003B; #100;
A = 16'h0096; B = 16'h003C; #100;
A = 16'h0096; B = 16'h003D; #100;
A = 16'h0096; B = 16'h003E; #100;
A = 16'h0096; B = 16'h003F; #100;
A = 16'h0096; B = 16'h0040; #100;
A = 16'h0096; B = 16'h0041; #100;
A = 16'h0096; B = 16'h0042; #100;
A = 16'h0096; B = 16'h0043; #100;
A = 16'h0096; B = 16'h0044; #100;
A = 16'h0096; B = 16'h0045; #100;
A = 16'h0096; B = 16'h0046; #100;
A = 16'h0096; B = 16'h0047; #100;
A = 16'h0096; B = 16'h0048; #100;
A = 16'h0096; B = 16'h0049; #100;
A = 16'h0096; B = 16'h004A; #100;
A = 16'h0096; B = 16'h004B; #100;
A = 16'h0096; B = 16'h004C; #100;
A = 16'h0096; B = 16'h004D; #100;
A = 16'h0096; B = 16'h004E; #100;
A = 16'h0096; B = 16'h004F; #100;
A = 16'h0096; B = 16'h0050; #100;
A = 16'h0096; B = 16'h0051; #100;
A = 16'h0096; B = 16'h0052; #100;
A = 16'h0096; B = 16'h0053; #100;
A = 16'h0096; B = 16'h0054; #100;
A = 16'h0096; B = 16'h0055; #100;
A = 16'h0096; B = 16'h0056; #100;
A = 16'h0096; B = 16'h0057; #100;
A = 16'h0096; B = 16'h0058; #100;
A = 16'h0096; B = 16'h0059; #100;
A = 16'h0096; B = 16'h005A; #100;
A = 16'h0096; B = 16'h005B; #100;
A = 16'h0096; B = 16'h005C; #100;
A = 16'h0096; B = 16'h005D; #100;
A = 16'h0096; B = 16'h005E; #100;
A = 16'h0096; B = 16'h005F; #100;
A = 16'h0096; B = 16'h0060; #100;
A = 16'h0096; B = 16'h0061; #100;
A = 16'h0096; B = 16'h0062; #100;
A = 16'h0096; B = 16'h0063; #100;
A = 16'h0096; B = 16'h0064; #100;
A = 16'h0096; B = 16'h0065; #100;
A = 16'h0096; B = 16'h0066; #100;
A = 16'h0096; B = 16'h0067; #100;
A = 16'h0096; B = 16'h0068; #100;
A = 16'h0096; B = 16'h0069; #100;
A = 16'h0096; B = 16'h006A; #100;
A = 16'h0096; B = 16'h006B; #100;
A = 16'h0096; B = 16'h006C; #100;
A = 16'h0096; B = 16'h006D; #100;
A = 16'h0096; B = 16'h006E; #100;
A = 16'h0096; B = 16'h006F; #100;
A = 16'h0096; B = 16'h0070; #100;
A = 16'h0096; B = 16'h0071; #100;
A = 16'h0096; B = 16'h0072; #100;
A = 16'h0096; B = 16'h0073; #100;
A = 16'h0096; B = 16'h0074; #100;
A = 16'h0096; B = 16'h0075; #100;
A = 16'h0096; B = 16'h0076; #100;
A = 16'h0096; B = 16'h0077; #100;
A = 16'h0096; B = 16'h0078; #100;
A = 16'h0096; B = 16'h0079; #100;
A = 16'h0096; B = 16'h007A; #100;
A = 16'h0096; B = 16'h007B; #100;
A = 16'h0096; B = 16'h007C; #100;
A = 16'h0096; B = 16'h007D; #100;
A = 16'h0096; B = 16'h007E; #100;
A = 16'h0096; B = 16'h007F; #100;
A = 16'h0096; B = 16'h0080; #100;
A = 16'h0096; B = 16'h0081; #100;
A = 16'h0096; B = 16'h0082; #100;
A = 16'h0096; B = 16'h0083; #100;
A = 16'h0096; B = 16'h0084; #100;
A = 16'h0096; B = 16'h0085; #100;
A = 16'h0096; B = 16'h0086; #100;
A = 16'h0096; B = 16'h0087; #100;
A = 16'h0096; B = 16'h0088; #100;
A = 16'h0096; B = 16'h0089; #100;
A = 16'h0096; B = 16'h008A; #100;
A = 16'h0096; B = 16'h008B; #100;
A = 16'h0096; B = 16'h008C; #100;
A = 16'h0096; B = 16'h008D; #100;
A = 16'h0096; B = 16'h008E; #100;
A = 16'h0096; B = 16'h008F; #100;
A = 16'h0096; B = 16'h0090; #100;
A = 16'h0096; B = 16'h0091; #100;
A = 16'h0096; B = 16'h0092; #100;
A = 16'h0096; B = 16'h0093; #100;
A = 16'h0096; B = 16'h0094; #100;
A = 16'h0096; B = 16'h0095; #100;
A = 16'h0096; B = 16'h0096; #100;
A = 16'h0096; B = 16'h0097; #100;
A = 16'h0096; B = 16'h0098; #100;
A = 16'h0096; B = 16'h0099; #100;
A = 16'h0096; B = 16'h009A; #100;
A = 16'h0096; B = 16'h009B; #100;
A = 16'h0096; B = 16'h009C; #100;
A = 16'h0096; B = 16'h009D; #100;
A = 16'h0096; B = 16'h009E; #100;
A = 16'h0096; B = 16'h009F; #100;
A = 16'h0096; B = 16'h00A0; #100;
A = 16'h0096; B = 16'h00A1; #100;
A = 16'h0096; B = 16'h00A2; #100;
A = 16'h0096; B = 16'h00A3; #100;
A = 16'h0096; B = 16'h00A4; #100;
A = 16'h0096; B = 16'h00A5; #100;
A = 16'h0096; B = 16'h00A6; #100;
A = 16'h0096; B = 16'h00A7; #100;
A = 16'h0096; B = 16'h00A8; #100;
A = 16'h0096; B = 16'h00A9; #100;
A = 16'h0096; B = 16'h00AA; #100;
A = 16'h0096; B = 16'h00AB; #100;
A = 16'h0096; B = 16'h00AC; #100;
A = 16'h0096; B = 16'h00AD; #100;
A = 16'h0096; B = 16'h00AE; #100;
A = 16'h0096; B = 16'h00AF; #100;
A = 16'h0096; B = 16'h00B0; #100;
A = 16'h0096; B = 16'h00B1; #100;
A = 16'h0096; B = 16'h00B2; #100;
A = 16'h0096; B = 16'h00B3; #100;
A = 16'h0096; B = 16'h00B4; #100;
A = 16'h0096; B = 16'h00B5; #100;
A = 16'h0096; B = 16'h00B6; #100;
A = 16'h0096; B = 16'h00B7; #100;
A = 16'h0096; B = 16'h00B8; #100;
A = 16'h0096; B = 16'h00B9; #100;
A = 16'h0096; B = 16'h00BA; #100;
A = 16'h0096; B = 16'h00BB; #100;
A = 16'h0096; B = 16'h00BC; #100;
A = 16'h0096; B = 16'h00BD; #100;
A = 16'h0096; B = 16'h00BE; #100;
A = 16'h0096; B = 16'h00BF; #100;
A = 16'h0096; B = 16'h00C0; #100;
A = 16'h0096; B = 16'h00C1; #100;
A = 16'h0096; B = 16'h00C2; #100;
A = 16'h0096; B = 16'h00C3; #100;
A = 16'h0096; B = 16'h00C4; #100;
A = 16'h0096; B = 16'h00C5; #100;
A = 16'h0096; B = 16'h00C6; #100;
A = 16'h0096; B = 16'h00C7; #100;
A = 16'h0096; B = 16'h00C8; #100;
A = 16'h0096; B = 16'h00C9; #100;
A = 16'h0096; B = 16'h00CA; #100;
A = 16'h0096; B = 16'h00CB; #100;
A = 16'h0096; B = 16'h00CC; #100;
A = 16'h0096; B = 16'h00CD; #100;
A = 16'h0096; B = 16'h00CE; #100;
A = 16'h0096; B = 16'h00CF; #100;
A = 16'h0096; B = 16'h00D0; #100;
A = 16'h0096; B = 16'h00D1; #100;
A = 16'h0096; B = 16'h00D2; #100;
A = 16'h0096; B = 16'h00D3; #100;
A = 16'h0096; B = 16'h00D4; #100;
A = 16'h0096; B = 16'h00D5; #100;
A = 16'h0096; B = 16'h00D6; #100;
A = 16'h0096; B = 16'h00D7; #100;
A = 16'h0096; B = 16'h00D8; #100;
A = 16'h0096; B = 16'h00D9; #100;
A = 16'h0096; B = 16'h00DA; #100;
A = 16'h0096; B = 16'h00DB; #100;
A = 16'h0096; B = 16'h00DC; #100;
A = 16'h0096; B = 16'h00DD; #100;
A = 16'h0096; B = 16'h00DE; #100;
A = 16'h0096; B = 16'h00DF; #100;
A = 16'h0096; B = 16'h00E0; #100;
A = 16'h0096; B = 16'h00E1; #100;
A = 16'h0096; B = 16'h00E2; #100;
A = 16'h0096; B = 16'h00E3; #100;
A = 16'h0096; B = 16'h00E4; #100;
A = 16'h0096; B = 16'h00E5; #100;
A = 16'h0096; B = 16'h00E6; #100;
A = 16'h0096; B = 16'h00E7; #100;
A = 16'h0096; B = 16'h00E8; #100;
A = 16'h0096; B = 16'h00E9; #100;
A = 16'h0096; B = 16'h00EA; #100;
A = 16'h0096; B = 16'h00EB; #100;
A = 16'h0096; B = 16'h00EC; #100;
A = 16'h0096; B = 16'h00ED; #100;
A = 16'h0096; B = 16'h00EE; #100;
A = 16'h0096; B = 16'h00EF; #100;
A = 16'h0096; B = 16'h00F0; #100;
A = 16'h0096; B = 16'h00F1; #100;
A = 16'h0096; B = 16'h00F2; #100;
A = 16'h0096; B = 16'h00F3; #100;
A = 16'h0096; B = 16'h00F4; #100;
A = 16'h0096; B = 16'h00F5; #100;
A = 16'h0096; B = 16'h00F6; #100;
A = 16'h0096; B = 16'h00F7; #100;
A = 16'h0096; B = 16'h00F8; #100;
A = 16'h0096; B = 16'h00F9; #100;
A = 16'h0096; B = 16'h00FA; #100;
A = 16'h0096; B = 16'h00FB; #100;
A = 16'h0096; B = 16'h00FC; #100;
A = 16'h0096; B = 16'h00FD; #100;
A = 16'h0096; B = 16'h00FE; #100;
A = 16'h0096; B = 16'h00FF; #100;
A = 16'h0097; B = 16'h000; #100;
A = 16'h0097; B = 16'h001; #100;
A = 16'h0097; B = 16'h002; #100;
A = 16'h0097; B = 16'h003; #100;
A = 16'h0097; B = 16'h004; #100;
A = 16'h0097; B = 16'h005; #100;
A = 16'h0097; B = 16'h006; #100;
A = 16'h0097; B = 16'h007; #100;
A = 16'h0097; B = 16'h008; #100;
A = 16'h0097; B = 16'h009; #100;
A = 16'h0097; B = 16'h00A; #100;
A = 16'h0097; B = 16'h00B; #100;
A = 16'h0097; B = 16'h00C; #100;
A = 16'h0097; B = 16'h00D; #100;
A = 16'h0097; B = 16'h00E; #100;
A = 16'h0097; B = 16'h00F; #100;
A = 16'h0097; B = 16'h0010; #100;
A = 16'h0097; B = 16'h0011; #100;
A = 16'h0097; B = 16'h0012; #100;
A = 16'h0097; B = 16'h0013; #100;
A = 16'h0097; B = 16'h0014; #100;
A = 16'h0097; B = 16'h0015; #100;
A = 16'h0097; B = 16'h0016; #100;
A = 16'h0097; B = 16'h0017; #100;
A = 16'h0097; B = 16'h0018; #100;
A = 16'h0097; B = 16'h0019; #100;
A = 16'h0097; B = 16'h001A; #100;
A = 16'h0097; B = 16'h001B; #100;
A = 16'h0097; B = 16'h001C; #100;
A = 16'h0097; B = 16'h001D; #100;
A = 16'h0097; B = 16'h001E; #100;
A = 16'h0097; B = 16'h001F; #100;
A = 16'h0097; B = 16'h0020; #100;
A = 16'h0097; B = 16'h0021; #100;
A = 16'h0097; B = 16'h0022; #100;
A = 16'h0097; B = 16'h0023; #100;
A = 16'h0097; B = 16'h0024; #100;
A = 16'h0097; B = 16'h0025; #100;
A = 16'h0097; B = 16'h0026; #100;
A = 16'h0097; B = 16'h0027; #100;
A = 16'h0097; B = 16'h0028; #100;
A = 16'h0097; B = 16'h0029; #100;
A = 16'h0097; B = 16'h002A; #100;
A = 16'h0097; B = 16'h002B; #100;
A = 16'h0097; B = 16'h002C; #100;
A = 16'h0097; B = 16'h002D; #100;
A = 16'h0097; B = 16'h002E; #100;
A = 16'h0097; B = 16'h002F; #100;
A = 16'h0097; B = 16'h0030; #100;
A = 16'h0097; B = 16'h0031; #100;
A = 16'h0097; B = 16'h0032; #100;
A = 16'h0097; B = 16'h0033; #100;
A = 16'h0097; B = 16'h0034; #100;
A = 16'h0097; B = 16'h0035; #100;
A = 16'h0097; B = 16'h0036; #100;
A = 16'h0097; B = 16'h0037; #100;
A = 16'h0097; B = 16'h0038; #100;
A = 16'h0097; B = 16'h0039; #100;
A = 16'h0097; B = 16'h003A; #100;
A = 16'h0097; B = 16'h003B; #100;
A = 16'h0097; B = 16'h003C; #100;
A = 16'h0097; B = 16'h003D; #100;
A = 16'h0097; B = 16'h003E; #100;
A = 16'h0097; B = 16'h003F; #100;
A = 16'h0097; B = 16'h0040; #100;
A = 16'h0097; B = 16'h0041; #100;
A = 16'h0097; B = 16'h0042; #100;
A = 16'h0097; B = 16'h0043; #100;
A = 16'h0097; B = 16'h0044; #100;
A = 16'h0097; B = 16'h0045; #100;
A = 16'h0097; B = 16'h0046; #100;
A = 16'h0097; B = 16'h0047; #100;
A = 16'h0097; B = 16'h0048; #100;
A = 16'h0097; B = 16'h0049; #100;
A = 16'h0097; B = 16'h004A; #100;
A = 16'h0097; B = 16'h004B; #100;
A = 16'h0097; B = 16'h004C; #100;
A = 16'h0097; B = 16'h004D; #100;
A = 16'h0097; B = 16'h004E; #100;
A = 16'h0097; B = 16'h004F; #100;
A = 16'h0097; B = 16'h0050; #100;
A = 16'h0097; B = 16'h0051; #100;
A = 16'h0097; B = 16'h0052; #100;
A = 16'h0097; B = 16'h0053; #100;
A = 16'h0097; B = 16'h0054; #100;
A = 16'h0097; B = 16'h0055; #100;
A = 16'h0097; B = 16'h0056; #100;
A = 16'h0097; B = 16'h0057; #100;
A = 16'h0097; B = 16'h0058; #100;
A = 16'h0097; B = 16'h0059; #100;
A = 16'h0097; B = 16'h005A; #100;
A = 16'h0097; B = 16'h005B; #100;
A = 16'h0097; B = 16'h005C; #100;
A = 16'h0097; B = 16'h005D; #100;
A = 16'h0097; B = 16'h005E; #100;
A = 16'h0097; B = 16'h005F; #100;
A = 16'h0097; B = 16'h0060; #100;
A = 16'h0097; B = 16'h0061; #100;
A = 16'h0097; B = 16'h0062; #100;
A = 16'h0097; B = 16'h0063; #100;
A = 16'h0097; B = 16'h0064; #100;
A = 16'h0097; B = 16'h0065; #100;
A = 16'h0097; B = 16'h0066; #100;
A = 16'h0097; B = 16'h0067; #100;
A = 16'h0097; B = 16'h0068; #100;
A = 16'h0097; B = 16'h0069; #100;
A = 16'h0097; B = 16'h006A; #100;
A = 16'h0097; B = 16'h006B; #100;
A = 16'h0097; B = 16'h006C; #100;
A = 16'h0097; B = 16'h006D; #100;
A = 16'h0097; B = 16'h006E; #100;
A = 16'h0097; B = 16'h006F; #100;
A = 16'h0097; B = 16'h0070; #100;
A = 16'h0097; B = 16'h0071; #100;
A = 16'h0097; B = 16'h0072; #100;
A = 16'h0097; B = 16'h0073; #100;
A = 16'h0097; B = 16'h0074; #100;
A = 16'h0097; B = 16'h0075; #100;
A = 16'h0097; B = 16'h0076; #100;
A = 16'h0097; B = 16'h0077; #100;
A = 16'h0097; B = 16'h0078; #100;
A = 16'h0097; B = 16'h0079; #100;
A = 16'h0097; B = 16'h007A; #100;
A = 16'h0097; B = 16'h007B; #100;
A = 16'h0097; B = 16'h007C; #100;
A = 16'h0097; B = 16'h007D; #100;
A = 16'h0097; B = 16'h007E; #100;
A = 16'h0097; B = 16'h007F; #100;
A = 16'h0097; B = 16'h0080; #100;
A = 16'h0097; B = 16'h0081; #100;
A = 16'h0097; B = 16'h0082; #100;
A = 16'h0097; B = 16'h0083; #100;
A = 16'h0097; B = 16'h0084; #100;
A = 16'h0097; B = 16'h0085; #100;
A = 16'h0097; B = 16'h0086; #100;
A = 16'h0097; B = 16'h0087; #100;
A = 16'h0097; B = 16'h0088; #100;
A = 16'h0097; B = 16'h0089; #100;
A = 16'h0097; B = 16'h008A; #100;
A = 16'h0097; B = 16'h008B; #100;
A = 16'h0097; B = 16'h008C; #100;
A = 16'h0097; B = 16'h008D; #100;
A = 16'h0097; B = 16'h008E; #100;
A = 16'h0097; B = 16'h008F; #100;
A = 16'h0097; B = 16'h0090; #100;
A = 16'h0097; B = 16'h0091; #100;
A = 16'h0097; B = 16'h0092; #100;
A = 16'h0097; B = 16'h0093; #100;
A = 16'h0097; B = 16'h0094; #100;
A = 16'h0097; B = 16'h0095; #100;
A = 16'h0097; B = 16'h0096; #100;
A = 16'h0097; B = 16'h0097; #100;
A = 16'h0097; B = 16'h0098; #100;
A = 16'h0097; B = 16'h0099; #100;
A = 16'h0097; B = 16'h009A; #100;
A = 16'h0097; B = 16'h009B; #100;
A = 16'h0097; B = 16'h009C; #100;
A = 16'h0097; B = 16'h009D; #100;
A = 16'h0097; B = 16'h009E; #100;
A = 16'h0097; B = 16'h009F; #100;
A = 16'h0097; B = 16'h00A0; #100;
A = 16'h0097; B = 16'h00A1; #100;
A = 16'h0097; B = 16'h00A2; #100;
A = 16'h0097; B = 16'h00A3; #100;
A = 16'h0097; B = 16'h00A4; #100;
A = 16'h0097; B = 16'h00A5; #100;
A = 16'h0097; B = 16'h00A6; #100;
A = 16'h0097; B = 16'h00A7; #100;
A = 16'h0097; B = 16'h00A8; #100;
A = 16'h0097; B = 16'h00A9; #100;
A = 16'h0097; B = 16'h00AA; #100;
A = 16'h0097; B = 16'h00AB; #100;
A = 16'h0097; B = 16'h00AC; #100;
A = 16'h0097; B = 16'h00AD; #100;
A = 16'h0097; B = 16'h00AE; #100;
A = 16'h0097; B = 16'h00AF; #100;
A = 16'h0097; B = 16'h00B0; #100;
A = 16'h0097; B = 16'h00B1; #100;
A = 16'h0097; B = 16'h00B2; #100;
A = 16'h0097; B = 16'h00B3; #100;
A = 16'h0097; B = 16'h00B4; #100;
A = 16'h0097; B = 16'h00B5; #100;
A = 16'h0097; B = 16'h00B6; #100;
A = 16'h0097; B = 16'h00B7; #100;
A = 16'h0097; B = 16'h00B8; #100;
A = 16'h0097; B = 16'h00B9; #100;
A = 16'h0097; B = 16'h00BA; #100;
A = 16'h0097; B = 16'h00BB; #100;
A = 16'h0097; B = 16'h00BC; #100;
A = 16'h0097; B = 16'h00BD; #100;
A = 16'h0097; B = 16'h00BE; #100;
A = 16'h0097; B = 16'h00BF; #100;
A = 16'h0097; B = 16'h00C0; #100;
A = 16'h0097; B = 16'h00C1; #100;
A = 16'h0097; B = 16'h00C2; #100;
A = 16'h0097; B = 16'h00C3; #100;
A = 16'h0097; B = 16'h00C4; #100;
A = 16'h0097; B = 16'h00C5; #100;
A = 16'h0097; B = 16'h00C6; #100;
A = 16'h0097; B = 16'h00C7; #100;
A = 16'h0097; B = 16'h00C8; #100;
A = 16'h0097; B = 16'h00C9; #100;
A = 16'h0097; B = 16'h00CA; #100;
A = 16'h0097; B = 16'h00CB; #100;
A = 16'h0097; B = 16'h00CC; #100;
A = 16'h0097; B = 16'h00CD; #100;
A = 16'h0097; B = 16'h00CE; #100;
A = 16'h0097; B = 16'h00CF; #100;
A = 16'h0097; B = 16'h00D0; #100;
A = 16'h0097; B = 16'h00D1; #100;
A = 16'h0097; B = 16'h00D2; #100;
A = 16'h0097; B = 16'h00D3; #100;
A = 16'h0097; B = 16'h00D4; #100;
A = 16'h0097; B = 16'h00D5; #100;
A = 16'h0097; B = 16'h00D6; #100;
A = 16'h0097; B = 16'h00D7; #100;
A = 16'h0097; B = 16'h00D8; #100;
A = 16'h0097; B = 16'h00D9; #100;
A = 16'h0097; B = 16'h00DA; #100;
A = 16'h0097; B = 16'h00DB; #100;
A = 16'h0097; B = 16'h00DC; #100;
A = 16'h0097; B = 16'h00DD; #100;
A = 16'h0097; B = 16'h00DE; #100;
A = 16'h0097; B = 16'h00DF; #100;
A = 16'h0097; B = 16'h00E0; #100;
A = 16'h0097; B = 16'h00E1; #100;
A = 16'h0097; B = 16'h00E2; #100;
A = 16'h0097; B = 16'h00E3; #100;
A = 16'h0097; B = 16'h00E4; #100;
A = 16'h0097; B = 16'h00E5; #100;
A = 16'h0097; B = 16'h00E6; #100;
A = 16'h0097; B = 16'h00E7; #100;
A = 16'h0097; B = 16'h00E8; #100;
A = 16'h0097; B = 16'h00E9; #100;
A = 16'h0097; B = 16'h00EA; #100;
A = 16'h0097; B = 16'h00EB; #100;
A = 16'h0097; B = 16'h00EC; #100;
A = 16'h0097; B = 16'h00ED; #100;
A = 16'h0097; B = 16'h00EE; #100;
A = 16'h0097; B = 16'h00EF; #100;
A = 16'h0097; B = 16'h00F0; #100;
A = 16'h0097; B = 16'h00F1; #100;
A = 16'h0097; B = 16'h00F2; #100;
A = 16'h0097; B = 16'h00F3; #100;
A = 16'h0097; B = 16'h00F4; #100;
A = 16'h0097; B = 16'h00F5; #100;
A = 16'h0097; B = 16'h00F6; #100;
A = 16'h0097; B = 16'h00F7; #100;
A = 16'h0097; B = 16'h00F8; #100;
A = 16'h0097; B = 16'h00F9; #100;
A = 16'h0097; B = 16'h00FA; #100;
A = 16'h0097; B = 16'h00FB; #100;
A = 16'h0097; B = 16'h00FC; #100;
A = 16'h0097; B = 16'h00FD; #100;
A = 16'h0097; B = 16'h00FE; #100;
A = 16'h0097; B = 16'h00FF; #100;
A = 16'h0098; B = 16'h000; #100;
A = 16'h0098; B = 16'h001; #100;
A = 16'h0098; B = 16'h002; #100;
A = 16'h0098; B = 16'h003; #100;
A = 16'h0098; B = 16'h004; #100;
A = 16'h0098; B = 16'h005; #100;
A = 16'h0098; B = 16'h006; #100;
A = 16'h0098; B = 16'h007; #100;
A = 16'h0098; B = 16'h008; #100;
A = 16'h0098; B = 16'h009; #100;
A = 16'h0098; B = 16'h00A; #100;
A = 16'h0098; B = 16'h00B; #100;
A = 16'h0098; B = 16'h00C; #100;
A = 16'h0098; B = 16'h00D; #100;
A = 16'h0098; B = 16'h00E; #100;
A = 16'h0098; B = 16'h00F; #100;
A = 16'h0098; B = 16'h0010; #100;
A = 16'h0098; B = 16'h0011; #100;
A = 16'h0098; B = 16'h0012; #100;
A = 16'h0098; B = 16'h0013; #100;
A = 16'h0098; B = 16'h0014; #100;
A = 16'h0098; B = 16'h0015; #100;
A = 16'h0098; B = 16'h0016; #100;
A = 16'h0098; B = 16'h0017; #100;
A = 16'h0098; B = 16'h0018; #100;
A = 16'h0098; B = 16'h0019; #100;
A = 16'h0098; B = 16'h001A; #100;
A = 16'h0098; B = 16'h001B; #100;
A = 16'h0098; B = 16'h001C; #100;
A = 16'h0098; B = 16'h001D; #100;
A = 16'h0098; B = 16'h001E; #100;
A = 16'h0098; B = 16'h001F; #100;
A = 16'h0098; B = 16'h0020; #100;
A = 16'h0098; B = 16'h0021; #100;
A = 16'h0098; B = 16'h0022; #100;
A = 16'h0098; B = 16'h0023; #100;
A = 16'h0098; B = 16'h0024; #100;
A = 16'h0098; B = 16'h0025; #100;
A = 16'h0098; B = 16'h0026; #100;
A = 16'h0098; B = 16'h0027; #100;
A = 16'h0098; B = 16'h0028; #100;
A = 16'h0098; B = 16'h0029; #100;
A = 16'h0098; B = 16'h002A; #100;
A = 16'h0098; B = 16'h002B; #100;
A = 16'h0098; B = 16'h002C; #100;
A = 16'h0098; B = 16'h002D; #100;
A = 16'h0098; B = 16'h002E; #100;
A = 16'h0098; B = 16'h002F; #100;
A = 16'h0098; B = 16'h0030; #100;
A = 16'h0098; B = 16'h0031; #100;
A = 16'h0098; B = 16'h0032; #100;
A = 16'h0098; B = 16'h0033; #100;
A = 16'h0098; B = 16'h0034; #100;
A = 16'h0098; B = 16'h0035; #100;
A = 16'h0098; B = 16'h0036; #100;
A = 16'h0098; B = 16'h0037; #100;
A = 16'h0098; B = 16'h0038; #100;
A = 16'h0098; B = 16'h0039; #100;
A = 16'h0098; B = 16'h003A; #100;
A = 16'h0098; B = 16'h003B; #100;
A = 16'h0098; B = 16'h003C; #100;
A = 16'h0098; B = 16'h003D; #100;
A = 16'h0098; B = 16'h003E; #100;
A = 16'h0098; B = 16'h003F; #100;
A = 16'h0098; B = 16'h0040; #100;
A = 16'h0098; B = 16'h0041; #100;
A = 16'h0098; B = 16'h0042; #100;
A = 16'h0098; B = 16'h0043; #100;
A = 16'h0098; B = 16'h0044; #100;
A = 16'h0098; B = 16'h0045; #100;
A = 16'h0098; B = 16'h0046; #100;
A = 16'h0098; B = 16'h0047; #100;
A = 16'h0098; B = 16'h0048; #100;
A = 16'h0098; B = 16'h0049; #100;
A = 16'h0098; B = 16'h004A; #100;
A = 16'h0098; B = 16'h004B; #100;
A = 16'h0098; B = 16'h004C; #100;
A = 16'h0098; B = 16'h004D; #100;
A = 16'h0098; B = 16'h004E; #100;
A = 16'h0098; B = 16'h004F; #100;
A = 16'h0098; B = 16'h0050; #100;
A = 16'h0098; B = 16'h0051; #100;
A = 16'h0098; B = 16'h0052; #100;
A = 16'h0098; B = 16'h0053; #100;
A = 16'h0098; B = 16'h0054; #100;
A = 16'h0098; B = 16'h0055; #100;
A = 16'h0098; B = 16'h0056; #100;
A = 16'h0098; B = 16'h0057; #100;
A = 16'h0098; B = 16'h0058; #100;
A = 16'h0098; B = 16'h0059; #100;
A = 16'h0098; B = 16'h005A; #100;
A = 16'h0098; B = 16'h005B; #100;
A = 16'h0098; B = 16'h005C; #100;
A = 16'h0098; B = 16'h005D; #100;
A = 16'h0098; B = 16'h005E; #100;
A = 16'h0098; B = 16'h005F; #100;
A = 16'h0098; B = 16'h0060; #100;
A = 16'h0098; B = 16'h0061; #100;
A = 16'h0098; B = 16'h0062; #100;
A = 16'h0098; B = 16'h0063; #100;
A = 16'h0098; B = 16'h0064; #100;
A = 16'h0098; B = 16'h0065; #100;
A = 16'h0098; B = 16'h0066; #100;
A = 16'h0098; B = 16'h0067; #100;
A = 16'h0098; B = 16'h0068; #100;
A = 16'h0098; B = 16'h0069; #100;
A = 16'h0098; B = 16'h006A; #100;
A = 16'h0098; B = 16'h006B; #100;
A = 16'h0098; B = 16'h006C; #100;
A = 16'h0098; B = 16'h006D; #100;
A = 16'h0098; B = 16'h006E; #100;
A = 16'h0098; B = 16'h006F; #100;
A = 16'h0098; B = 16'h0070; #100;
A = 16'h0098; B = 16'h0071; #100;
A = 16'h0098; B = 16'h0072; #100;
A = 16'h0098; B = 16'h0073; #100;
A = 16'h0098; B = 16'h0074; #100;
A = 16'h0098; B = 16'h0075; #100;
A = 16'h0098; B = 16'h0076; #100;
A = 16'h0098; B = 16'h0077; #100;
A = 16'h0098; B = 16'h0078; #100;
A = 16'h0098; B = 16'h0079; #100;
A = 16'h0098; B = 16'h007A; #100;
A = 16'h0098; B = 16'h007B; #100;
A = 16'h0098; B = 16'h007C; #100;
A = 16'h0098; B = 16'h007D; #100;
A = 16'h0098; B = 16'h007E; #100;
A = 16'h0098; B = 16'h007F; #100;
A = 16'h0098; B = 16'h0080; #100;
A = 16'h0098; B = 16'h0081; #100;
A = 16'h0098; B = 16'h0082; #100;
A = 16'h0098; B = 16'h0083; #100;
A = 16'h0098; B = 16'h0084; #100;
A = 16'h0098; B = 16'h0085; #100;
A = 16'h0098; B = 16'h0086; #100;
A = 16'h0098; B = 16'h0087; #100;
A = 16'h0098; B = 16'h0088; #100;
A = 16'h0098; B = 16'h0089; #100;
A = 16'h0098; B = 16'h008A; #100;
A = 16'h0098; B = 16'h008B; #100;
A = 16'h0098; B = 16'h008C; #100;
A = 16'h0098; B = 16'h008D; #100;
A = 16'h0098; B = 16'h008E; #100;
A = 16'h0098; B = 16'h008F; #100;
A = 16'h0098; B = 16'h0090; #100;
A = 16'h0098; B = 16'h0091; #100;
A = 16'h0098; B = 16'h0092; #100;
A = 16'h0098; B = 16'h0093; #100;
A = 16'h0098; B = 16'h0094; #100;
A = 16'h0098; B = 16'h0095; #100;
A = 16'h0098; B = 16'h0096; #100;
A = 16'h0098; B = 16'h0097; #100;
A = 16'h0098; B = 16'h0098; #100;
A = 16'h0098; B = 16'h0099; #100;
A = 16'h0098; B = 16'h009A; #100;
A = 16'h0098; B = 16'h009B; #100;
A = 16'h0098; B = 16'h009C; #100;
A = 16'h0098; B = 16'h009D; #100;
A = 16'h0098; B = 16'h009E; #100;
A = 16'h0098; B = 16'h009F; #100;
A = 16'h0098; B = 16'h00A0; #100;
A = 16'h0098; B = 16'h00A1; #100;
A = 16'h0098; B = 16'h00A2; #100;
A = 16'h0098; B = 16'h00A3; #100;
A = 16'h0098; B = 16'h00A4; #100;
A = 16'h0098; B = 16'h00A5; #100;
A = 16'h0098; B = 16'h00A6; #100;
A = 16'h0098; B = 16'h00A7; #100;
A = 16'h0098; B = 16'h00A8; #100;
A = 16'h0098; B = 16'h00A9; #100;
A = 16'h0098; B = 16'h00AA; #100;
A = 16'h0098; B = 16'h00AB; #100;
A = 16'h0098; B = 16'h00AC; #100;
A = 16'h0098; B = 16'h00AD; #100;
A = 16'h0098; B = 16'h00AE; #100;
A = 16'h0098; B = 16'h00AF; #100;
A = 16'h0098; B = 16'h00B0; #100;
A = 16'h0098; B = 16'h00B1; #100;
A = 16'h0098; B = 16'h00B2; #100;
A = 16'h0098; B = 16'h00B3; #100;
A = 16'h0098; B = 16'h00B4; #100;
A = 16'h0098; B = 16'h00B5; #100;
A = 16'h0098; B = 16'h00B6; #100;
A = 16'h0098; B = 16'h00B7; #100;
A = 16'h0098; B = 16'h00B8; #100;
A = 16'h0098; B = 16'h00B9; #100;
A = 16'h0098; B = 16'h00BA; #100;
A = 16'h0098; B = 16'h00BB; #100;
A = 16'h0098; B = 16'h00BC; #100;
A = 16'h0098; B = 16'h00BD; #100;
A = 16'h0098; B = 16'h00BE; #100;
A = 16'h0098; B = 16'h00BF; #100;
A = 16'h0098; B = 16'h00C0; #100;
A = 16'h0098; B = 16'h00C1; #100;
A = 16'h0098; B = 16'h00C2; #100;
A = 16'h0098; B = 16'h00C3; #100;
A = 16'h0098; B = 16'h00C4; #100;
A = 16'h0098; B = 16'h00C5; #100;
A = 16'h0098; B = 16'h00C6; #100;
A = 16'h0098; B = 16'h00C7; #100;
A = 16'h0098; B = 16'h00C8; #100;
A = 16'h0098; B = 16'h00C9; #100;
A = 16'h0098; B = 16'h00CA; #100;
A = 16'h0098; B = 16'h00CB; #100;
A = 16'h0098; B = 16'h00CC; #100;
A = 16'h0098; B = 16'h00CD; #100;
A = 16'h0098; B = 16'h00CE; #100;
A = 16'h0098; B = 16'h00CF; #100;
A = 16'h0098; B = 16'h00D0; #100;
A = 16'h0098; B = 16'h00D1; #100;
A = 16'h0098; B = 16'h00D2; #100;
A = 16'h0098; B = 16'h00D3; #100;
A = 16'h0098; B = 16'h00D4; #100;
A = 16'h0098; B = 16'h00D5; #100;
A = 16'h0098; B = 16'h00D6; #100;
A = 16'h0098; B = 16'h00D7; #100;
A = 16'h0098; B = 16'h00D8; #100;
A = 16'h0098; B = 16'h00D9; #100;
A = 16'h0098; B = 16'h00DA; #100;
A = 16'h0098; B = 16'h00DB; #100;
A = 16'h0098; B = 16'h00DC; #100;
A = 16'h0098; B = 16'h00DD; #100;
A = 16'h0098; B = 16'h00DE; #100;
A = 16'h0098; B = 16'h00DF; #100;
A = 16'h0098; B = 16'h00E0; #100;
A = 16'h0098; B = 16'h00E1; #100;
A = 16'h0098; B = 16'h00E2; #100;
A = 16'h0098; B = 16'h00E3; #100;
A = 16'h0098; B = 16'h00E4; #100;
A = 16'h0098; B = 16'h00E5; #100;
A = 16'h0098; B = 16'h00E6; #100;
A = 16'h0098; B = 16'h00E7; #100;
A = 16'h0098; B = 16'h00E8; #100;
A = 16'h0098; B = 16'h00E9; #100;
A = 16'h0098; B = 16'h00EA; #100;
A = 16'h0098; B = 16'h00EB; #100;
A = 16'h0098; B = 16'h00EC; #100;
A = 16'h0098; B = 16'h00ED; #100;
A = 16'h0098; B = 16'h00EE; #100;
A = 16'h0098; B = 16'h00EF; #100;
A = 16'h0098; B = 16'h00F0; #100;
A = 16'h0098; B = 16'h00F1; #100;
A = 16'h0098; B = 16'h00F2; #100;
A = 16'h0098; B = 16'h00F3; #100;
A = 16'h0098; B = 16'h00F4; #100;
A = 16'h0098; B = 16'h00F5; #100;
A = 16'h0098; B = 16'h00F6; #100;
A = 16'h0098; B = 16'h00F7; #100;
A = 16'h0098; B = 16'h00F8; #100;
A = 16'h0098; B = 16'h00F9; #100;
A = 16'h0098; B = 16'h00FA; #100;
A = 16'h0098; B = 16'h00FB; #100;
A = 16'h0098; B = 16'h00FC; #100;
A = 16'h0098; B = 16'h00FD; #100;
A = 16'h0098; B = 16'h00FE; #100;
A = 16'h0098; B = 16'h00FF; #100;
A = 16'h0099; B = 16'h000; #100;
A = 16'h0099; B = 16'h001; #100;
A = 16'h0099; B = 16'h002; #100;
A = 16'h0099; B = 16'h003; #100;
A = 16'h0099; B = 16'h004; #100;
A = 16'h0099; B = 16'h005; #100;
A = 16'h0099; B = 16'h006; #100;
A = 16'h0099; B = 16'h007; #100;
A = 16'h0099; B = 16'h008; #100;
A = 16'h0099; B = 16'h009; #100;
A = 16'h0099; B = 16'h00A; #100;
A = 16'h0099; B = 16'h00B; #100;
A = 16'h0099; B = 16'h00C; #100;
A = 16'h0099; B = 16'h00D; #100;
A = 16'h0099; B = 16'h00E; #100;
A = 16'h0099; B = 16'h00F; #100;
A = 16'h0099; B = 16'h0010; #100;
A = 16'h0099; B = 16'h0011; #100;
A = 16'h0099; B = 16'h0012; #100;
A = 16'h0099; B = 16'h0013; #100;
A = 16'h0099; B = 16'h0014; #100;
A = 16'h0099; B = 16'h0015; #100;
A = 16'h0099; B = 16'h0016; #100;
A = 16'h0099; B = 16'h0017; #100;
A = 16'h0099; B = 16'h0018; #100;
A = 16'h0099; B = 16'h0019; #100;
A = 16'h0099; B = 16'h001A; #100;
A = 16'h0099; B = 16'h001B; #100;
A = 16'h0099; B = 16'h001C; #100;
A = 16'h0099; B = 16'h001D; #100;
A = 16'h0099; B = 16'h001E; #100;
A = 16'h0099; B = 16'h001F; #100;
A = 16'h0099; B = 16'h0020; #100;
A = 16'h0099; B = 16'h0021; #100;
A = 16'h0099; B = 16'h0022; #100;
A = 16'h0099; B = 16'h0023; #100;
A = 16'h0099; B = 16'h0024; #100;
A = 16'h0099; B = 16'h0025; #100;
A = 16'h0099; B = 16'h0026; #100;
A = 16'h0099; B = 16'h0027; #100;
A = 16'h0099; B = 16'h0028; #100;
A = 16'h0099; B = 16'h0029; #100;
A = 16'h0099; B = 16'h002A; #100;
A = 16'h0099; B = 16'h002B; #100;
A = 16'h0099; B = 16'h002C; #100;
A = 16'h0099; B = 16'h002D; #100;
A = 16'h0099; B = 16'h002E; #100;
A = 16'h0099; B = 16'h002F; #100;
A = 16'h0099; B = 16'h0030; #100;
A = 16'h0099; B = 16'h0031; #100;
A = 16'h0099; B = 16'h0032; #100;
A = 16'h0099; B = 16'h0033; #100;
A = 16'h0099; B = 16'h0034; #100;
A = 16'h0099; B = 16'h0035; #100;
A = 16'h0099; B = 16'h0036; #100;
A = 16'h0099; B = 16'h0037; #100;
A = 16'h0099; B = 16'h0038; #100;
A = 16'h0099; B = 16'h0039; #100;
A = 16'h0099; B = 16'h003A; #100;
A = 16'h0099; B = 16'h003B; #100;
A = 16'h0099; B = 16'h003C; #100;
A = 16'h0099; B = 16'h003D; #100;
A = 16'h0099; B = 16'h003E; #100;
A = 16'h0099; B = 16'h003F; #100;
A = 16'h0099; B = 16'h0040; #100;
A = 16'h0099; B = 16'h0041; #100;
A = 16'h0099; B = 16'h0042; #100;
A = 16'h0099; B = 16'h0043; #100;
A = 16'h0099; B = 16'h0044; #100;
A = 16'h0099; B = 16'h0045; #100;
A = 16'h0099; B = 16'h0046; #100;
A = 16'h0099; B = 16'h0047; #100;
A = 16'h0099; B = 16'h0048; #100;
A = 16'h0099; B = 16'h0049; #100;
A = 16'h0099; B = 16'h004A; #100;
A = 16'h0099; B = 16'h004B; #100;
A = 16'h0099; B = 16'h004C; #100;
A = 16'h0099; B = 16'h004D; #100;
A = 16'h0099; B = 16'h004E; #100;
A = 16'h0099; B = 16'h004F; #100;
A = 16'h0099; B = 16'h0050; #100;
A = 16'h0099; B = 16'h0051; #100;
A = 16'h0099; B = 16'h0052; #100;
A = 16'h0099; B = 16'h0053; #100;
A = 16'h0099; B = 16'h0054; #100;
A = 16'h0099; B = 16'h0055; #100;
A = 16'h0099; B = 16'h0056; #100;
A = 16'h0099; B = 16'h0057; #100;
A = 16'h0099; B = 16'h0058; #100;
A = 16'h0099; B = 16'h0059; #100;
A = 16'h0099; B = 16'h005A; #100;
A = 16'h0099; B = 16'h005B; #100;
A = 16'h0099; B = 16'h005C; #100;
A = 16'h0099; B = 16'h005D; #100;
A = 16'h0099; B = 16'h005E; #100;
A = 16'h0099; B = 16'h005F; #100;
A = 16'h0099; B = 16'h0060; #100;
A = 16'h0099; B = 16'h0061; #100;
A = 16'h0099; B = 16'h0062; #100;
A = 16'h0099; B = 16'h0063; #100;
A = 16'h0099; B = 16'h0064; #100;
A = 16'h0099; B = 16'h0065; #100;
A = 16'h0099; B = 16'h0066; #100;
A = 16'h0099; B = 16'h0067; #100;
A = 16'h0099; B = 16'h0068; #100;
A = 16'h0099; B = 16'h0069; #100;
A = 16'h0099; B = 16'h006A; #100;
A = 16'h0099; B = 16'h006B; #100;
A = 16'h0099; B = 16'h006C; #100;
A = 16'h0099; B = 16'h006D; #100;
A = 16'h0099; B = 16'h006E; #100;
A = 16'h0099; B = 16'h006F; #100;
A = 16'h0099; B = 16'h0070; #100;
A = 16'h0099; B = 16'h0071; #100;
A = 16'h0099; B = 16'h0072; #100;
A = 16'h0099; B = 16'h0073; #100;
A = 16'h0099; B = 16'h0074; #100;
A = 16'h0099; B = 16'h0075; #100;
A = 16'h0099; B = 16'h0076; #100;
A = 16'h0099; B = 16'h0077; #100;
A = 16'h0099; B = 16'h0078; #100;
A = 16'h0099; B = 16'h0079; #100;
A = 16'h0099; B = 16'h007A; #100;
A = 16'h0099; B = 16'h007B; #100;
A = 16'h0099; B = 16'h007C; #100;
A = 16'h0099; B = 16'h007D; #100;
A = 16'h0099; B = 16'h007E; #100;
A = 16'h0099; B = 16'h007F; #100;
A = 16'h0099; B = 16'h0080; #100;
A = 16'h0099; B = 16'h0081; #100;
A = 16'h0099; B = 16'h0082; #100;
A = 16'h0099; B = 16'h0083; #100;
A = 16'h0099; B = 16'h0084; #100;
A = 16'h0099; B = 16'h0085; #100;
A = 16'h0099; B = 16'h0086; #100;
A = 16'h0099; B = 16'h0087; #100;
A = 16'h0099; B = 16'h0088; #100;
A = 16'h0099; B = 16'h0089; #100;
A = 16'h0099; B = 16'h008A; #100;
A = 16'h0099; B = 16'h008B; #100;
A = 16'h0099; B = 16'h008C; #100;
A = 16'h0099; B = 16'h008D; #100;
A = 16'h0099; B = 16'h008E; #100;
A = 16'h0099; B = 16'h008F; #100;
A = 16'h0099; B = 16'h0090; #100;
A = 16'h0099; B = 16'h0091; #100;
A = 16'h0099; B = 16'h0092; #100;
A = 16'h0099; B = 16'h0093; #100;
A = 16'h0099; B = 16'h0094; #100;
A = 16'h0099; B = 16'h0095; #100;
A = 16'h0099; B = 16'h0096; #100;
A = 16'h0099; B = 16'h0097; #100;
A = 16'h0099; B = 16'h0098; #100;
A = 16'h0099; B = 16'h0099; #100;
A = 16'h0099; B = 16'h009A; #100;
A = 16'h0099; B = 16'h009B; #100;
A = 16'h0099; B = 16'h009C; #100;
A = 16'h0099; B = 16'h009D; #100;
A = 16'h0099; B = 16'h009E; #100;
A = 16'h0099; B = 16'h009F; #100;
A = 16'h0099; B = 16'h00A0; #100;
A = 16'h0099; B = 16'h00A1; #100;
A = 16'h0099; B = 16'h00A2; #100;
A = 16'h0099; B = 16'h00A3; #100;
A = 16'h0099; B = 16'h00A4; #100;
A = 16'h0099; B = 16'h00A5; #100;
A = 16'h0099; B = 16'h00A6; #100;
A = 16'h0099; B = 16'h00A7; #100;
A = 16'h0099; B = 16'h00A8; #100;
A = 16'h0099; B = 16'h00A9; #100;
A = 16'h0099; B = 16'h00AA; #100;
A = 16'h0099; B = 16'h00AB; #100;
A = 16'h0099; B = 16'h00AC; #100;
A = 16'h0099; B = 16'h00AD; #100;
A = 16'h0099; B = 16'h00AE; #100;
A = 16'h0099; B = 16'h00AF; #100;
A = 16'h0099; B = 16'h00B0; #100;
A = 16'h0099; B = 16'h00B1; #100;
A = 16'h0099; B = 16'h00B2; #100;
A = 16'h0099; B = 16'h00B3; #100;
A = 16'h0099; B = 16'h00B4; #100;
A = 16'h0099; B = 16'h00B5; #100;
A = 16'h0099; B = 16'h00B6; #100;
A = 16'h0099; B = 16'h00B7; #100;
A = 16'h0099; B = 16'h00B8; #100;
A = 16'h0099; B = 16'h00B9; #100;
A = 16'h0099; B = 16'h00BA; #100;
A = 16'h0099; B = 16'h00BB; #100;
A = 16'h0099; B = 16'h00BC; #100;
A = 16'h0099; B = 16'h00BD; #100;
A = 16'h0099; B = 16'h00BE; #100;
A = 16'h0099; B = 16'h00BF; #100;
A = 16'h0099; B = 16'h00C0; #100;
A = 16'h0099; B = 16'h00C1; #100;
A = 16'h0099; B = 16'h00C2; #100;
A = 16'h0099; B = 16'h00C3; #100;
A = 16'h0099; B = 16'h00C4; #100;
A = 16'h0099; B = 16'h00C5; #100;
A = 16'h0099; B = 16'h00C6; #100;
A = 16'h0099; B = 16'h00C7; #100;
A = 16'h0099; B = 16'h00C8; #100;
A = 16'h0099; B = 16'h00C9; #100;
A = 16'h0099; B = 16'h00CA; #100;
A = 16'h0099; B = 16'h00CB; #100;
A = 16'h0099; B = 16'h00CC; #100;
A = 16'h0099; B = 16'h00CD; #100;
A = 16'h0099; B = 16'h00CE; #100;
A = 16'h0099; B = 16'h00CF; #100;
A = 16'h0099; B = 16'h00D0; #100;
A = 16'h0099; B = 16'h00D1; #100;
A = 16'h0099; B = 16'h00D2; #100;
A = 16'h0099; B = 16'h00D3; #100;
A = 16'h0099; B = 16'h00D4; #100;
A = 16'h0099; B = 16'h00D5; #100;
A = 16'h0099; B = 16'h00D6; #100;
A = 16'h0099; B = 16'h00D7; #100;
A = 16'h0099; B = 16'h00D8; #100;
A = 16'h0099; B = 16'h00D9; #100;
A = 16'h0099; B = 16'h00DA; #100;
A = 16'h0099; B = 16'h00DB; #100;
A = 16'h0099; B = 16'h00DC; #100;
A = 16'h0099; B = 16'h00DD; #100;
A = 16'h0099; B = 16'h00DE; #100;
A = 16'h0099; B = 16'h00DF; #100;
A = 16'h0099; B = 16'h00E0; #100;
A = 16'h0099; B = 16'h00E1; #100;
A = 16'h0099; B = 16'h00E2; #100;
A = 16'h0099; B = 16'h00E3; #100;
A = 16'h0099; B = 16'h00E4; #100;
A = 16'h0099; B = 16'h00E5; #100;
A = 16'h0099; B = 16'h00E6; #100;
A = 16'h0099; B = 16'h00E7; #100;
A = 16'h0099; B = 16'h00E8; #100;
A = 16'h0099; B = 16'h00E9; #100;
A = 16'h0099; B = 16'h00EA; #100;
A = 16'h0099; B = 16'h00EB; #100;
A = 16'h0099; B = 16'h00EC; #100;
A = 16'h0099; B = 16'h00ED; #100;
A = 16'h0099; B = 16'h00EE; #100;
A = 16'h0099; B = 16'h00EF; #100;
A = 16'h0099; B = 16'h00F0; #100;
A = 16'h0099; B = 16'h00F1; #100;
A = 16'h0099; B = 16'h00F2; #100;
A = 16'h0099; B = 16'h00F3; #100;
A = 16'h0099; B = 16'h00F4; #100;
A = 16'h0099; B = 16'h00F5; #100;
A = 16'h0099; B = 16'h00F6; #100;
A = 16'h0099; B = 16'h00F7; #100;
A = 16'h0099; B = 16'h00F8; #100;
A = 16'h0099; B = 16'h00F9; #100;
A = 16'h0099; B = 16'h00FA; #100;
A = 16'h0099; B = 16'h00FB; #100;
A = 16'h0099; B = 16'h00FC; #100;
A = 16'h0099; B = 16'h00FD; #100;
A = 16'h0099; B = 16'h00FE; #100;
A = 16'h0099; B = 16'h00FF; #100;
A = 16'h009A; B = 16'h000; #100;
A = 16'h009A; B = 16'h001; #100;
A = 16'h009A; B = 16'h002; #100;
A = 16'h009A; B = 16'h003; #100;
A = 16'h009A; B = 16'h004; #100;
A = 16'h009A; B = 16'h005; #100;
A = 16'h009A; B = 16'h006; #100;
A = 16'h009A; B = 16'h007; #100;
A = 16'h009A; B = 16'h008; #100;
A = 16'h009A; B = 16'h009; #100;
A = 16'h009A; B = 16'h00A; #100;
A = 16'h009A; B = 16'h00B; #100;
A = 16'h009A; B = 16'h00C; #100;
A = 16'h009A; B = 16'h00D; #100;
A = 16'h009A; B = 16'h00E; #100;
A = 16'h009A; B = 16'h00F; #100;
A = 16'h009A; B = 16'h0010; #100;
A = 16'h009A; B = 16'h0011; #100;
A = 16'h009A; B = 16'h0012; #100;
A = 16'h009A; B = 16'h0013; #100;
A = 16'h009A; B = 16'h0014; #100;
A = 16'h009A; B = 16'h0015; #100;
A = 16'h009A; B = 16'h0016; #100;
A = 16'h009A; B = 16'h0017; #100;
A = 16'h009A; B = 16'h0018; #100;
A = 16'h009A; B = 16'h0019; #100;
A = 16'h009A; B = 16'h001A; #100;
A = 16'h009A; B = 16'h001B; #100;
A = 16'h009A; B = 16'h001C; #100;
A = 16'h009A; B = 16'h001D; #100;
A = 16'h009A; B = 16'h001E; #100;
A = 16'h009A; B = 16'h001F; #100;
A = 16'h009A; B = 16'h0020; #100;
A = 16'h009A; B = 16'h0021; #100;
A = 16'h009A; B = 16'h0022; #100;
A = 16'h009A; B = 16'h0023; #100;
A = 16'h009A; B = 16'h0024; #100;
A = 16'h009A; B = 16'h0025; #100;
A = 16'h009A; B = 16'h0026; #100;
A = 16'h009A; B = 16'h0027; #100;
A = 16'h009A; B = 16'h0028; #100;
A = 16'h009A; B = 16'h0029; #100;
A = 16'h009A; B = 16'h002A; #100;
A = 16'h009A; B = 16'h002B; #100;
A = 16'h009A; B = 16'h002C; #100;
A = 16'h009A; B = 16'h002D; #100;
A = 16'h009A; B = 16'h002E; #100;
A = 16'h009A; B = 16'h002F; #100;
A = 16'h009A; B = 16'h0030; #100;
A = 16'h009A; B = 16'h0031; #100;
A = 16'h009A; B = 16'h0032; #100;
A = 16'h009A; B = 16'h0033; #100;
A = 16'h009A; B = 16'h0034; #100;
A = 16'h009A; B = 16'h0035; #100;
A = 16'h009A; B = 16'h0036; #100;
A = 16'h009A; B = 16'h0037; #100;
A = 16'h009A; B = 16'h0038; #100;
A = 16'h009A; B = 16'h0039; #100;
A = 16'h009A; B = 16'h003A; #100;
A = 16'h009A; B = 16'h003B; #100;
A = 16'h009A; B = 16'h003C; #100;
A = 16'h009A; B = 16'h003D; #100;
A = 16'h009A; B = 16'h003E; #100;
A = 16'h009A; B = 16'h003F; #100;
A = 16'h009A; B = 16'h0040; #100;
A = 16'h009A; B = 16'h0041; #100;
A = 16'h009A; B = 16'h0042; #100;
A = 16'h009A; B = 16'h0043; #100;
A = 16'h009A; B = 16'h0044; #100;
A = 16'h009A; B = 16'h0045; #100;
A = 16'h009A; B = 16'h0046; #100;
A = 16'h009A; B = 16'h0047; #100;
A = 16'h009A; B = 16'h0048; #100;
A = 16'h009A; B = 16'h0049; #100;
A = 16'h009A; B = 16'h004A; #100;
A = 16'h009A; B = 16'h004B; #100;
A = 16'h009A; B = 16'h004C; #100;
A = 16'h009A; B = 16'h004D; #100;
A = 16'h009A; B = 16'h004E; #100;
A = 16'h009A; B = 16'h004F; #100;
A = 16'h009A; B = 16'h0050; #100;
A = 16'h009A; B = 16'h0051; #100;
A = 16'h009A; B = 16'h0052; #100;
A = 16'h009A; B = 16'h0053; #100;
A = 16'h009A; B = 16'h0054; #100;
A = 16'h009A; B = 16'h0055; #100;
A = 16'h009A; B = 16'h0056; #100;
A = 16'h009A; B = 16'h0057; #100;
A = 16'h009A; B = 16'h0058; #100;
A = 16'h009A; B = 16'h0059; #100;
A = 16'h009A; B = 16'h005A; #100;
A = 16'h009A; B = 16'h005B; #100;
A = 16'h009A; B = 16'h005C; #100;
A = 16'h009A; B = 16'h005D; #100;
A = 16'h009A; B = 16'h005E; #100;
A = 16'h009A; B = 16'h005F; #100;
A = 16'h009A; B = 16'h0060; #100;
A = 16'h009A; B = 16'h0061; #100;
A = 16'h009A; B = 16'h0062; #100;
A = 16'h009A; B = 16'h0063; #100;
A = 16'h009A; B = 16'h0064; #100;
A = 16'h009A; B = 16'h0065; #100;
A = 16'h009A; B = 16'h0066; #100;
A = 16'h009A; B = 16'h0067; #100;
A = 16'h009A; B = 16'h0068; #100;
A = 16'h009A; B = 16'h0069; #100;
A = 16'h009A; B = 16'h006A; #100;
A = 16'h009A; B = 16'h006B; #100;
A = 16'h009A; B = 16'h006C; #100;
A = 16'h009A; B = 16'h006D; #100;
A = 16'h009A; B = 16'h006E; #100;
A = 16'h009A; B = 16'h006F; #100;
A = 16'h009A; B = 16'h0070; #100;
A = 16'h009A; B = 16'h0071; #100;
A = 16'h009A; B = 16'h0072; #100;
A = 16'h009A; B = 16'h0073; #100;
A = 16'h009A; B = 16'h0074; #100;
A = 16'h009A; B = 16'h0075; #100;
A = 16'h009A; B = 16'h0076; #100;
A = 16'h009A; B = 16'h0077; #100;
A = 16'h009A; B = 16'h0078; #100;
A = 16'h009A; B = 16'h0079; #100;
A = 16'h009A; B = 16'h007A; #100;
A = 16'h009A; B = 16'h007B; #100;
A = 16'h009A; B = 16'h007C; #100;
A = 16'h009A; B = 16'h007D; #100;
A = 16'h009A; B = 16'h007E; #100;
A = 16'h009A; B = 16'h007F; #100;
A = 16'h009A; B = 16'h0080; #100;
A = 16'h009A; B = 16'h0081; #100;
A = 16'h009A; B = 16'h0082; #100;
A = 16'h009A; B = 16'h0083; #100;
A = 16'h009A; B = 16'h0084; #100;
A = 16'h009A; B = 16'h0085; #100;
A = 16'h009A; B = 16'h0086; #100;
A = 16'h009A; B = 16'h0087; #100;
A = 16'h009A; B = 16'h0088; #100;
A = 16'h009A; B = 16'h0089; #100;
A = 16'h009A; B = 16'h008A; #100;
A = 16'h009A; B = 16'h008B; #100;
A = 16'h009A; B = 16'h008C; #100;
A = 16'h009A; B = 16'h008D; #100;
A = 16'h009A; B = 16'h008E; #100;
A = 16'h009A; B = 16'h008F; #100;
A = 16'h009A; B = 16'h0090; #100;
A = 16'h009A; B = 16'h0091; #100;
A = 16'h009A; B = 16'h0092; #100;
A = 16'h009A; B = 16'h0093; #100;
A = 16'h009A; B = 16'h0094; #100;
A = 16'h009A; B = 16'h0095; #100;
A = 16'h009A; B = 16'h0096; #100;
A = 16'h009A; B = 16'h0097; #100;
A = 16'h009A; B = 16'h0098; #100;
A = 16'h009A; B = 16'h0099; #100;
A = 16'h009A; B = 16'h009A; #100;
A = 16'h009A; B = 16'h009B; #100;
A = 16'h009A; B = 16'h009C; #100;
A = 16'h009A; B = 16'h009D; #100;
A = 16'h009A; B = 16'h009E; #100;
A = 16'h009A; B = 16'h009F; #100;
A = 16'h009A; B = 16'h00A0; #100;
A = 16'h009A; B = 16'h00A1; #100;
A = 16'h009A; B = 16'h00A2; #100;
A = 16'h009A; B = 16'h00A3; #100;
A = 16'h009A; B = 16'h00A4; #100;
A = 16'h009A; B = 16'h00A5; #100;
A = 16'h009A; B = 16'h00A6; #100;
A = 16'h009A; B = 16'h00A7; #100;
A = 16'h009A; B = 16'h00A8; #100;
A = 16'h009A; B = 16'h00A9; #100;
A = 16'h009A; B = 16'h00AA; #100;
A = 16'h009A; B = 16'h00AB; #100;
A = 16'h009A; B = 16'h00AC; #100;
A = 16'h009A; B = 16'h00AD; #100;
A = 16'h009A; B = 16'h00AE; #100;
A = 16'h009A; B = 16'h00AF; #100;
A = 16'h009A; B = 16'h00B0; #100;
A = 16'h009A; B = 16'h00B1; #100;
A = 16'h009A; B = 16'h00B2; #100;
A = 16'h009A; B = 16'h00B3; #100;
A = 16'h009A; B = 16'h00B4; #100;
A = 16'h009A; B = 16'h00B5; #100;
A = 16'h009A; B = 16'h00B6; #100;
A = 16'h009A; B = 16'h00B7; #100;
A = 16'h009A; B = 16'h00B8; #100;
A = 16'h009A; B = 16'h00B9; #100;
A = 16'h009A; B = 16'h00BA; #100;
A = 16'h009A; B = 16'h00BB; #100;
A = 16'h009A; B = 16'h00BC; #100;
A = 16'h009A; B = 16'h00BD; #100;
A = 16'h009A; B = 16'h00BE; #100;
A = 16'h009A; B = 16'h00BF; #100;
A = 16'h009A; B = 16'h00C0; #100;
A = 16'h009A; B = 16'h00C1; #100;
A = 16'h009A; B = 16'h00C2; #100;
A = 16'h009A; B = 16'h00C3; #100;
A = 16'h009A; B = 16'h00C4; #100;
A = 16'h009A; B = 16'h00C5; #100;
A = 16'h009A; B = 16'h00C6; #100;
A = 16'h009A; B = 16'h00C7; #100;
A = 16'h009A; B = 16'h00C8; #100;
A = 16'h009A; B = 16'h00C9; #100;
A = 16'h009A; B = 16'h00CA; #100;
A = 16'h009A; B = 16'h00CB; #100;
A = 16'h009A; B = 16'h00CC; #100;
A = 16'h009A; B = 16'h00CD; #100;
A = 16'h009A; B = 16'h00CE; #100;
A = 16'h009A; B = 16'h00CF; #100;
A = 16'h009A; B = 16'h00D0; #100;
A = 16'h009A; B = 16'h00D1; #100;
A = 16'h009A; B = 16'h00D2; #100;
A = 16'h009A; B = 16'h00D3; #100;
A = 16'h009A; B = 16'h00D4; #100;
A = 16'h009A; B = 16'h00D5; #100;
A = 16'h009A; B = 16'h00D6; #100;
A = 16'h009A; B = 16'h00D7; #100;
A = 16'h009A; B = 16'h00D8; #100;
A = 16'h009A; B = 16'h00D9; #100;
A = 16'h009A; B = 16'h00DA; #100;
A = 16'h009A; B = 16'h00DB; #100;
A = 16'h009A; B = 16'h00DC; #100;
A = 16'h009A; B = 16'h00DD; #100;
A = 16'h009A; B = 16'h00DE; #100;
A = 16'h009A; B = 16'h00DF; #100;
A = 16'h009A; B = 16'h00E0; #100;
A = 16'h009A; B = 16'h00E1; #100;
A = 16'h009A; B = 16'h00E2; #100;
A = 16'h009A; B = 16'h00E3; #100;
A = 16'h009A; B = 16'h00E4; #100;
A = 16'h009A; B = 16'h00E5; #100;
A = 16'h009A; B = 16'h00E6; #100;
A = 16'h009A; B = 16'h00E7; #100;
A = 16'h009A; B = 16'h00E8; #100;
A = 16'h009A; B = 16'h00E9; #100;
A = 16'h009A; B = 16'h00EA; #100;
A = 16'h009A; B = 16'h00EB; #100;
A = 16'h009A; B = 16'h00EC; #100;
A = 16'h009A; B = 16'h00ED; #100;
A = 16'h009A; B = 16'h00EE; #100;
A = 16'h009A; B = 16'h00EF; #100;
A = 16'h009A; B = 16'h00F0; #100;
A = 16'h009A; B = 16'h00F1; #100;
A = 16'h009A; B = 16'h00F2; #100;
A = 16'h009A; B = 16'h00F3; #100;
A = 16'h009A; B = 16'h00F4; #100;
A = 16'h009A; B = 16'h00F5; #100;
A = 16'h009A; B = 16'h00F6; #100;
A = 16'h009A; B = 16'h00F7; #100;
A = 16'h009A; B = 16'h00F8; #100;
A = 16'h009A; B = 16'h00F9; #100;
A = 16'h009A; B = 16'h00FA; #100;
A = 16'h009A; B = 16'h00FB; #100;
A = 16'h009A; B = 16'h00FC; #100;
A = 16'h009A; B = 16'h00FD; #100;
A = 16'h009A; B = 16'h00FE; #100;
A = 16'h009A; B = 16'h00FF; #100;
A = 16'h009B; B = 16'h000; #100;
A = 16'h009B; B = 16'h001; #100;
A = 16'h009B; B = 16'h002; #100;
A = 16'h009B; B = 16'h003; #100;
A = 16'h009B; B = 16'h004; #100;
A = 16'h009B; B = 16'h005; #100;
A = 16'h009B; B = 16'h006; #100;
A = 16'h009B; B = 16'h007; #100;
A = 16'h009B; B = 16'h008; #100;
A = 16'h009B; B = 16'h009; #100;
A = 16'h009B; B = 16'h00A; #100;
A = 16'h009B; B = 16'h00B; #100;
A = 16'h009B; B = 16'h00C; #100;
A = 16'h009B; B = 16'h00D; #100;
A = 16'h009B; B = 16'h00E; #100;
A = 16'h009B; B = 16'h00F; #100;
A = 16'h009B; B = 16'h0010; #100;
A = 16'h009B; B = 16'h0011; #100;
A = 16'h009B; B = 16'h0012; #100;
A = 16'h009B; B = 16'h0013; #100;
A = 16'h009B; B = 16'h0014; #100;
A = 16'h009B; B = 16'h0015; #100;
A = 16'h009B; B = 16'h0016; #100;
A = 16'h009B; B = 16'h0017; #100;
A = 16'h009B; B = 16'h0018; #100;
A = 16'h009B; B = 16'h0019; #100;
A = 16'h009B; B = 16'h001A; #100;
A = 16'h009B; B = 16'h001B; #100;
A = 16'h009B; B = 16'h001C; #100;
A = 16'h009B; B = 16'h001D; #100;
A = 16'h009B; B = 16'h001E; #100;
A = 16'h009B; B = 16'h001F; #100;
A = 16'h009B; B = 16'h0020; #100;
A = 16'h009B; B = 16'h0021; #100;
A = 16'h009B; B = 16'h0022; #100;
A = 16'h009B; B = 16'h0023; #100;
A = 16'h009B; B = 16'h0024; #100;
A = 16'h009B; B = 16'h0025; #100;
A = 16'h009B; B = 16'h0026; #100;
A = 16'h009B; B = 16'h0027; #100;
A = 16'h009B; B = 16'h0028; #100;
A = 16'h009B; B = 16'h0029; #100;
A = 16'h009B; B = 16'h002A; #100;
A = 16'h009B; B = 16'h002B; #100;
A = 16'h009B; B = 16'h002C; #100;
A = 16'h009B; B = 16'h002D; #100;
A = 16'h009B; B = 16'h002E; #100;
A = 16'h009B; B = 16'h002F; #100;
A = 16'h009B; B = 16'h0030; #100;
A = 16'h009B; B = 16'h0031; #100;
A = 16'h009B; B = 16'h0032; #100;
A = 16'h009B; B = 16'h0033; #100;
A = 16'h009B; B = 16'h0034; #100;
A = 16'h009B; B = 16'h0035; #100;
A = 16'h009B; B = 16'h0036; #100;
A = 16'h009B; B = 16'h0037; #100;
A = 16'h009B; B = 16'h0038; #100;
A = 16'h009B; B = 16'h0039; #100;
A = 16'h009B; B = 16'h003A; #100;
A = 16'h009B; B = 16'h003B; #100;
A = 16'h009B; B = 16'h003C; #100;
A = 16'h009B; B = 16'h003D; #100;
A = 16'h009B; B = 16'h003E; #100;
A = 16'h009B; B = 16'h003F; #100;
A = 16'h009B; B = 16'h0040; #100;
A = 16'h009B; B = 16'h0041; #100;
A = 16'h009B; B = 16'h0042; #100;
A = 16'h009B; B = 16'h0043; #100;
A = 16'h009B; B = 16'h0044; #100;
A = 16'h009B; B = 16'h0045; #100;
A = 16'h009B; B = 16'h0046; #100;
A = 16'h009B; B = 16'h0047; #100;
A = 16'h009B; B = 16'h0048; #100;
A = 16'h009B; B = 16'h0049; #100;
A = 16'h009B; B = 16'h004A; #100;
A = 16'h009B; B = 16'h004B; #100;
A = 16'h009B; B = 16'h004C; #100;
A = 16'h009B; B = 16'h004D; #100;
A = 16'h009B; B = 16'h004E; #100;
A = 16'h009B; B = 16'h004F; #100;
A = 16'h009B; B = 16'h0050; #100;
A = 16'h009B; B = 16'h0051; #100;
A = 16'h009B; B = 16'h0052; #100;
A = 16'h009B; B = 16'h0053; #100;
A = 16'h009B; B = 16'h0054; #100;
A = 16'h009B; B = 16'h0055; #100;
A = 16'h009B; B = 16'h0056; #100;
A = 16'h009B; B = 16'h0057; #100;
A = 16'h009B; B = 16'h0058; #100;
A = 16'h009B; B = 16'h0059; #100;
A = 16'h009B; B = 16'h005A; #100;
A = 16'h009B; B = 16'h005B; #100;
A = 16'h009B; B = 16'h005C; #100;
A = 16'h009B; B = 16'h005D; #100;
A = 16'h009B; B = 16'h005E; #100;
A = 16'h009B; B = 16'h005F; #100;
A = 16'h009B; B = 16'h0060; #100;
A = 16'h009B; B = 16'h0061; #100;
A = 16'h009B; B = 16'h0062; #100;
A = 16'h009B; B = 16'h0063; #100;
A = 16'h009B; B = 16'h0064; #100;
A = 16'h009B; B = 16'h0065; #100;
A = 16'h009B; B = 16'h0066; #100;
A = 16'h009B; B = 16'h0067; #100;
A = 16'h009B; B = 16'h0068; #100;
A = 16'h009B; B = 16'h0069; #100;
A = 16'h009B; B = 16'h006A; #100;
A = 16'h009B; B = 16'h006B; #100;
A = 16'h009B; B = 16'h006C; #100;
A = 16'h009B; B = 16'h006D; #100;
A = 16'h009B; B = 16'h006E; #100;
A = 16'h009B; B = 16'h006F; #100;
A = 16'h009B; B = 16'h0070; #100;
A = 16'h009B; B = 16'h0071; #100;
A = 16'h009B; B = 16'h0072; #100;
A = 16'h009B; B = 16'h0073; #100;
A = 16'h009B; B = 16'h0074; #100;
A = 16'h009B; B = 16'h0075; #100;
A = 16'h009B; B = 16'h0076; #100;
A = 16'h009B; B = 16'h0077; #100;
A = 16'h009B; B = 16'h0078; #100;
A = 16'h009B; B = 16'h0079; #100;
A = 16'h009B; B = 16'h007A; #100;
A = 16'h009B; B = 16'h007B; #100;
A = 16'h009B; B = 16'h007C; #100;
A = 16'h009B; B = 16'h007D; #100;
A = 16'h009B; B = 16'h007E; #100;
A = 16'h009B; B = 16'h007F; #100;
A = 16'h009B; B = 16'h0080; #100;
A = 16'h009B; B = 16'h0081; #100;
A = 16'h009B; B = 16'h0082; #100;
A = 16'h009B; B = 16'h0083; #100;
A = 16'h009B; B = 16'h0084; #100;
A = 16'h009B; B = 16'h0085; #100;
A = 16'h009B; B = 16'h0086; #100;
A = 16'h009B; B = 16'h0087; #100;
A = 16'h009B; B = 16'h0088; #100;
A = 16'h009B; B = 16'h0089; #100;
A = 16'h009B; B = 16'h008A; #100;
A = 16'h009B; B = 16'h008B; #100;
A = 16'h009B; B = 16'h008C; #100;
A = 16'h009B; B = 16'h008D; #100;
A = 16'h009B; B = 16'h008E; #100;
A = 16'h009B; B = 16'h008F; #100;
A = 16'h009B; B = 16'h0090; #100;
A = 16'h009B; B = 16'h0091; #100;
A = 16'h009B; B = 16'h0092; #100;
A = 16'h009B; B = 16'h0093; #100;
A = 16'h009B; B = 16'h0094; #100;
A = 16'h009B; B = 16'h0095; #100;
A = 16'h009B; B = 16'h0096; #100;
A = 16'h009B; B = 16'h0097; #100;
A = 16'h009B; B = 16'h0098; #100;
A = 16'h009B; B = 16'h0099; #100;
A = 16'h009B; B = 16'h009A; #100;
A = 16'h009B; B = 16'h009B; #100;
A = 16'h009B; B = 16'h009C; #100;
A = 16'h009B; B = 16'h009D; #100;
A = 16'h009B; B = 16'h009E; #100;
A = 16'h009B; B = 16'h009F; #100;
A = 16'h009B; B = 16'h00A0; #100;
A = 16'h009B; B = 16'h00A1; #100;
A = 16'h009B; B = 16'h00A2; #100;
A = 16'h009B; B = 16'h00A3; #100;
A = 16'h009B; B = 16'h00A4; #100;
A = 16'h009B; B = 16'h00A5; #100;
A = 16'h009B; B = 16'h00A6; #100;
A = 16'h009B; B = 16'h00A7; #100;
A = 16'h009B; B = 16'h00A8; #100;
A = 16'h009B; B = 16'h00A9; #100;
A = 16'h009B; B = 16'h00AA; #100;
A = 16'h009B; B = 16'h00AB; #100;
A = 16'h009B; B = 16'h00AC; #100;
A = 16'h009B; B = 16'h00AD; #100;
A = 16'h009B; B = 16'h00AE; #100;
A = 16'h009B; B = 16'h00AF; #100;
A = 16'h009B; B = 16'h00B0; #100;
A = 16'h009B; B = 16'h00B1; #100;
A = 16'h009B; B = 16'h00B2; #100;
A = 16'h009B; B = 16'h00B3; #100;
A = 16'h009B; B = 16'h00B4; #100;
A = 16'h009B; B = 16'h00B5; #100;
A = 16'h009B; B = 16'h00B6; #100;
A = 16'h009B; B = 16'h00B7; #100;
A = 16'h009B; B = 16'h00B8; #100;
A = 16'h009B; B = 16'h00B9; #100;
A = 16'h009B; B = 16'h00BA; #100;
A = 16'h009B; B = 16'h00BB; #100;
A = 16'h009B; B = 16'h00BC; #100;
A = 16'h009B; B = 16'h00BD; #100;
A = 16'h009B; B = 16'h00BE; #100;
A = 16'h009B; B = 16'h00BF; #100;
A = 16'h009B; B = 16'h00C0; #100;
A = 16'h009B; B = 16'h00C1; #100;
A = 16'h009B; B = 16'h00C2; #100;
A = 16'h009B; B = 16'h00C3; #100;
A = 16'h009B; B = 16'h00C4; #100;
A = 16'h009B; B = 16'h00C5; #100;
A = 16'h009B; B = 16'h00C6; #100;
A = 16'h009B; B = 16'h00C7; #100;
A = 16'h009B; B = 16'h00C8; #100;
A = 16'h009B; B = 16'h00C9; #100;
A = 16'h009B; B = 16'h00CA; #100;
A = 16'h009B; B = 16'h00CB; #100;
A = 16'h009B; B = 16'h00CC; #100;
A = 16'h009B; B = 16'h00CD; #100;
A = 16'h009B; B = 16'h00CE; #100;
A = 16'h009B; B = 16'h00CF; #100;
A = 16'h009B; B = 16'h00D0; #100;
A = 16'h009B; B = 16'h00D1; #100;
A = 16'h009B; B = 16'h00D2; #100;
A = 16'h009B; B = 16'h00D3; #100;
A = 16'h009B; B = 16'h00D4; #100;
A = 16'h009B; B = 16'h00D5; #100;
A = 16'h009B; B = 16'h00D6; #100;
A = 16'h009B; B = 16'h00D7; #100;
A = 16'h009B; B = 16'h00D8; #100;
A = 16'h009B; B = 16'h00D9; #100;
A = 16'h009B; B = 16'h00DA; #100;
A = 16'h009B; B = 16'h00DB; #100;
A = 16'h009B; B = 16'h00DC; #100;
A = 16'h009B; B = 16'h00DD; #100;
A = 16'h009B; B = 16'h00DE; #100;
A = 16'h009B; B = 16'h00DF; #100;
A = 16'h009B; B = 16'h00E0; #100;
A = 16'h009B; B = 16'h00E1; #100;
A = 16'h009B; B = 16'h00E2; #100;
A = 16'h009B; B = 16'h00E3; #100;
A = 16'h009B; B = 16'h00E4; #100;
A = 16'h009B; B = 16'h00E5; #100;
A = 16'h009B; B = 16'h00E6; #100;
A = 16'h009B; B = 16'h00E7; #100;
A = 16'h009B; B = 16'h00E8; #100;
A = 16'h009B; B = 16'h00E9; #100;
A = 16'h009B; B = 16'h00EA; #100;
A = 16'h009B; B = 16'h00EB; #100;
A = 16'h009B; B = 16'h00EC; #100;
A = 16'h009B; B = 16'h00ED; #100;
A = 16'h009B; B = 16'h00EE; #100;
A = 16'h009B; B = 16'h00EF; #100;
A = 16'h009B; B = 16'h00F0; #100;
A = 16'h009B; B = 16'h00F1; #100;
A = 16'h009B; B = 16'h00F2; #100;
A = 16'h009B; B = 16'h00F3; #100;
A = 16'h009B; B = 16'h00F4; #100;
A = 16'h009B; B = 16'h00F5; #100;
A = 16'h009B; B = 16'h00F6; #100;
A = 16'h009B; B = 16'h00F7; #100;
A = 16'h009B; B = 16'h00F8; #100;
A = 16'h009B; B = 16'h00F9; #100;
A = 16'h009B; B = 16'h00FA; #100;
A = 16'h009B; B = 16'h00FB; #100;
A = 16'h009B; B = 16'h00FC; #100;
A = 16'h009B; B = 16'h00FD; #100;
A = 16'h009B; B = 16'h00FE; #100;
A = 16'h009B; B = 16'h00FF; #100;
A = 16'h009C; B = 16'h000; #100;
A = 16'h009C; B = 16'h001; #100;
A = 16'h009C; B = 16'h002; #100;
A = 16'h009C; B = 16'h003; #100;
A = 16'h009C; B = 16'h004; #100;
A = 16'h009C; B = 16'h005; #100;
A = 16'h009C; B = 16'h006; #100;
A = 16'h009C; B = 16'h007; #100;
A = 16'h009C; B = 16'h008; #100;
A = 16'h009C; B = 16'h009; #100;
A = 16'h009C; B = 16'h00A; #100;
A = 16'h009C; B = 16'h00B; #100;
A = 16'h009C; B = 16'h00C; #100;
A = 16'h009C; B = 16'h00D; #100;
A = 16'h009C; B = 16'h00E; #100;
A = 16'h009C; B = 16'h00F; #100;
A = 16'h009C; B = 16'h0010; #100;
A = 16'h009C; B = 16'h0011; #100;
A = 16'h009C; B = 16'h0012; #100;
A = 16'h009C; B = 16'h0013; #100;
A = 16'h009C; B = 16'h0014; #100;
A = 16'h009C; B = 16'h0015; #100;
A = 16'h009C; B = 16'h0016; #100;
A = 16'h009C; B = 16'h0017; #100;
A = 16'h009C; B = 16'h0018; #100;
A = 16'h009C; B = 16'h0019; #100;
A = 16'h009C; B = 16'h001A; #100;
A = 16'h009C; B = 16'h001B; #100;
A = 16'h009C; B = 16'h001C; #100;
A = 16'h009C; B = 16'h001D; #100;
A = 16'h009C; B = 16'h001E; #100;
A = 16'h009C; B = 16'h001F; #100;
A = 16'h009C; B = 16'h0020; #100;
A = 16'h009C; B = 16'h0021; #100;
A = 16'h009C; B = 16'h0022; #100;
A = 16'h009C; B = 16'h0023; #100;
A = 16'h009C; B = 16'h0024; #100;
A = 16'h009C; B = 16'h0025; #100;
A = 16'h009C; B = 16'h0026; #100;
A = 16'h009C; B = 16'h0027; #100;
A = 16'h009C; B = 16'h0028; #100;
A = 16'h009C; B = 16'h0029; #100;
A = 16'h009C; B = 16'h002A; #100;
A = 16'h009C; B = 16'h002B; #100;
A = 16'h009C; B = 16'h002C; #100;
A = 16'h009C; B = 16'h002D; #100;
A = 16'h009C; B = 16'h002E; #100;
A = 16'h009C; B = 16'h002F; #100;
A = 16'h009C; B = 16'h0030; #100;
A = 16'h009C; B = 16'h0031; #100;
A = 16'h009C; B = 16'h0032; #100;
A = 16'h009C; B = 16'h0033; #100;
A = 16'h009C; B = 16'h0034; #100;
A = 16'h009C; B = 16'h0035; #100;
A = 16'h009C; B = 16'h0036; #100;
A = 16'h009C; B = 16'h0037; #100;
A = 16'h009C; B = 16'h0038; #100;
A = 16'h009C; B = 16'h0039; #100;
A = 16'h009C; B = 16'h003A; #100;
A = 16'h009C; B = 16'h003B; #100;
A = 16'h009C; B = 16'h003C; #100;
A = 16'h009C; B = 16'h003D; #100;
A = 16'h009C; B = 16'h003E; #100;
A = 16'h009C; B = 16'h003F; #100;
A = 16'h009C; B = 16'h0040; #100;
A = 16'h009C; B = 16'h0041; #100;
A = 16'h009C; B = 16'h0042; #100;
A = 16'h009C; B = 16'h0043; #100;
A = 16'h009C; B = 16'h0044; #100;
A = 16'h009C; B = 16'h0045; #100;
A = 16'h009C; B = 16'h0046; #100;
A = 16'h009C; B = 16'h0047; #100;
A = 16'h009C; B = 16'h0048; #100;
A = 16'h009C; B = 16'h0049; #100;
A = 16'h009C; B = 16'h004A; #100;
A = 16'h009C; B = 16'h004B; #100;
A = 16'h009C; B = 16'h004C; #100;
A = 16'h009C; B = 16'h004D; #100;
A = 16'h009C; B = 16'h004E; #100;
A = 16'h009C; B = 16'h004F; #100;
A = 16'h009C; B = 16'h0050; #100;
A = 16'h009C; B = 16'h0051; #100;
A = 16'h009C; B = 16'h0052; #100;
A = 16'h009C; B = 16'h0053; #100;
A = 16'h009C; B = 16'h0054; #100;
A = 16'h009C; B = 16'h0055; #100;
A = 16'h009C; B = 16'h0056; #100;
A = 16'h009C; B = 16'h0057; #100;
A = 16'h009C; B = 16'h0058; #100;
A = 16'h009C; B = 16'h0059; #100;
A = 16'h009C; B = 16'h005A; #100;
A = 16'h009C; B = 16'h005B; #100;
A = 16'h009C; B = 16'h005C; #100;
A = 16'h009C; B = 16'h005D; #100;
A = 16'h009C; B = 16'h005E; #100;
A = 16'h009C; B = 16'h005F; #100;
A = 16'h009C; B = 16'h0060; #100;
A = 16'h009C; B = 16'h0061; #100;
A = 16'h009C; B = 16'h0062; #100;
A = 16'h009C; B = 16'h0063; #100;
A = 16'h009C; B = 16'h0064; #100;
A = 16'h009C; B = 16'h0065; #100;
A = 16'h009C; B = 16'h0066; #100;
A = 16'h009C; B = 16'h0067; #100;
A = 16'h009C; B = 16'h0068; #100;
A = 16'h009C; B = 16'h0069; #100;
A = 16'h009C; B = 16'h006A; #100;
A = 16'h009C; B = 16'h006B; #100;
A = 16'h009C; B = 16'h006C; #100;
A = 16'h009C; B = 16'h006D; #100;
A = 16'h009C; B = 16'h006E; #100;
A = 16'h009C; B = 16'h006F; #100;
A = 16'h009C; B = 16'h0070; #100;
A = 16'h009C; B = 16'h0071; #100;
A = 16'h009C; B = 16'h0072; #100;
A = 16'h009C; B = 16'h0073; #100;
A = 16'h009C; B = 16'h0074; #100;
A = 16'h009C; B = 16'h0075; #100;
A = 16'h009C; B = 16'h0076; #100;
A = 16'h009C; B = 16'h0077; #100;
A = 16'h009C; B = 16'h0078; #100;
A = 16'h009C; B = 16'h0079; #100;
A = 16'h009C; B = 16'h007A; #100;
A = 16'h009C; B = 16'h007B; #100;
A = 16'h009C; B = 16'h007C; #100;
A = 16'h009C; B = 16'h007D; #100;
A = 16'h009C; B = 16'h007E; #100;
A = 16'h009C; B = 16'h007F; #100;
A = 16'h009C; B = 16'h0080; #100;
A = 16'h009C; B = 16'h0081; #100;
A = 16'h009C; B = 16'h0082; #100;
A = 16'h009C; B = 16'h0083; #100;
A = 16'h009C; B = 16'h0084; #100;
A = 16'h009C; B = 16'h0085; #100;
A = 16'h009C; B = 16'h0086; #100;
A = 16'h009C; B = 16'h0087; #100;
A = 16'h009C; B = 16'h0088; #100;
A = 16'h009C; B = 16'h0089; #100;
A = 16'h009C; B = 16'h008A; #100;
A = 16'h009C; B = 16'h008B; #100;
A = 16'h009C; B = 16'h008C; #100;
A = 16'h009C; B = 16'h008D; #100;
A = 16'h009C; B = 16'h008E; #100;
A = 16'h009C; B = 16'h008F; #100;
A = 16'h009C; B = 16'h0090; #100;
A = 16'h009C; B = 16'h0091; #100;
A = 16'h009C; B = 16'h0092; #100;
A = 16'h009C; B = 16'h0093; #100;
A = 16'h009C; B = 16'h0094; #100;
A = 16'h009C; B = 16'h0095; #100;
A = 16'h009C; B = 16'h0096; #100;
A = 16'h009C; B = 16'h0097; #100;
A = 16'h009C; B = 16'h0098; #100;
A = 16'h009C; B = 16'h0099; #100;
A = 16'h009C; B = 16'h009A; #100;
A = 16'h009C; B = 16'h009B; #100;
A = 16'h009C; B = 16'h009C; #100;
A = 16'h009C; B = 16'h009D; #100;
A = 16'h009C; B = 16'h009E; #100;
A = 16'h009C; B = 16'h009F; #100;
A = 16'h009C; B = 16'h00A0; #100;
A = 16'h009C; B = 16'h00A1; #100;
A = 16'h009C; B = 16'h00A2; #100;
A = 16'h009C; B = 16'h00A3; #100;
A = 16'h009C; B = 16'h00A4; #100;
A = 16'h009C; B = 16'h00A5; #100;
A = 16'h009C; B = 16'h00A6; #100;
A = 16'h009C; B = 16'h00A7; #100;
A = 16'h009C; B = 16'h00A8; #100;
A = 16'h009C; B = 16'h00A9; #100;
A = 16'h009C; B = 16'h00AA; #100;
A = 16'h009C; B = 16'h00AB; #100;
A = 16'h009C; B = 16'h00AC; #100;
A = 16'h009C; B = 16'h00AD; #100;
A = 16'h009C; B = 16'h00AE; #100;
A = 16'h009C; B = 16'h00AF; #100;
A = 16'h009C; B = 16'h00B0; #100;
A = 16'h009C; B = 16'h00B1; #100;
A = 16'h009C; B = 16'h00B2; #100;
A = 16'h009C; B = 16'h00B3; #100;
A = 16'h009C; B = 16'h00B4; #100;
A = 16'h009C; B = 16'h00B5; #100;
A = 16'h009C; B = 16'h00B6; #100;
A = 16'h009C; B = 16'h00B7; #100;
A = 16'h009C; B = 16'h00B8; #100;
A = 16'h009C; B = 16'h00B9; #100;
A = 16'h009C; B = 16'h00BA; #100;
A = 16'h009C; B = 16'h00BB; #100;
A = 16'h009C; B = 16'h00BC; #100;
A = 16'h009C; B = 16'h00BD; #100;
A = 16'h009C; B = 16'h00BE; #100;
A = 16'h009C; B = 16'h00BF; #100;
A = 16'h009C; B = 16'h00C0; #100;
A = 16'h009C; B = 16'h00C1; #100;
A = 16'h009C; B = 16'h00C2; #100;
A = 16'h009C; B = 16'h00C3; #100;
A = 16'h009C; B = 16'h00C4; #100;
A = 16'h009C; B = 16'h00C5; #100;
A = 16'h009C; B = 16'h00C6; #100;
A = 16'h009C; B = 16'h00C7; #100;
A = 16'h009C; B = 16'h00C8; #100;
A = 16'h009C; B = 16'h00C9; #100;
A = 16'h009C; B = 16'h00CA; #100;
A = 16'h009C; B = 16'h00CB; #100;
A = 16'h009C; B = 16'h00CC; #100;
A = 16'h009C; B = 16'h00CD; #100;
A = 16'h009C; B = 16'h00CE; #100;
A = 16'h009C; B = 16'h00CF; #100;
A = 16'h009C; B = 16'h00D0; #100;
A = 16'h009C; B = 16'h00D1; #100;
A = 16'h009C; B = 16'h00D2; #100;
A = 16'h009C; B = 16'h00D3; #100;
A = 16'h009C; B = 16'h00D4; #100;
A = 16'h009C; B = 16'h00D5; #100;
A = 16'h009C; B = 16'h00D6; #100;
A = 16'h009C; B = 16'h00D7; #100;
A = 16'h009C; B = 16'h00D8; #100;
A = 16'h009C; B = 16'h00D9; #100;
A = 16'h009C; B = 16'h00DA; #100;
A = 16'h009C; B = 16'h00DB; #100;
A = 16'h009C; B = 16'h00DC; #100;
A = 16'h009C; B = 16'h00DD; #100;
A = 16'h009C; B = 16'h00DE; #100;
A = 16'h009C; B = 16'h00DF; #100;
A = 16'h009C; B = 16'h00E0; #100;
A = 16'h009C; B = 16'h00E1; #100;
A = 16'h009C; B = 16'h00E2; #100;
A = 16'h009C; B = 16'h00E3; #100;
A = 16'h009C; B = 16'h00E4; #100;
A = 16'h009C; B = 16'h00E5; #100;
A = 16'h009C; B = 16'h00E6; #100;
A = 16'h009C; B = 16'h00E7; #100;
A = 16'h009C; B = 16'h00E8; #100;
A = 16'h009C; B = 16'h00E9; #100;
A = 16'h009C; B = 16'h00EA; #100;
A = 16'h009C; B = 16'h00EB; #100;
A = 16'h009C; B = 16'h00EC; #100;
A = 16'h009C; B = 16'h00ED; #100;
A = 16'h009C; B = 16'h00EE; #100;
A = 16'h009C; B = 16'h00EF; #100;
A = 16'h009C; B = 16'h00F0; #100;
A = 16'h009C; B = 16'h00F1; #100;
A = 16'h009C; B = 16'h00F2; #100;
A = 16'h009C; B = 16'h00F3; #100;
A = 16'h009C; B = 16'h00F4; #100;
A = 16'h009C; B = 16'h00F5; #100;
A = 16'h009C; B = 16'h00F6; #100;
A = 16'h009C; B = 16'h00F7; #100;
A = 16'h009C; B = 16'h00F8; #100;
A = 16'h009C; B = 16'h00F9; #100;
A = 16'h009C; B = 16'h00FA; #100;
A = 16'h009C; B = 16'h00FB; #100;
A = 16'h009C; B = 16'h00FC; #100;
A = 16'h009C; B = 16'h00FD; #100;
A = 16'h009C; B = 16'h00FE; #100;
A = 16'h009C; B = 16'h00FF; #100;
A = 16'h009D; B = 16'h000; #100;
A = 16'h009D; B = 16'h001; #100;
A = 16'h009D; B = 16'h002; #100;
A = 16'h009D; B = 16'h003; #100;
A = 16'h009D; B = 16'h004; #100;
A = 16'h009D; B = 16'h005; #100;
A = 16'h009D; B = 16'h006; #100;
A = 16'h009D; B = 16'h007; #100;
A = 16'h009D; B = 16'h008; #100;
A = 16'h009D; B = 16'h009; #100;
A = 16'h009D; B = 16'h00A; #100;
A = 16'h009D; B = 16'h00B; #100;
A = 16'h009D; B = 16'h00C; #100;
A = 16'h009D; B = 16'h00D; #100;
A = 16'h009D; B = 16'h00E; #100;
A = 16'h009D; B = 16'h00F; #100;
A = 16'h009D; B = 16'h0010; #100;
A = 16'h009D; B = 16'h0011; #100;
A = 16'h009D; B = 16'h0012; #100;
A = 16'h009D; B = 16'h0013; #100;
A = 16'h009D; B = 16'h0014; #100;
A = 16'h009D; B = 16'h0015; #100;
A = 16'h009D; B = 16'h0016; #100;
A = 16'h009D; B = 16'h0017; #100;
A = 16'h009D; B = 16'h0018; #100;
A = 16'h009D; B = 16'h0019; #100;
A = 16'h009D; B = 16'h001A; #100;
A = 16'h009D; B = 16'h001B; #100;
A = 16'h009D; B = 16'h001C; #100;
A = 16'h009D; B = 16'h001D; #100;
A = 16'h009D; B = 16'h001E; #100;
A = 16'h009D; B = 16'h001F; #100;
A = 16'h009D; B = 16'h0020; #100;
A = 16'h009D; B = 16'h0021; #100;
A = 16'h009D; B = 16'h0022; #100;
A = 16'h009D; B = 16'h0023; #100;
A = 16'h009D; B = 16'h0024; #100;
A = 16'h009D; B = 16'h0025; #100;
A = 16'h009D; B = 16'h0026; #100;
A = 16'h009D; B = 16'h0027; #100;
A = 16'h009D; B = 16'h0028; #100;
A = 16'h009D; B = 16'h0029; #100;
A = 16'h009D; B = 16'h002A; #100;
A = 16'h009D; B = 16'h002B; #100;
A = 16'h009D; B = 16'h002C; #100;
A = 16'h009D; B = 16'h002D; #100;
A = 16'h009D; B = 16'h002E; #100;
A = 16'h009D; B = 16'h002F; #100;
A = 16'h009D; B = 16'h0030; #100;
A = 16'h009D; B = 16'h0031; #100;
A = 16'h009D; B = 16'h0032; #100;
A = 16'h009D; B = 16'h0033; #100;
A = 16'h009D; B = 16'h0034; #100;
A = 16'h009D; B = 16'h0035; #100;
A = 16'h009D; B = 16'h0036; #100;
A = 16'h009D; B = 16'h0037; #100;
A = 16'h009D; B = 16'h0038; #100;
A = 16'h009D; B = 16'h0039; #100;
A = 16'h009D; B = 16'h003A; #100;
A = 16'h009D; B = 16'h003B; #100;
A = 16'h009D; B = 16'h003C; #100;
A = 16'h009D; B = 16'h003D; #100;
A = 16'h009D; B = 16'h003E; #100;
A = 16'h009D; B = 16'h003F; #100;
A = 16'h009D; B = 16'h0040; #100;
A = 16'h009D; B = 16'h0041; #100;
A = 16'h009D; B = 16'h0042; #100;
A = 16'h009D; B = 16'h0043; #100;
A = 16'h009D; B = 16'h0044; #100;
A = 16'h009D; B = 16'h0045; #100;
A = 16'h009D; B = 16'h0046; #100;
A = 16'h009D; B = 16'h0047; #100;
A = 16'h009D; B = 16'h0048; #100;
A = 16'h009D; B = 16'h0049; #100;
A = 16'h009D; B = 16'h004A; #100;
A = 16'h009D; B = 16'h004B; #100;
A = 16'h009D; B = 16'h004C; #100;
A = 16'h009D; B = 16'h004D; #100;
A = 16'h009D; B = 16'h004E; #100;
A = 16'h009D; B = 16'h004F; #100;
A = 16'h009D; B = 16'h0050; #100;
A = 16'h009D; B = 16'h0051; #100;
A = 16'h009D; B = 16'h0052; #100;
A = 16'h009D; B = 16'h0053; #100;
A = 16'h009D; B = 16'h0054; #100;
A = 16'h009D; B = 16'h0055; #100;
A = 16'h009D; B = 16'h0056; #100;
A = 16'h009D; B = 16'h0057; #100;
A = 16'h009D; B = 16'h0058; #100;
A = 16'h009D; B = 16'h0059; #100;
A = 16'h009D; B = 16'h005A; #100;
A = 16'h009D; B = 16'h005B; #100;
A = 16'h009D; B = 16'h005C; #100;
A = 16'h009D; B = 16'h005D; #100;
A = 16'h009D; B = 16'h005E; #100;
A = 16'h009D; B = 16'h005F; #100;
A = 16'h009D; B = 16'h0060; #100;
A = 16'h009D; B = 16'h0061; #100;
A = 16'h009D; B = 16'h0062; #100;
A = 16'h009D; B = 16'h0063; #100;
A = 16'h009D; B = 16'h0064; #100;
A = 16'h009D; B = 16'h0065; #100;
A = 16'h009D; B = 16'h0066; #100;
A = 16'h009D; B = 16'h0067; #100;
A = 16'h009D; B = 16'h0068; #100;
A = 16'h009D; B = 16'h0069; #100;
A = 16'h009D; B = 16'h006A; #100;
A = 16'h009D; B = 16'h006B; #100;
A = 16'h009D; B = 16'h006C; #100;
A = 16'h009D; B = 16'h006D; #100;
A = 16'h009D; B = 16'h006E; #100;
A = 16'h009D; B = 16'h006F; #100;
A = 16'h009D; B = 16'h0070; #100;
A = 16'h009D; B = 16'h0071; #100;
A = 16'h009D; B = 16'h0072; #100;
A = 16'h009D; B = 16'h0073; #100;
A = 16'h009D; B = 16'h0074; #100;
A = 16'h009D; B = 16'h0075; #100;
A = 16'h009D; B = 16'h0076; #100;
A = 16'h009D; B = 16'h0077; #100;
A = 16'h009D; B = 16'h0078; #100;
A = 16'h009D; B = 16'h0079; #100;
A = 16'h009D; B = 16'h007A; #100;
A = 16'h009D; B = 16'h007B; #100;
A = 16'h009D; B = 16'h007C; #100;
A = 16'h009D; B = 16'h007D; #100;
A = 16'h009D; B = 16'h007E; #100;
A = 16'h009D; B = 16'h007F; #100;
A = 16'h009D; B = 16'h0080; #100;
A = 16'h009D; B = 16'h0081; #100;
A = 16'h009D; B = 16'h0082; #100;
A = 16'h009D; B = 16'h0083; #100;
A = 16'h009D; B = 16'h0084; #100;
A = 16'h009D; B = 16'h0085; #100;
A = 16'h009D; B = 16'h0086; #100;
A = 16'h009D; B = 16'h0087; #100;
A = 16'h009D; B = 16'h0088; #100;
A = 16'h009D; B = 16'h0089; #100;
A = 16'h009D; B = 16'h008A; #100;
A = 16'h009D; B = 16'h008B; #100;
A = 16'h009D; B = 16'h008C; #100;
A = 16'h009D; B = 16'h008D; #100;
A = 16'h009D; B = 16'h008E; #100;
A = 16'h009D; B = 16'h008F; #100;
A = 16'h009D; B = 16'h0090; #100;
A = 16'h009D; B = 16'h0091; #100;
A = 16'h009D; B = 16'h0092; #100;
A = 16'h009D; B = 16'h0093; #100;
A = 16'h009D; B = 16'h0094; #100;
A = 16'h009D; B = 16'h0095; #100;
A = 16'h009D; B = 16'h0096; #100;
A = 16'h009D; B = 16'h0097; #100;
A = 16'h009D; B = 16'h0098; #100;
A = 16'h009D; B = 16'h0099; #100;
A = 16'h009D; B = 16'h009A; #100;
A = 16'h009D; B = 16'h009B; #100;
A = 16'h009D; B = 16'h009C; #100;
A = 16'h009D; B = 16'h009D; #100;
A = 16'h009D; B = 16'h009E; #100;
A = 16'h009D; B = 16'h009F; #100;
A = 16'h009D; B = 16'h00A0; #100;
A = 16'h009D; B = 16'h00A1; #100;
A = 16'h009D; B = 16'h00A2; #100;
A = 16'h009D; B = 16'h00A3; #100;
A = 16'h009D; B = 16'h00A4; #100;
A = 16'h009D; B = 16'h00A5; #100;
A = 16'h009D; B = 16'h00A6; #100;
A = 16'h009D; B = 16'h00A7; #100;
A = 16'h009D; B = 16'h00A8; #100;
A = 16'h009D; B = 16'h00A9; #100;
A = 16'h009D; B = 16'h00AA; #100;
A = 16'h009D; B = 16'h00AB; #100;
A = 16'h009D; B = 16'h00AC; #100;
A = 16'h009D; B = 16'h00AD; #100;
A = 16'h009D; B = 16'h00AE; #100;
A = 16'h009D; B = 16'h00AF; #100;
A = 16'h009D; B = 16'h00B0; #100;
A = 16'h009D; B = 16'h00B1; #100;
A = 16'h009D; B = 16'h00B2; #100;
A = 16'h009D; B = 16'h00B3; #100;
A = 16'h009D; B = 16'h00B4; #100;
A = 16'h009D; B = 16'h00B5; #100;
A = 16'h009D; B = 16'h00B6; #100;
A = 16'h009D; B = 16'h00B7; #100;
A = 16'h009D; B = 16'h00B8; #100;
A = 16'h009D; B = 16'h00B9; #100;
A = 16'h009D; B = 16'h00BA; #100;
A = 16'h009D; B = 16'h00BB; #100;
A = 16'h009D; B = 16'h00BC; #100;
A = 16'h009D; B = 16'h00BD; #100;
A = 16'h009D; B = 16'h00BE; #100;
A = 16'h009D; B = 16'h00BF; #100;
A = 16'h009D; B = 16'h00C0; #100;
A = 16'h009D; B = 16'h00C1; #100;
A = 16'h009D; B = 16'h00C2; #100;
A = 16'h009D; B = 16'h00C3; #100;
A = 16'h009D; B = 16'h00C4; #100;
A = 16'h009D; B = 16'h00C5; #100;
A = 16'h009D; B = 16'h00C6; #100;
A = 16'h009D; B = 16'h00C7; #100;
A = 16'h009D; B = 16'h00C8; #100;
A = 16'h009D; B = 16'h00C9; #100;
A = 16'h009D; B = 16'h00CA; #100;
A = 16'h009D; B = 16'h00CB; #100;
A = 16'h009D; B = 16'h00CC; #100;
A = 16'h009D; B = 16'h00CD; #100;
A = 16'h009D; B = 16'h00CE; #100;
A = 16'h009D; B = 16'h00CF; #100;
A = 16'h009D; B = 16'h00D0; #100;
A = 16'h009D; B = 16'h00D1; #100;
A = 16'h009D; B = 16'h00D2; #100;
A = 16'h009D; B = 16'h00D3; #100;
A = 16'h009D; B = 16'h00D4; #100;
A = 16'h009D; B = 16'h00D5; #100;
A = 16'h009D; B = 16'h00D6; #100;
A = 16'h009D; B = 16'h00D7; #100;
A = 16'h009D; B = 16'h00D8; #100;
A = 16'h009D; B = 16'h00D9; #100;
A = 16'h009D; B = 16'h00DA; #100;
A = 16'h009D; B = 16'h00DB; #100;
A = 16'h009D; B = 16'h00DC; #100;
A = 16'h009D; B = 16'h00DD; #100;
A = 16'h009D; B = 16'h00DE; #100;
A = 16'h009D; B = 16'h00DF; #100;
A = 16'h009D; B = 16'h00E0; #100;
A = 16'h009D; B = 16'h00E1; #100;
A = 16'h009D; B = 16'h00E2; #100;
A = 16'h009D; B = 16'h00E3; #100;
A = 16'h009D; B = 16'h00E4; #100;
A = 16'h009D; B = 16'h00E5; #100;
A = 16'h009D; B = 16'h00E6; #100;
A = 16'h009D; B = 16'h00E7; #100;
A = 16'h009D; B = 16'h00E8; #100;
A = 16'h009D; B = 16'h00E9; #100;
A = 16'h009D; B = 16'h00EA; #100;
A = 16'h009D; B = 16'h00EB; #100;
A = 16'h009D; B = 16'h00EC; #100;
A = 16'h009D; B = 16'h00ED; #100;
A = 16'h009D; B = 16'h00EE; #100;
A = 16'h009D; B = 16'h00EF; #100;
A = 16'h009D; B = 16'h00F0; #100;
A = 16'h009D; B = 16'h00F1; #100;
A = 16'h009D; B = 16'h00F2; #100;
A = 16'h009D; B = 16'h00F3; #100;
A = 16'h009D; B = 16'h00F4; #100;
A = 16'h009D; B = 16'h00F5; #100;
A = 16'h009D; B = 16'h00F6; #100;
A = 16'h009D; B = 16'h00F7; #100;
A = 16'h009D; B = 16'h00F8; #100;
A = 16'h009D; B = 16'h00F9; #100;
A = 16'h009D; B = 16'h00FA; #100;
A = 16'h009D; B = 16'h00FB; #100;
A = 16'h009D; B = 16'h00FC; #100;
A = 16'h009D; B = 16'h00FD; #100;
A = 16'h009D; B = 16'h00FE; #100;
A = 16'h009D; B = 16'h00FF; #100;
A = 16'h009E; B = 16'h000; #100;
A = 16'h009E; B = 16'h001; #100;
A = 16'h009E; B = 16'h002; #100;
A = 16'h009E; B = 16'h003; #100;
A = 16'h009E; B = 16'h004; #100;
A = 16'h009E; B = 16'h005; #100;
A = 16'h009E; B = 16'h006; #100;
A = 16'h009E; B = 16'h007; #100;
A = 16'h009E; B = 16'h008; #100;
A = 16'h009E; B = 16'h009; #100;
A = 16'h009E; B = 16'h00A; #100;
A = 16'h009E; B = 16'h00B; #100;
A = 16'h009E; B = 16'h00C; #100;
A = 16'h009E; B = 16'h00D; #100;
A = 16'h009E; B = 16'h00E; #100;
A = 16'h009E; B = 16'h00F; #100;
A = 16'h009E; B = 16'h0010; #100;
A = 16'h009E; B = 16'h0011; #100;
A = 16'h009E; B = 16'h0012; #100;
A = 16'h009E; B = 16'h0013; #100;
A = 16'h009E; B = 16'h0014; #100;
A = 16'h009E; B = 16'h0015; #100;
A = 16'h009E; B = 16'h0016; #100;
A = 16'h009E; B = 16'h0017; #100;
A = 16'h009E; B = 16'h0018; #100;
A = 16'h009E; B = 16'h0019; #100;
A = 16'h009E; B = 16'h001A; #100;
A = 16'h009E; B = 16'h001B; #100;
A = 16'h009E; B = 16'h001C; #100;
A = 16'h009E; B = 16'h001D; #100;
A = 16'h009E; B = 16'h001E; #100;
A = 16'h009E; B = 16'h001F; #100;
A = 16'h009E; B = 16'h0020; #100;
A = 16'h009E; B = 16'h0021; #100;
A = 16'h009E; B = 16'h0022; #100;
A = 16'h009E; B = 16'h0023; #100;
A = 16'h009E; B = 16'h0024; #100;
A = 16'h009E; B = 16'h0025; #100;
A = 16'h009E; B = 16'h0026; #100;
A = 16'h009E; B = 16'h0027; #100;
A = 16'h009E; B = 16'h0028; #100;
A = 16'h009E; B = 16'h0029; #100;
A = 16'h009E; B = 16'h002A; #100;
A = 16'h009E; B = 16'h002B; #100;
A = 16'h009E; B = 16'h002C; #100;
A = 16'h009E; B = 16'h002D; #100;
A = 16'h009E; B = 16'h002E; #100;
A = 16'h009E; B = 16'h002F; #100;
A = 16'h009E; B = 16'h0030; #100;
A = 16'h009E; B = 16'h0031; #100;
A = 16'h009E; B = 16'h0032; #100;
A = 16'h009E; B = 16'h0033; #100;
A = 16'h009E; B = 16'h0034; #100;
A = 16'h009E; B = 16'h0035; #100;
A = 16'h009E; B = 16'h0036; #100;
A = 16'h009E; B = 16'h0037; #100;
A = 16'h009E; B = 16'h0038; #100;
A = 16'h009E; B = 16'h0039; #100;
A = 16'h009E; B = 16'h003A; #100;
A = 16'h009E; B = 16'h003B; #100;
A = 16'h009E; B = 16'h003C; #100;
A = 16'h009E; B = 16'h003D; #100;
A = 16'h009E; B = 16'h003E; #100;
A = 16'h009E; B = 16'h003F; #100;
A = 16'h009E; B = 16'h0040; #100;
A = 16'h009E; B = 16'h0041; #100;
A = 16'h009E; B = 16'h0042; #100;
A = 16'h009E; B = 16'h0043; #100;
A = 16'h009E; B = 16'h0044; #100;
A = 16'h009E; B = 16'h0045; #100;
A = 16'h009E; B = 16'h0046; #100;
A = 16'h009E; B = 16'h0047; #100;
A = 16'h009E; B = 16'h0048; #100;
A = 16'h009E; B = 16'h0049; #100;
A = 16'h009E; B = 16'h004A; #100;
A = 16'h009E; B = 16'h004B; #100;
A = 16'h009E; B = 16'h004C; #100;
A = 16'h009E; B = 16'h004D; #100;
A = 16'h009E; B = 16'h004E; #100;
A = 16'h009E; B = 16'h004F; #100;
A = 16'h009E; B = 16'h0050; #100;
A = 16'h009E; B = 16'h0051; #100;
A = 16'h009E; B = 16'h0052; #100;
A = 16'h009E; B = 16'h0053; #100;
A = 16'h009E; B = 16'h0054; #100;
A = 16'h009E; B = 16'h0055; #100;
A = 16'h009E; B = 16'h0056; #100;
A = 16'h009E; B = 16'h0057; #100;
A = 16'h009E; B = 16'h0058; #100;
A = 16'h009E; B = 16'h0059; #100;
A = 16'h009E; B = 16'h005A; #100;
A = 16'h009E; B = 16'h005B; #100;
A = 16'h009E; B = 16'h005C; #100;
A = 16'h009E; B = 16'h005D; #100;
A = 16'h009E; B = 16'h005E; #100;
A = 16'h009E; B = 16'h005F; #100;
A = 16'h009E; B = 16'h0060; #100;
A = 16'h009E; B = 16'h0061; #100;
A = 16'h009E; B = 16'h0062; #100;
A = 16'h009E; B = 16'h0063; #100;
A = 16'h009E; B = 16'h0064; #100;
A = 16'h009E; B = 16'h0065; #100;
A = 16'h009E; B = 16'h0066; #100;
A = 16'h009E; B = 16'h0067; #100;
A = 16'h009E; B = 16'h0068; #100;
A = 16'h009E; B = 16'h0069; #100;
A = 16'h009E; B = 16'h006A; #100;
A = 16'h009E; B = 16'h006B; #100;
A = 16'h009E; B = 16'h006C; #100;
A = 16'h009E; B = 16'h006D; #100;
A = 16'h009E; B = 16'h006E; #100;
A = 16'h009E; B = 16'h006F; #100;
A = 16'h009E; B = 16'h0070; #100;
A = 16'h009E; B = 16'h0071; #100;
A = 16'h009E; B = 16'h0072; #100;
A = 16'h009E; B = 16'h0073; #100;
A = 16'h009E; B = 16'h0074; #100;
A = 16'h009E; B = 16'h0075; #100;
A = 16'h009E; B = 16'h0076; #100;
A = 16'h009E; B = 16'h0077; #100;
A = 16'h009E; B = 16'h0078; #100;
A = 16'h009E; B = 16'h0079; #100;
A = 16'h009E; B = 16'h007A; #100;
A = 16'h009E; B = 16'h007B; #100;
A = 16'h009E; B = 16'h007C; #100;
A = 16'h009E; B = 16'h007D; #100;
A = 16'h009E; B = 16'h007E; #100;
A = 16'h009E; B = 16'h007F; #100;
A = 16'h009E; B = 16'h0080; #100;
A = 16'h009E; B = 16'h0081; #100;
A = 16'h009E; B = 16'h0082; #100;
A = 16'h009E; B = 16'h0083; #100;
A = 16'h009E; B = 16'h0084; #100;
A = 16'h009E; B = 16'h0085; #100;
A = 16'h009E; B = 16'h0086; #100;
A = 16'h009E; B = 16'h0087; #100;
A = 16'h009E; B = 16'h0088; #100;
A = 16'h009E; B = 16'h0089; #100;
A = 16'h009E; B = 16'h008A; #100;
A = 16'h009E; B = 16'h008B; #100;
A = 16'h009E; B = 16'h008C; #100;
A = 16'h009E; B = 16'h008D; #100;
A = 16'h009E; B = 16'h008E; #100;
A = 16'h009E; B = 16'h008F; #100;
A = 16'h009E; B = 16'h0090; #100;
A = 16'h009E; B = 16'h0091; #100;
A = 16'h009E; B = 16'h0092; #100;
A = 16'h009E; B = 16'h0093; #100;
A = 16'h009E; B = 16'h0094; #100;
A = 16'h009E; B = 16'h0095; #100;
A = 16'h009E; B = 16'h0096; #100;
A = 16'h009E; B = 16'h0097; #100;
A = 16'h009E; B = 16'h0098; #100;
A = 16'h009E; B = 16'h0099; #100;
A = 16'h009E; B = 16'h009A; #100;
A = 16'h009E; B = 16'h009B; #100;
A = 16'h009E; B = 16'h009C; #100;
A = 16'h009E; B = 16'h009D; #100;
A = 16'h009E; B = 16'h009E; #100;
A = 16'h009E; B = 16'h009F; #100;
A = 16'h009E; B = 16'h00A0; #100;
A = 16'h009E; B = 16'h00A1; #100;
A = 16'h009E; B = 16'h00A2; #100;
A = 16'h009E; B = 16'h00A3; #100;
A = 16'h009E; B = 16'h00A4; #100;
A = 16'h009E; B = 16'h00A5; #100;
A = 16'h009E; B = 16'h00A6; #100;
A = 16'h009E; B = 16'h00A7; #100;
A = 16'h009E; B = 16'h00A8; #100;
A = 16'h009E; B = 16'h00A9; #100;
A = 16'h009E; B = 16'h00AA; #100;
A = 16'h009E; B = 16'h00AB; #100;
A = 16'h009E; B = 16'h00AC; #100;
A = 16'h009E; B = 16'h00AD; #100;
A = 16'h009E; B = 16'h00AE; #100;
A = 16'h009E; B = 16'h00AF; #100;
A = 16'h009E; B = 16'h00B0; #100;
A = 16'h009E; B = 16'h00B1; #100;
A = 16'h009E; B = 16'h00B2; #100;
A = 16'h009E; B = 16'h00B3; #100;
A = 16'h009E; B = 16'h00B4; #100;
A = 16'h009E; B = 16'h00B5; #100;
A = 16'h009E; B = 16'h00B6; #100;
A = 16'h009E; B = 16'h00B7; #100;
A = 16'h009E; B = 16'h00B8; #100;
A = 16'h009E; B = 16'h00B9; #100;
A = 16'h009E; B = 16'h00BA; #100;
A = 16'h009E; B = 16'h00BB; #100;
A = 16'h009E; B = 16'h00BC; #100;
A = 16'h009E; B = 16'h00BD; #100;
A = 16'h009E; B = 16'h00BE; #100;
A = 16'h009E; B = 16'h00BF; #100;
A = 16'h009E; B = 16'h00C0; #100;
A = 16'h009E; B = 16'h00C1; #100;
A = 16'h009E; B = 16'h00C2; #100;
A = 16'h009E; B = 16'h00C3; #100;
A = 16'h009E; B = 16'h00C4; #100;
A = 16'h009E; B = 16'h00C5; #100;
A = 16'h009E; B = 16'h00C6; #100;
A = 16'h009E; B = 16'h00C7; #100;
A = 16'h009E; B = 16'h00C8; #100;
A = 16'h009E; B = 16'h00C9; #100;
A = 16'h009E; B = 16'h00CA; #100;
A = 16'h009E; B = 16'h00CB; #100;
A = 16'h009E; B = 16'h00CC; #100;
A = 16'h009E; B = 16'h00CD; #100;
A = 16'h009E; B = 16'h00CE; #100;
A = 16'h009E; B = 16'h00CF; #100;
A = 16'h009E; B = 16'h00D0; #100;
A = 16'h009E; B = 16'h00D1; #100;
A = 16'h009E; B = 16'h00D2; #100;
A = 16'h009E; B = 16'h00D3; #100;
A = 16'h009E; B = 16'h00D4; #100;
A = 16'h009E; B = 16'h00D5; #100;
A = 16'h009E; B = 16'h00D6; #100;
A = 16'h009E; B = 16'h00D7; #100;
A = 16'h009E; B = 16'h00D8; #100;
A = 16'h009E; B = 16'h00D9; #100;
A = 16'h009E; B = 16'h00DA; #100;
A = 16'h009E; B = 16'h00DB; #100;
A = 16'h009E; B = 16'h00DC; #100;
A = 16'h009E; B = 16'h00DD; #100;
A = 16'h009E; B = 16'h00DE; #100;
A = 16'h009E; B = 16'h00DF; #100;
A = 16'h009E; B = 16'h00E0; #100;
A = 16'h009E; B = 16'h00E1; #100;
A = 16'h009E; B = 16'h00E2; #100;
A = 16'h009E; B = 16'h00E3; #100;
A = 16'h009E; B = 16'h00E4; #100;
A = 16'h009E; B = 16'h00E5; #100;
A = 16'h009E; B = 16'h00E6; #100;
A = 16'h009E; B = 16'h00E7; #100;
A = 16'h009E; B = 16'h00E8; #100;
A = 16'h009E; B = 16'h00E9; #100;
A = 16'h009E; B = 16'h00EA; #100;
A = 16'h009E; B = 16'h00EB; #100;
A = 16'h009E; B = 16'h00EC; #100;
A = 16'h009E; B = 16'h00ED; #100;
A = 16'h009E; B = 16'h00EE; #100;
A = 16'h009E; B = 16'h00EF; #100;
A = 16'h009E; B = 16'h00F0; #100;
A = 16'h009E; B = 16'h00F1; #100;
A = 16'h009E; B = 16'h00F2; #100;
A = 16'h009E; B = 16'h00F3; #100;
A = 16'h009E; B = 16'h00F4; #100;
A = 16'h009E; B = 16'h00F5; #100;
A = 16'h009E; B = 16'h00F6; #100;
A = 16'h009E; B = 16'h00F7; #100;
A = 16'h009E; B = 16'h00F8; #100;
A = 16'h009E; B = 16'h00F9; #100;
A = 16'h009E; B = 16'h00FA; #100;
A = 16'h009E; B = 16'h00FB; #100;
A = 16'h009E; B = 16'h00FC; #100;
A = 16'h009E; B = 16'h00FD; #100;
A = 16'h009E; B = 16'h00FE; #100;
A = 16'h009E; B = 16'h00FF; #100;
A = 16'h009F; B = 16'h000; #100;
A = 16'h009F; B = 16'h001; #100;
A = 16'h009F; B = 16'h002; #100;
A = 16'h009F; B = 16'h003; #100;
A = 16'h009F; B = 16'h004; #100;
A = 16'h009F; B = 16'h005; #100;
A = 16'h009F; B = 16'h006; #100;
A = 16'h009F; B = 16'h007; #100;
A = 16'h009F; B = 16'h008; #100;
A = 16'h009F; B = 16'h009; #100;
A = 16'h009F; B = 16'h00A; #100;
A = 16'h009F; B = 16'h00B; #100;
A = 16'h009F; B = 16'h00C; #100;
A = 16'h009F; B = 16'h00D; #100;
A = 16'h009F; B = 16'h00E; #100;
A = 16'h009F; B = 16'h00F; #100;
A = 16'h009F; B = 16'h0010; #100;
A = 16'h009F; B = 16'h0011; #100;
A = 16'h009F; B = 16'h0012; #100;
A = 16'h009F; B = 16'h0013; #100;
A = 16'h009F; B = 16'h0014; #100;
A = 16'h009F; B = 16'h0015; #100;
A = 16'h009F; B = 16'h0016; #100;
A = 16'h009F; B = 16'h0017; #100;
A = 16'h009F; B = 16'h0018; #100;
A = 16'h009F; B = 16'h0019; #100;
A = 16'h009F; B = 16'h001A; #100;
A = 16'h009F; B = 16'h001B; #100;
A = 16'h009F; B = 16'h001C; #100;
A = 16'h009F; B = 16'h001D; #100;
A = 16'h009F; B = 16'h001E; #100;
A = 16'h009F; B = 16'h001F; #100;
A = 16'h009F; B = 16'h0020; #100;
A = 16'h009F; B = 16'h0021; #100;
A = 16'h009F; B = 16'h0022; #100;
A = 16'h009F; B = 16'h0023; #100;
A = 16'h009F; B = 16'h0024; #100;
A = 16'h009F; B = 16'h0025; #100;
A = 16'h009F; B = 16'h0026; #100;
A = 16'h009F; B = 16'h0027; #100;
A = 16'h009F; B = 16'h0028; #100;
A = 16'h009F; B = 16'h0029; #100;
A = 16'h009F; B = 16'h002A; #100;
A = 16'h009F; B = 16'h002B; #100;
A = 16'h009F; B = 16'h002C; #100;
A = 16'h009F; B = 16'h002D; #100;
A = 16'h009F; B = 16'h002E; #100;
A = 16'h009F; B = 16'h002F; #100;
A = 16'h009F; B = 16'h0030; #100;
A = 16'h009F; B = 16'h0031; #100;
A = 16'h009F; B = 16'h0032; #100;
A = 16'h009F; B = 16'h0033; #100;
A = 16'h009F; B = 16'h0034; #100;
A = 16'h009F; B = 16'h0035; #100;
A = 16'h009F; B = 16'h0036; #100;
A = 16'h009F; B = 16'h0037; #100;
A = 16'h009F; B = 16'h0038; #100;
A = 16'h009F; B = 16'h0039; #100;
A = 16'h009F; B = 16'h003A; #100;
A = 16'h009F; B = 16'h003B; #100;
A = 16'h009F; B = 16'h003C; #100;
A = 16'h009F; B = 16'h003D; #100;
A = 16'h009F; B = 16'h003E; #100;
A = 16'h009F; B = 16'h003F; #100;
A = 16'h009F; B = 16'h0040; #100;
A = 16'h009F; B = 16'h0041; #100;
A = 16'h009F; B = 16'h0042; #100;
A = 16'h009F; B = 16'h0043; #100;
A = 16'h009F; B = 16'h0044; #100;
A = 16'h009F; B = 16'h0045; #100;
A = 16'h009F; B = 16'h0046; #100;
A = 16'h009F; B = 16'h0047; #100;
A = 16'h009F; B = 16'h0048; #100;
A = 16'h009F; B = 16'h0049; #100;
A = 16'h009F; B = 16'h004A; #100;
A = 16'h009F; B = 16'h004B; #100;
A = 16'h009F; B = 16'h004C; #100;
A = 16'h009F; B = 16'h004D; #100;
A = 16'h009F; B = 16'h004E; #100;
A = 16'h009F; B = 16'h004F; #100;
A = 16'h009F; B = 16'h0050; #100;
A = 16'h009F; B = 16'h0051; #100;
A = 16'h009F; B = 16'h0052; #100;
A = 16'h009F; B = 16'h0053; #100;
A = 16'h009F; B = 16'h0054; #100;
A = 16'h009F; B = 16'h0055; #100;
A = 16'h009F; B = 16'h0056; #100;
A = 16'h009F; B = 16'h0057; #100;
A = 16'h009F; B = 16'h0058; #100;
A = 16'h009F; B = 16'h0059; #100;
A = 16'h009F; B = 16'h005A; #100;
A = 16'h009F; B = 16'h005B; #100;
A = 16'h009F; B = 16'h005C; #100;
A = 16'h009F; B = 16'h005D; #100;
A = 16'h009F; B = 16'h005E; #100;
A = 16'h009F; B = 16'h005F; #100;
A = 16'h009F; B = 16'h0060; #100;
A = 16'h009F; B = 16'h0061; #100;
A = 16'h009F; B = 16'h0062; #100;
A = 16'h009F; B = 16'h0063; #100;
A = 16'h009F; B = 16'h0064; #100;
A = 16'h009F; B = 16'h0065; #100;
A = 16'h009F; B = 16'h0066; #100;
A = 16'h009F; B = 16'h0067; #100;
A = 16'h009F; B = 16'h0068; #100;
A = 16'h009F; B = 16'h0069; #100;
A = 16'h009F; B = 16'h006A; #100;
A = 16'h009F; B = 16'h006B; #100;
A = 16'h009F; B = 16'h006C; #100;
A = 16'h009F; B = 16'h006D; #100;
A = 16'h009F; B = 16'h006E; #100;
A = 16'h009F; B = 16'h006F; #100;
A = 16'h009F; B = 16'h0070; #100;
A = 16'h009F; B = 16'h0071; #100;
A = 16'h009F; B = 16'h0072; #100;
A = 16'h009F; B = 16'h0073; #100;
A = 16'h009F; B = 16'h0074; #100;
A = 16'h009F; B = 16'h0075; #100;
A = 16'h009F; B = 16'h0076; #100;
A = 16'h009F; B = 16'h0077; #100;
A = 16'h009F; B = 16'h0078; #100;
A = 16'h009F; B = 16'h0079; #100;
A = 16'h009F; B = 16'h007A; #100;
A = 16'h009F; B = 16'h007B; #100;
A = 16'h009F; B = 16'h007C; #100;
A = 16'h009F; B = 16'h007D; #100;
A = 16'h009F; B = 16'h007E; #100;
A = 16'h009F; B = 16'h007F; #100;
A = 16'h009F; B = 16'h0080; #100;
A = 16'h009F; B = 16'h0081; #100;
A = 16'h009F; B = 16'h0082; #100;
A = 16'h009F; B = 16'h0083; #100;
A = 16'h009F; B = 16'h0084; #100;
A = 16'h009F; B = 16'h0085; #100;
A = 16'h009F; B = 16'h0086; #100;
A = 16'h009F; B = 16'h0087; #100;
A = 16'h009F; B = 16'h0088; #100;
A = 16'h009F; B = 16'h0089; #100;
A = 16'h009F; B = 16'h008A; #100;
A = 16'h009F; B = 16'h008B; #100;
A = 16'h009F; B = 16'h008C; #100;
A = 16'h009F; B = 16'h008D; #100;
A = 16'h009F; B = 16'h008E; #100;
A = 16'h009F; B = 16'h008F; #100;
A = 16'h009F; B = 16'h0090; #100;
A = 16'h009F; B = 16'h0091; #100;
A = 16'h009F; B = 16'h0092; #100;
A = 16'h009F; B = 16'h0093; #100;
A = 16'h009F; B = 16'h0094; #100;
A = 16'h009F; B = 16'h0095; #100;
A = 16'h009F; B = 16'h0096; #100;
A = 16'h009F; B = 16'h0097; #100;
A = 16'h009F; B = 16'h0098; #100;
A = 16'h009F; B = 16'h0099; #100;
A = 16'h009F; B = 16'h009A; #100;
A = 16'h009F; B = 16'h009B; #100;
A = 16'h009F; B = 16'h009C; #100;
A = 16'h009F; B = 16'h009D; #100;
A = 16'h009F; B = 16'h009E; #100;
A = 16'h009F; B = 16'h009F; #100;
A = 16'h009F; B = 16'h00A0; #100;
A = 16'h009F; B = 16'h00A1; #100;
A = 16'h009F; B = 16'h00A2; #100;
A = 16'h009F; B = 16'h00A3; #100;
A = 16'h009F; B = 16'h00A4; #100;
A = 16'h009F; B = 16'h00A5; #100;
A = 16'h009F; B = 16'h00A6; #100;
A = 16'h009F; B = 16'h00A7; #100;
A = 16'h009F; B = 16'h00A8; #100;
A = 16'h009F; B = 16'h00A9; #100;
A = 16'h009F; B = 16'h00AA; #100;
A = 16'h009F; B = 16'h00AB; #100;
A = 16'h009F; B = 16'h00AC; #100;
A = 16'h009F; B = 16'h00AD; #100;
A = 16'h009F; B = 16'h00AE; #100;
A = 16'h009F; B = 16'h00AF; #100;
A = 16'h009F; B = 16'h00B0; #100;
A = 16'h009F; B = 16'h00B1; #100;
A = 16'h009F; B = 16'h00B2; #100;
A = 16'h009F; B = 16'h00B3; #100;
A = 16'h009F; B = 16'h00B4; #100;
A = 16'h009F; B = 16'h00B5; #100;
A = 16'h009F; B = 16'h00B6; #100;
A = 16'h009F; B = 16'h00B7; #100;
A = 16'h009F; B = 16'h00B8; #100;
A = 16'h009F; B = 16'h00B9; #100;
A = 16'h009F; B = 16'h00BA; #100;
A = 16'h009F; B = 16'h00BB; #100;
A = 16'h009F; B = 16'h00BC; #100;
A = 16'h009F; B = 16'h00BD; #100;
A = 16'h009F; B = 16'h00BE; #100;
A = 16'h009F; B = 16'h00BF; #100;
A = 16'h009F; B = 16'h00C0; #100;
A = 16'h009F; B = 16'h00C1; #100;
A = 16'h009F; B = 16'h00C2; #100;
A = 16'h009F; B = 16'h00C3; #100;
A = 16'h009F; B = 16'h00C4; #100;
A = 16'h009F; B = 16'h00C5; #100;
A = 16'h009F; B = 16'h00C6; #100;
A = 16'h009F; B = 16'h00C7; #100;
A = 16'h009F; B = 16'h00C8; #100;
A = 16'h009F; B = 16'h00C9; #100;
A = 16'h009F; B = 16'h00CA; #100;
A = 16'h009F; B = 16'h00CB; #100;
A = 16'h009F; B = 16'h00CC; #100;
A = 16'h009F; B = 16'h00CD; #100;
A = 16'h009F; B = 16'h00CE; #100;
A = 16'h009F; B = 16'h00CF; #100;
A = 16'h009F; B = 16'h00D0; #100;
A = 16'h009F; B = 16'h00D1; #100;
A = 16'h009F; B = 16'h00D2; #100;
A = 16'h009F; B = 16'h00D3; #100;
A = 16'h009F; B = 16'h00D4; #100;
A = 16'h009F; B = 16'h00D5; #100;
A = 16'h009F; B = 16'h00D6; #100;
A = 16'h009F; B = 16'h00D7; #100;
A = 16'h009F; B = 16'h00D8; #100;
A = 16'h009F; B = 16'h00D9; #100;
A = 16'h009F; B = 16'h00DA; #100;
A = 16'h009F; B = 16'h00DB; #100;
A = 16'h009F; B = 16'h00DC; #100;
A = 16'h009F; B = 16'h00DD; #100;
A = 16'h009F; B = 16'h00DE; #100;
A = 16'h009F; B = 16'h00DF; #100;
A = 16'h009F; B = 16'h00E0; #100;
A = 16'h009F; B = 16'h00E1; #100;
A = 16'h009F; B = 16'h00E2; #100;
A = 16'h009F; B = 16'h00E3; #100;
A = 16'h009F; B = 16'h00E4; #100;
A = 16'h009F; B = 16'h00E5; #100;
A = 16'h009F; B = 16'h00E6; #100;
A = 16'h009F; B = 16'h00E7; #100;
A = 16'h009F; B = 16'h00E8; #100;
A = 16'h009F; B = 16'h00E9; #100;
A = 16'h009F; B = 16'h00EA; #100;
A = 16'h009F; B = 16'h00EB; #100;
A = 16'h009F; B = 16'h00EC; #100;
A = 16'h009F; B = 16'h00ED; #100;
A = 16'h009F; B = 16'h00EE; #100;
A = 16'h009F; B = 16'h00EF; #100;
A = 16'h009F; B = 16'h00F0; #100;
A = 16'h009F; B = 16'h00F1; #100;
A = 16'h009F; B = 16'h00F2; #100;
A = 16'h009F; B = 16'h00F3; #100;
A = 16'h009F; B = 16'h00F4; #100;
A = 16'h009F; B = 16'h00F5; #100;
A = 16'h009F; B = 16'h00F6; #100;
A = 16'h009F; B = 16'h00F7; #100;
A = 16'h009F; B = 16'h00F8; #100;
A = 16'h009F; B = 16'h00F9; #100;
A = 16'h009F; B = 16'h00FA; #100;
A = 16'h009F; B = 16'h00FB; #100;
A = 16'h009F; B = 16'h00FC; #100;
A = 16'h009F; B = 16'h00FD; #100;
A = 16'h009F; B = 16'h00FE; #100;
A = 16'h009F; B = 16'h00FF; #100;
A = 16'h00A0; B = 16'h000; #100;
A = 16'h00A0; B = 16'h001; #100;
A = 16'h00A0; B = 16'h002; #100;
A = 16'h00A0; B = 16'h003; #100;
A = 16'h00A0; B = 16'h004; #100;
A = 16'h00A0; B = 16'h005; #100;
A = 16'h00A0; B = 16'h006; #100;
A = 16'h00A0; B = 16'h007; #100;
A = 16'h00A0; B = 16'h008; #100;
A = 16'h00A0; B = 16'h009; #100;
A = 16'h00A0; B = 16'h00A; #100;
A = 16'h00A0; B = 16'h00B; #100;
A = 16'h00A0; B = 16'h00C; #100;
A = 16'h00A0; B = 16'h00D; #100;
A = 16'h00A0; B = 16'h00E; #100;
A = 16'h00A0; B = 16'h00F; #100;
A = 16'h00A0; B = 16'h0010; #100;
A = 16'h00A0; B = 16'h0011; #100;
A = 16'h00A0; B = 16'h0012; #100;
A = 16'h00A0; B = 16'h0013; #100;
A = 16'h00A0; B = 16'h0014; #100;
A = 16'h00A0; B = 16'h0015; #100;
A = 16'h00A0; B = 16'h0016; #100;
A = 16'h00A0; B = 16'h0017; #100;
A = 16'h00A0; B = 16'h0018; #100;
A = 16'h00A0; B = 16'h0019; #100;
A = 16'h00A0; B = 16'h001A; #100;
A = 16'h00A0; B = 16'h001B; #100;
A = 16'h00A0; B = 16'h001C; #100;
A = 16'h00A0; B = 16'h001D; #100;
A = 16'h00A0; B = 16'h001E; #100;
A = 16'h00A0; B = 16'h001F; #100;
A = 16'h00A0; B = 16'h0020; #100;
A = 16'h00A0; B = 16'h0021; #100;
A = 16'h00A0; B = 16'h0022; #100;
A = 16'h00A0; B = 16'h0023; #100;
A = 16'h00A0; B = 16'h0024; #100;
A = 16'h00A0; B = 16'h0025; #100;
A = 16'h00A0; B = 16'h0026; #100;
A = 16'h00A0; B = 16'h0027; #100;
A = 16'h00A0; B = 16'h0028; #100;
A = 16'h00A0; B = 16'h0029; #100;
A = 16'h00A0; B = 16'h002A; #100;
A = 16'h00A0; B = 16'h002B; #100;
A = 16'h00A0; B = 16'h002C; #100;
A = 16'h00A0; B = 16'h002D; #100;
A = 16'h00A0; B = 16'h002E; #100;
A = 16'h00A0; B = 16'h002F; #100;
A = 16'h00A0; B = 16'h0030; #100;
A = 16'h00A0; B = 16'h0031; #100;
A = 16'h00A0; B = 16'h0032; #100;
A = 16'h00A0; B = 16'h0033; #100;
A = 16'h00A0; B = 16'h0034; #100;
A = 16'h00A0; B = 16'h0035; #100;
A = 16'h00A0; B = 16'h0036; #100;
A = 16'h00A0; B = 16'h0037; #100;
A = 16'h00A0; B = 16'h0038; #100;
A = 16'h00A0; B = 16'h0039; #100;
A = 16'h00A0; B = 16'h003A; #100;
A = 16'h00A0; B = 16'h003B; #100;
A = 16'h00A0; B = 16'h003C; #100;
A = 16'h00A0; B = 16'h003D; #100;
A = 16'h00A0; B = 16'h003E; #100;
A = 16'h00A0; B = 16'h003F; #100;
A = 16'h00A0; B = 16'h0040; #100;
A = 16'h00A0; B = 16'h0041; #100;
A = 16'h00A0; B = 16'h0042; #100;
A = 16'h00A0; B = 16'h0043; #100;
A = 16'h00A0; B = 16'h0044; #100;
A = 16'h00A0; B = 16'h0045; #100;
A = 16'h00A0; B = 16'h0046; #100;
A = 16'h00A0; B = 16'h0047; #100;
A = 16'h00A0; B = 16'h0048; #100;
A = 16'h00A0; B = 16'h0049; #100;
A = 16'h00A0; B = 16'h004A; #100;
A = 16'h00A0; B = 16'h004B; #100;
A = 16'h00A0; B = 16'h004C; #100;
A = 16'h00A0; B = 16'h004D; #100;
A = 16'h00A0; B = 16'h004E; #100;
A = 16'h00A0; B = 16'h004F; #100;
A = 16'h00A0; B = 16'h0050; #100;
A = 16'h00A0; B = 16'h0051; #100;
A = 16'h00A0; B = 16'h0052; #100;
A = 16'h00A0; B = 16'h0053; #100;
A = 16'h00A0; B = 16'h0054; #100;
A = 16'h00A0; B = 16'h0055; #100;
A = 16'h00A0; B = 16'h0056; #100;
A = 16'h00A0; B = 16'h0057; #100;
A = 16'h00A0; B = 16'h0058; #100;
A = 16'h00A0; B = 16'h0059; #100;
A = 16'h00A0; B = 16'h005A; #100;
A = 16'h00A0; B = 16'h005B; #100;
A = 16'h00A0; B = 16'h005C; #100;
A = 16'h00A0; B = 16'h005D; #100;
A = 16'h00A0; B = 16'h005E; #100;
A = 16'h00A0; B = 16'h005F; #100;
A = 16'h00A0; B = 16'h0060; #100;
A = 16'h00A0; B = 16'h0061; #100;
A = 16'h00A0; B = 16'h0062; #100;
A = 16'h00A0; B = 16'h0063; #100;
A = 16'h00A0; B = 16'h0064; #100;
A = 16'h00A0; B = 16'h0065; #100;
A = 16'h00A0; B = 16'h0066; #100;
A = 16'h00A0; B = 16'h0067; #100;
A = 16'h00A0; B = 16'h0068; #100;
A = 16'h00A0; B = 16'h0069; #100;
A = 16'h00A0; B = 16'h006A; #100;
A = 16'h00A0; B = 16'h006B; #100;
A = 16'h00A0; B = 16'h006C; #100;
A = 16'h00A0; B = 16'h006D; #100;
A = 16'h00A0; B = 16'h006E; #100;
A = 16'h00A0; B = 16'h006F; #100;
A = 16'h00A0; B = 16'h0070; #100;
A = 16'h00A0; B = 16'h0071; #100;
A = 16'h00A0; B = 16'h0072; #100;
A = 16'h00A0; B = 16'h0073; #100;
A = 16'h00A0; B = 16'h0074; #100;
A = 16'h00A0; B = 16'h0075; #100;
A = 16'h00A0; B = 16'h0076; #100;
A = 16'h00A0; B = 16'h0077; #100;
A = 16'h00A0; B = 16'h0078; #100;
A = 16'h00A0; B = 16'h0079; #100;
A = 16'h00A0; B = 16'h007A; #100;
A = 16'h00A0; B = 16'h007B; #100;
A = 16'h00A0; B = 16'h007C; #100;
A = 16'h00A0; B = 16'h007D; #100;
A = 16'h00A0; B = 16'h007E; #100;
A = 16'h00A0; B = 16'h007F; #100;
A = 16'h00A0; B = 16'h0080; #100;
A = 16'h00A0; B = 16'h0081; #100;
A = 16'h00A0; B = 16'h0082; #100;
A = 16'h00A0; B = 16'h0083; #100;
A = 16'h00A0; B = 16'h0084; #100;
A = 16'h00A0; B = 16'h0085; #100;
A = 16'h00A0; B = 16'h0086; #100;
A = 16'h00A0; B = 16'h0087; #100;
A = 16'h00A0; B = 16'h0088; #100;
A = 16'h00A0; B = 16'h0089; #100;
A = 16'h00A0; B = 16'h008A; #100;
A = 16'h00A0; B = 16'h008B; #100;
A = 16'h00A0; B = 16'h008C; #100;
A = 16'h00A0; B = 16'h008D; #100;
A = 16'h00A0; B = 16'h008E; #100;
A = 16'h00A0; B = 16'h008F; #100;
A = 16'h00A0; B = 16'h0090; #100;
A = 16'h00A0; B = 16'h0091; #100;
A = 16'h00A0; B = 16'h0092; #100;
A = 16'h00A0; B = 16'h0093; #100;
A = 16'h00A0; B = 16'h0094; #100;
A = 16'h00A0; B = 16'h0095; #100;
A = 16'h00A0; B = 16'h0096; #100;
A = 16'h00A0; B = 16'h0097; #100;
A = 16'h00A0; B = 16'h0098; #100;
A = 16'h00A0; B = 16'h0099; #100;
A = 16'h00A0; B = 16'h009A; #100;
A = 16'h00A0; B = 16'h009B; #100;
A = 16'h00A0; B = 16'h009C; #100;
A = 16'h00A0; B = 16'h009D; #100;
A = 16'h00A0; B = 16'h009E; #100;
A = 16'h00A0; B = 16'h009F; #100;
A = 16'h00A0; B = 16'h00A0; #100;
A = 16'h00A0; B = 16'h00A1; #100;
A = 16'h00A0; B = 16'h00A2; #100;
A = 16'h00A0; B = 16'h00A3; #100;
A = 16'h00A0; B = 16'h00A4; #100;
A = 16'h00A0; B = 16'h00A5; #100;
A = 16'h00A0; B = 16'h00A6; #100;
A = 16'h00A0; B = 16'h00A7; #100;
A = 16'h00A0; B = 16'h00A8; #100;
A = 16'h00A0; B = 16'h00A9; #100;
A = 16'h00A0; B = 16'h00AA; #100;
A = 16'h00A0; B = 16'h00AB; #100;
A = 16'h00A0; B = 16'h00AC; #100;
A = 16'h00A0; B = 16'h00AD; #100;
A = 16'h00A0; B = 16'h00AE; #100;
A = 16'h00A0; B = 16'h00AF; #100;
A = 16'h00A0; B = 16'h00B0; #100;
A = 16'h00A0; B = 16'h00B1; #100;
A = 16'h00A0; B = 16'h00B2; #100;
A = 16'h00A0; B = 16'h00B3; #100;
A = 16'h00A0; B = 16'h00B4; #100;
A = 16'h00A0; B = 16'h00B5; #100;
A = 16'h00A0; B = 16'h00B6; #100;
A = 16'h00A0; B = 16'h00B7; #100;
A = 16'h00A0; B = 16'h00B8; #100;
A = 16'h00A0; B = 16'h00B9; #100;
A = 16'h00A0; B = 16'h00BA; #100;
A = 16'h00A0; B = 16'h00BB; #100;
A = 16'h00A0; B = 16'h00BC; #100;
A = 16'h00A0; B = 16'h00BD; #100;
A = 16'h00A0; B = 16'h00BE; #100;
A = 16'h00A0; B = 16'h00BF; #100;
A = 16'h00A0; B = 16'h00C0; #100;
A = 16'h00A0; B = 16'h00C1; #100;
A = 16'h00A0; B = 16'h00C2; #100;
A = 16'h00A0; B = 16'h00C3; #100;
A = 16'h00A0; B = 16'h00C4; #100;
A = 16'h00A0; B = 16'h00C5; #100;
A = 16'h00A0; B = 16'h00C6; #100;
A = 16'h00A0; B = 16'h00C7; #100;
A = 16'h00A0; B = 16'h00C8; #100;
A = 16'h00A0; B = 16'h00C9; #100;
A = 16'h00A0; B = 16'h00CA; #100;
A = 16'h00A0; B = 16'h00CB; #100;
A = 16'h00A0; B = 16'h00CC; #100;
A = 16'h00A0; B = 16'h00CD; #100;
A = 16'h00A0; B = 16'h00CE; #100;
A = 16'h00A0; B = 16'h00CF; #100;
A = 16'h00A0; B = 16'h00D0; #100;
A = 16'h00A0; B = 16'h00D1; #100;
A = 16'h00A0; B = 16'h00D2; #100;
A = 16'h00A0; B = 16'h00D3; #100;
A = 16'h00A0; B = 16'h00D4; #100;
A = 16'h00A0; B = 16'h00D5; #100;
A = 16'h00A0; B = 16'h00D6; #100;
A = 16'h00A0; B = 16'h00D7; #100;
A = 16'h00A0; B = 16'h00D8; #100;
A = 16'h00A0; B = 16'h00D9; #100;
A = 16'h00A0; B = 16'h00DA; #100;
A = 16'h00A0; B = 16'h00DB; #100;
A = 16'h00A0; B = 16'h00DC; #100;
A = 16'h00A0; B = 16'h00DD; #100;
A = 16'h00A0; B = 16'h00DE; #100;
A = 16'h00A0; B = 16'h00DF; #100;
A = 16'h00A0; B = 16'h00E0; #100;
A = 16'h00A0; B = 16'h00E1; #100;
A = 16'h00A0; B = 16'h00E2; #100;
A = 16'h00A0; B = 16'h00E3; #100;
A = 16'h00A0; B = 16'h00E4; #100;
A = 16'h00A0; B = 16'h00E5; #100;
A = 16'h00A0; B = 16'h00E6; #100;
A = 16'h00A0; B = 16'h00E7; #100;
A = 16'h00A0; B = 16'h00E8; #100;
A = 16'h00A0; B = 16'h00E9; #100;
A = 16'h00A0; B = 16'h00EA; #100;
A = 16'h00A0; B = 16'h00EB; #100;
A = 16'h00A0; B = 16'h00EC; #100;
A = 16'h00A0; B = 16'h00ED; #100;
A = 16'h00A0; B = 16'h00EE; #100;
A = 16'h00A0; B = 16'h00EF; #100;
A = 16'h00A0; B = 16'h00F0; #100;
A = 16'h00A0; B = 16'h00F1; #100;
A = 16'h00A0; B = 16'h00F2; #100;
A = 16'h00A0; B = 16'h00F3; #100;
A = 16'h00A0; B = 16'h00F4; #100;
A = 16'h00A0; B = 16'h00F5; #100;
A = 16'h00A0; B = 16'h00F6; #100;
A = 16'h00A0; B = 16'h00F7; #100;
A = 16'h00A0; B = 16'h00F8; #100;
A = 16'h00A0; B = 16'h00F9; #100;
A = 16'h00A0; B = 16'h00FA; #100;
A = 16'h00A0; B = 16'h00FB; #100;
A = 16'h00A0; B = 16'h00FC; #100;
A = 16'h00A0; B = 16'h00FD; #100;
A = 16'h00A0; B = 16'h00FE; #100;
A = 16'h00A0; B = 16'h00FF; #100;
A = 16'h00A1; B = 16'h000; #100;
A = 16'h00A1; B = 16'h001; #100;
A = 16'h00A1; B = 16'h002; #100;
A = 16'h00A1; B = 16'h003; #100;
A = 16'h00A1; B = 16'h004; #100;
A = 16'h00A1; B = 16'h005; #100;
A = 16'h00A1; B = 16'h006; #100;
A = 16'h00A1; B = 16'h007; #100;
A = 16'h00A1; B = 16'h008; #100;
A = 16'h00A1; B = 16'h009; #100;
A = 16'h00A1; B = 16'h00A; #100;
A = 16'h00A1; B = 16'h00B; #100;
A = 16'h00A1; B = 16'h00C; #100;
A = 16'h00A1; B = 16'h00D; #100;
A = 16'h00A1; B = 16'h00E; #100;
A = 16'h00A1; B = 16'h00F; #100;
A = 16'h00A1; B = 16'h0010; #100;
A = 16'h00A1; B = 16'h0011; #100;
A = 16'h00A1; B = 16'h0012; #100;
A = 16'h00A1; B = 16'h0013; #100;
A = 16'h00A1; B = 16'h0014; #100;
A = 16'h00A1; B = 16'h0015; #100;
A = 16'h00A1; B = 16'h0016; #100;
A = 16'h00A1; B = 16'h0017; #100;
A = 16'h00A1; B = 16'h0018; #100;
A = 16'h00A1; B = 16'h0019; #100;
A = 16'h00A1; B = 16'h001A; #100;
A = 16'h00A1; B = 16'h001B; #100;
A = 16'h00A1; B = 16'h001C; #100;
A = 16'h00A1; B = 16'h001D; #100;
A = 16'h00A1; B = 16'h001E; #100;
A = 16'h00A1; B = 16'h001F; #100;
A = 16'h00A1; B = 16'h0020; #100;
A = 16'h00A1; B = 16'h0021; #100;
A = 16'h00A1; B = 16'h0022; #100;
A = 16'h00A1; B = 16'h0023; #100;
A = 16'h00A1; B = 16'h0024; #100;
A = 16'h00A1; B = 16'h0025; #100;
A = 16'h00A1; B = 16'h0026; #100;
A = 16'h00A1; B = 16'h0027; #100;
A = 16'h00A1; B = 16'h0028; #100;
A = 16'h00A1; B = 16'h0029; #100;
A = 16'h00A1; B = 16'h002A; #100;
A = 16'h00A1; B = 16'h002B; #100;
A = 16'h00A1; B = 16'h002C; #100;
A = 16'h00A1; B = 16'h002D; #100;
A = 16'h00A1; B = 16'h002E; #100;
A = 16'h00A1; B = 16'h002F; #100;
A = 16'h00A1; B = 16'h0030; #100;
A = 16'h00A1; B = 16'h0031; #100;
A = 16'h00A1; B = 16'h0032; #100;
A = 16'h00A1; B = 16'h0033; #100;
A = 16'h00A1; B = 16'h0034; #100;
A = 16'h00A1; B = 16'h0035; #100;
A = 16'h00A1; B = 16'h0036; #100;
A = 16'h00A1; B = 16'h0037; #100;
A = 16'h00A1; B = 16'h0038; #100;
A = 16'h00A1; B = 16'h0039; #100;
A = 16'h00A1; B = 16'h003A; #100;
A = 16'h00A1; B = 16'h003B; #100;
A = 16'h00A1; B = 16'h003C; #100;
A = 16'h00A1; B = 16'h003D; #100;
A = 16'h00A1; B = 16'h003E; #100;
A = 16'h00A1; B = 16'h003F; #100;
A = 16'h00A1; B = 16'h0040; #100;
A = 16'h00A1; B = 16'h0041; #100;
A = 16'h00A1; B = 16'h0042; #100;
A = 16'h00A1; B = 16'h0043; #100;
A = 16'h00A1; B = 16'h0044; #100;
A = 16'h00A1; B = 16'h0045; #100;
A = 16'h00A1; B = 16'h0046; #100;
A = 16'h00A1; B = 16'h0047; #100;
A = 16'h00A1; B = 16'h0048; #100;
A = 16'h00A1; B = 16'h0049; #100;
A = 16'h00A1; B = 16'h004A; #100;
A = 16'h00A1; B = 16'h004B; #100;
A = 16'h00A1; B = 16'h004C; #100;
A = 16'h00A1; B = 16'h004D; #100;
A = 16'h00A1; B = 16'h004E; #100;
A = 16'h00A1; B = 16'h004F; #100;
A = 16'h00A1; B = 16'h0050; #100;
A = 16'h00A1; B = 16'h0051; #100;
A = 16'h00A1; B = 16'h0052; #100;
A = 16'h00A1; B = 16'h0053; #100;
A = 16'h00A1; B = 16'h0054; #100;
A = 16'h00A1; B = 16'h0055; #100;
A = 16'h00A1; B = 16'h0056; #100;
A = 16'h00A1; B = 16'h0057; #100;
A = 16'h00A1; B = 16'h0058; #100;
A = 16'h00A1; B = 16'h0059; #100;
A = 16'h00A1; B = 16'h005A; #100;
A = 16'h00A1; B = 16'h005B; #100;
A = 16'h00A1; B = 16'h005C; #100;
A = 16'h00A1; B = 16'h005D; #100;
A = 16'h00A1; B = 16'h005E; #100;
A = 16'h00A1; B = 16'h005F; #100;
A = 16'h00A1; B = 16'h0060; #100;
A = 16'h00A1; B = 16'h0061; #100;
A = 16'h00A1; B = 16'h0062; #100;
A = 16'h00A1; B = 16'h0063; #100;
A = 16'h00A1; B = 16'h0064; #100;
A = 16'h00A1; B = 16'h0065; #100;
A = 16'h00A1; B = 16'h0066; #100;
A = 16'h00A1; B = 16'h0067; #100;
A = 16'h00A1; B = 16'h0068; #100;
A = 16'h00A1; B = 16'h0069; #100;
A = 16'h00A1; B = 16'h006A; #100;
A = 16'h00A1; B = 16'h006B; #100;
A = 16'h00A1; B = 16'h006C; #100;
A = 16'h00A1; B = 16'h006D; #100;
A = 16'h00A1; B = 16'h006E; #100;
A = 16'h00A1; B = 16'h006F; #100;
A = 16'h00A1; B = 16'h0070; #100;
A = 16'h00A1; B = 16'h0071; #100;
A = 16'h00A1; B = 16'h0072; #100;
A = 16'h00A1; B = 16'h0073; #100;
A = 16'h00A1; B = 16'h0074; #100;
A = 16'h00A1; B = 16'h0075; #100;
A = 16'h00A1; B = 16'h0076; #100;
A = 16'h00A1; B = 16'h0077; #100;
A = 16'h00A1; B = 16'h0078; #100;
A = 16'h00A1; B = 16'h0079; #100;
A = 16'h00A1; B = 16'h007A; #100;
A = 16'h00A1; B = 16'h007B; #100;
A = 16'h00A1; B = 16'h007C; #100;
A = 16'h00A1; B = 16'h007D; #100;
A = 16'h00A1; B = 16'h007E; #100;
A = 16'h00A1; B = 16'h007F; #100;
A = 16'h00A1; B = 16'h0080; #100;
A = 16'h00A1; B = 16'h0081; #100;
A = 16'h00A1; B = 16'h0082; #100;
A = 16'h00A1; B = 16'h0083; #100;
A = 16'h00A1; B = 16'h0084; #100;
A = 16'h00A1; B = 16'h0085; #100;
A = 16'h00A1; B = 16'h0086; #100;
A = 16'h00A1; B = 16'h0087; #100;
A = 16'h00A1; B = 16'h0088; #100;
A = 16'h00A1; B = 16'h0089; #100;
A = 16'h00A1; B = 16'h008A; #100;
A = 16'h00A1; B = 16'h008B; #100;
A = 16'h00A1; B = 16'h008C; #100;
A = 16'h00A1; B = 16'h008D; #100;
A = 16'h00A1; B = 16'h008E; #100;
A = 16'h00A1; B = 16'h008F; #100;
A = 16'h00A1; B = 16'h0090; #100;
A = 16'h00A1; B = 16'h0091; #100;
A = 16'h00A1; B = 16'h0092; #100;
A = 16'h00A1; B = 16'h0093; #100;
A = 16'h00A1; B = 16'h0094; #100;
A = 16'h00A1; B = 16'h0095; #100;
A = 16'h00A1; B = 16'h0096; #100;
A = 16'h00A1; B = 16'h0097; #100;
A = 16'h00A1; B = 16'h0098; #100;
A = 16'h00A1; B = 16'h0099; #100;
A = 16'h00A1; B = 16'h009A; #100;
A = 16'h00A1; B = 16'h009B; #100;
A = 16'h00A1; B = 16'h009C; #100;
A = 16'h00A1; B = 16'h009D; #100;
A = 16'h00A1; B = 16'h009E; #100;
A = 16'h00A1; B = 16'h009F; #100;
A = 16'h00A1; B = 16'h00A0; #100;
A = 16'h00A1; B = 16'h00A1; #100;
A = 16'h00A1; B = 16'h00A2; #100;
A = 16'h00A1; B = 16'h00A3; #100;
A = 16'h00A1; B = 16'h00A4; #100;
A = 16'h00A1; B = 16'h00A5; #100;
A = 16'h00A1; B = 16'h00A6; #100;
A = 16'h00A1; B = 16'h00A7; #100;
A = 16'h00A1; B = 16'h00A8; #100;
A = 16'h00A1; B = 16'h00A9; #100;
A = 16'h00A1; B = 16'h00AA; #100;
A = 16'h00A1; B = 16'h00AB; #100;
A = 16'h00A1; B = 16'h00AC; #100;
A = 16'h00A1; B = 16'h00AD; #100;
A = 16'h00A1; B = 16'h00AE; #100;
A = 16'h00A1; B = 16'h00AF; #100;
A = 16'h00A1; B = 16'h00B0; #100;
A = 16'h00A1; B = 16'h00B1; #100;
A = 16'h00A1; B = 16'h00B2; #100;
A = 16'h00A1; B = 16'h00B3; #100;
A = 16'h00A1; B = 16'h00B4; #100;
A = 16'h00A1; B = 16'h00B5; #100;
A = 16'h00A1; B = 16'h00B6; #100;
A = 16'h00A1; B = 16'h00B7; #100;
A = 16'h00A1; B = 16'h00B8; #100;
A = 16'h00A1; B = 16'h00B9; #100;
A = 16'h00A1; B = 16'h00BA; #100;
A = 16'h00A1; B = 16'h00BB; #100;
A = 16'h00A1; B = 16'h00BC; #100;
A = 16'h00A1; B = 16'h00BD; #100;
A = 16'h00A1; B = 16'h00BE; #100;
A = 16'h00A1; B = 16'h00BF; #100;
A = 16'h00A1; B = 16'h00C0; #100;
A = 16'h00A1; B = 16'h00C1; #100;
A = 16'h00A1; B = 16'h00C2; #100;
A = 16'h00A1; B = 16'h00C3; #100;
A = 16'h00A1; B = 16'h00C4; #100;
A = 16'h00A1; B = 16'h00C5; #100;
A = 16'h00A1; B = 16'h00C6; #100;
A = 16'h00A1; B = 16'h00C7; #100;
A = 16'h00A1; B = 16'h00C8; #100;
A = 16'h00A1; B = 16'h00C9; #100;
A = 16'h00A1; B = 16'h00CA; #100;
A = 16'h00A1; B = 16'h00CB; #100;
A = 16'h00A1; B = 16'h00CC; #100;
A = 16'h00A1; B = 16'h00CD; #100;
A = 16'h00A1; B = 16'h00CE; #100;
A = 16'h00A1; B = 16'h00CF; #100;
A = 16'h00A1; B = 16'h00D0; #100;
A = 16'h00A1; B = 16'h00D1; #100;
A = 16'h00A1; B = 16'h00D2; #100;
A = 16'h00A1; B = 16'h00D3; #100;
A = 16'h00A1; B = 16'h00D4; #100;
A = 16'h00A1; B = 16'h00D5; #100;
A = 16'h00A1; B = 16'h00D6; #100;
A = 16'h00A1; B = 16'h00D7; #100;
A = 16'h00A1; B = 16'h00D8; #100;
A = 16'h00A1; B = 16'h00D9; #100;
A = 16'h00A1; B = 16'h00DA; #100;
A = 16'h00A1; B = 16'h00DB; #100;
A = 16'h00A1; B = 16'h00DC; #100;
A = 16'h00A1; B = 16'h00DD; #100;
A = 16'h00A1; B = 16'h00DE; #100;
A = 16'h00A1; B = 16'h00DF; #100;
A = 16'h00A1; B = 16'h00E0; #100;
A = 16'h00A1; B = 16'h00E1; #100;
A = 16'h00A1; B = 16'h00E2; #100;
A = 16'h00A1; B = 16'h00E3; #100;
A = 16'h00A1; B = 16'h00E4; #100;
A = 16'h00A1; B = 16'h00E5; #100;
A = 16'h00A1; B = 16'h00E6; #100;
A = 16'h00A1; B = 16'h00E7; #100;
A = 16'h00A1; B = 16'h00E8; #100;
A = 16'h00A1; B = 16'h00E9; #100;
A = 16'h00A1; B = 16'h00EA; #100;
A = 16'h00A1; B = 16'h00EB; #100;
A = 16'h00A1; B = 16'h00EC; #100;
A = 16'h00A1; B = 16'h00ED; #100;
A = 16'h00A1; B = 16'h00EE; #100;
A = 16'h00A1; B = 16'h00EF; #100;
A = 16'h00A1; B = 16'h00F0; #100;
A = 16'h00A1; B = 16'h00F1; #100;
A = 16'h00A1; B = 16'h00F2; #100;
A = 16'h00A1; B = 16'h00F3; #100;
A = 16'h00A1; B = 16'h00F4; #100;
A = 16'h00A1; B = 16'h00F5; #100;
A = 16'h00A1; B = 16'h00F6; #100;
A = 16'h00A1; B = 16'h00F7; #100;
A = 16'h00A1; B = 16'h00F8; #100;
A = 16'h00A1; B = 16'h00F9; #100;
A = 16'h00A1; B = 16'h00FA; #100;
A = 16'h00A1; B = 16'h00FB; #100;
A = 16'h00A1; B = 16'h00FC; #100;
A = 16'h00A1; B = 16'h00FD; #100;
A = 16'h00A1; B = 16'h00FE; #100;
A = 16'h00A1; B = 16'h00FF; #100;
A = 16'h00A2; B = 16'h000; #100;
A = 16'h00A2; B = 16'h001; #100;
A = 16'h00A2; B = 16'h002; #100;
A = 16'h00A2; B = 16'h003; #100;
A = 16'h00A2; B = 16'h004; #100;
A = 16'h00A2; B = 16'h005; #100;
A = 16'h00A2; B = 16'h006; #100;
A = 16'h00A2; B = 16'h007; #100;
A = 16'h00A2; B = 16'h008; #100;
A = 16'h00A2; B = 16'h009; #100;
A = 16'h00A2; B = 16'h00A; #100;
A = 16'h00A2; B = 16'h00B; #100;
A = 16'h00A2; B = 16'h00C; #100;
A = 16'h00A2; B = 16'h00D; #100;
A = 16'h00A2; B = 16'h00E; #100;
A = 16'h00A2; B = 16'h00F; #100;
A = 16'h00A2; B = 16'h0010; #100;
A = 16'h00A2; B = 16'h0011; #100;
A = 16'h00A2; B = 16'h0012; #100;
A = 16'h00A2; B = 16'h0013; #100;
A = 16'h00A2; B = 16'h0014; #100;
A = 16'h00A2; B = 16'h0015; #100;
A = 16'h00A2; B = 16'h0016; #100;
A = 16'h00A2; B = 16'h0017; #100;
A = 16'h00A2; B = 16'h0018; #100;
A = 16'h00A2; B = 16'h0019; #100;
A = 16'h00A2; B = 16'h001A; #100;
A = 16'h00A2; B = 16'h001B; #100;
A = 16'h00A2; B = 16'h001C; #100;
A = 16'h00A2; B = 16'h001D; #100;
A = 16'h00A2; B = 16'h001E; #100;
A = 16'h00A2; B = 16'h001F; #100;
A = 16'h00A2; B = 16'h0020; #100;
A = 16'h00A2; B = 16'h0021; #100;
A = 16'h00A2; B = 16'h0022; #100;
A = 16'h00A2; B = 16'h0023; #100;
A = 16'h00A2; B = 16'h0024; #100;
A = 16'h00A2; B = 16'h0025; #100;
A = 16'h00A2; B = 16'h0026; #100;
A = 16'h00A2; B = 16'h0027; #100;
A = 16'h00A2; B = 16'h0028; #100;
A = 16'h00A2; B = 16'h0029; #100;
A = 16'h00A2; B = 16'h002A; #100;
A = 16'h00A2; B = 16'h002B; #100;
A = 16'h00A2; B = 16'h002C; #100;
A = 16'h00A2; B = 16'h002D; #100;
A = 16'h00A2; B = 16'h002E; #100;
A = 16'h00A2; B = 16'h002F; #100;
A = 16'h00A2; B = 16'h0030; #100;
A = 16'h00A2; B = 16'h0031; #100;
A = 16'h00A2; B = 16'h0032; #100;
A = 16'h00A2; B = 16'h0033; #100;
A = 16'h00A2; B = 16'h0034; #100;
A = 16'h00A2; B = 16'h0035; #100;
A = 16'h00A2; B = 16'h0036; #100;
A = 16'h00A2; B = 16'h0037; #100;
A = 16'h00A2; B = 16'h0038; #100;
A = 16'h00A2; B = 16'h0039; #100;
A = 16'h00A2; B = 16'h003A; #100;
A = 16'h00A2; B = 16'h003B; #100;
A = 16'h00A2; B = 16'h003C; #100;
A = 16'h00A2; B = 16'h003D; #100;
A = 16'h00A2; B = 16'h003E; #100;
A = 16'h00A2; B = 16'h003F; #100;
A = 16'h00A2; B = 16'h0040; #100;
A = 16'h00A2; B = 16'h0041; #100;
A = 16'h00A2; B = 16'h0042; #100;
A = 16'h00A2; B = 16'h0043; #100;
A = 16'h00A2; B = 16'h0044; #100;
A = 16'h00A2; B = 16'h0045; #100;
A = 16'h00A2; B = 16'h0046; #100;
A = 16'h00A2; B = 16'h0047; #100;
A = 16'h00A2; B = 16'h0048; #100;
A = 16'h00A2; B = 16'h0049; #100;
A = 16'h00A2; B = 16'h004A; #100;
A = 16'h00A2; B = 16'h004B; #100;
A = 16'h00A2; B = 16'h004C; #100;
A = 16'h00A2; B = 16'h004D; #100;
A = 16'h00A2; B = 16'h004E; #100;
A = 16'h00A2; B = 16'h004F; #100;
A = 16'h00A2; B = 16'h0050; #100;
A = 16'h00A2; B = 16'h0051; #100;
A = 16'h00A2; B = 16'h0052; #100;
A = 16'h00A2; B = 16'h0053; #100;
A = 16'h00A2; B = 16'h0054; #100;
A = 16'h00A2; B = 16'h0055; #100;
A = 16'h00A2; B = 16'h0056; #100;
A = 16'h00A2; B = 16'h0057; #100;
A = 16'h00A2; B = 16'h0058; #100;
A = 16'h00A2; B = 16'h0059; #100;
A = 16'h00A2; B = 16'h005A; #100;
A = 16'h00A2; B = 16'h005B; #100;
A = 16'h00A2; B = 16'h005C; #100;
A = 16'h00A2; B = 16'h005D; #100;
A = 16'h00A2; B = 16'h005E; #100;
A = 16'h00A2; B = 16'h005F; #100;
A = 16'h00A2; B = 16'h0060; #100;
A = 16'h00A2; B = 16'h0061; #100;
A = 16'h00A2; B = 16'h0062; #100;
A = 16'h00A2; B = 16'h0063; #100;
A = 16'h00A2; B = 16'h0064; #100;
A = 16'h00A2; B = 16'h0065; #100;
A = 16'h00A2; B = 16'h0066; #100;
A = 16'h00A2; B = 16'h0067; #100;
A = 16'h00A2; B = 16'h0068; #100;
A = 16'h00A2; B = 16'h0069; #100;
A = 16'h00A2; B = 16'h006A; #100;
A = 16'h00A2; B = 16'h006B; #100;
A = 16'h00A2; B = 16'h006C; #100;
A = 16'h00A2; B = 16'h006D; #100;
A = 16'h00A2; B = 16'h006E; #100;
A = 16'h00A2; B = 16'h006F; #100;
A = 16'h00A2; B = 16'h0070; #100;
A = 16'h00A2; B = 16'h0071; #100;
A = 16'h00A2; B = 16'h0072; #100;
A = 16'h00A2; B = 16'h0073; #100;
A = 16'h00A2; B = 16'h0074; #100;
A = 16'h00A2; B = 16'h0075; #100;
A = 16'h00A2; B = 16'h0076; #100;
A = 16'h00A2; B = 16'h0077; #100;
A = 16'h00A2; B = 16'h0078; #100;
A = 16'h00A2; B = 16'h0079; #100;
A = 16'h00A2; B = 16'h007A; #100;
A = 16'h00A2; B = 16'h007B; #100;
A = 16'h00A2; B = 16'h007C; #100;
A = 16'h00A2; B = 16'h007D; #100;
A = 16'h00A2; B = 16'h007E; #100;
A = 16'h00A2; B = 16'h007F; #100;
A = 16'h00A2; B = 16'h0080; #100;
A = 16'h00A2; B = 16'h0081; #100;
A = 16'h00A2; B = 16'h0082; #100;
A = 16'h00A2; B = 16'h0083; #100;
A = 16'h00A2; B = 16'h0084; #100;
A = 16'h00A2; B = 16'h0085; #100;
A = 16'h00A2; B = 16'h0086; #100;
A = 16'h00A2; B = 16'h0087; #100;
A = 16'h00A2; B = 16'h0088; #100;
A = 16'h00A2; B = 16'h0089; #100;
A = 16'h00A2; B = 16'h008A; #100;
A = 16'h00A2; B = 16'h008B; #100;
A = 16'h00A2; B = 16'h008C; #100;
A = 16'h00A2; B = 16'h008D; #100;
A = 16'h00A2; B = 16'h008E; #100;
A = 16'h00A2; B = 16'h008F; #100;
A = 16'h00A2; B = 16'h0090; #100;
A = 16'h00A2; B = 16'h0091; #100;
A = 16'h00A2; B = 16'h0092; #100;
A = 16'h00A2; B = 16'h0093; #100;
A = 16'h00A2; B = 16'h0094; #100;
A = 16'h00A2; B = 16'h0095; #100;
A = 16'h00A2; B = 16'h0096; #100;
A = 16'h00A2; B = 16'h0097; #100;
A = 16'h00A2; B = 16'h0098; #100;
A = 16'h00A2; B = 16'h0099; #100;
A = 16'h00A2; B = 16'h009A; #100;
A = 16'h00A2; B = 16'h009B; #100;
A = 16'h00A2; B = 16'h009C; #100;
A = 16'h00A2; B = 16'h009D; #100;
A = 16'h00A2; B = 16'h009E; #100;
A = 16'h00A2; B = 16'h009F; #100;
A = 16'h00A2; B = 16'h00A0; #100;
A = 16'h00A2; B = 16'h00A1; #100;
A = 16'h00A2; B = 16'h00A2; #100;
A = 16'h00A2; B = 16'h00A3; #100;
A = 16'h00A2; B = 16'h00A4; #100;
A = 16'h00A2; B = 16'h00A5; #100;
A = 16'h00A2; B = 16'h00A6; #100;
A = 16'h00A2; B = 16'h00A7; #100;
A = 16'h00A2; B = 16'h00A8; #100;
A = 16'h00A2; B = 16'h00A9; #100;
A = 16'h00A2; B = 16'h00AA; #100;
A = 16'h00A2; B = 16'h00AB; #100;
A = 16'h00A2; B = 16'h00AC; #100;
A = 16'h00A2; B = 16'h00AD; #100;
A = 16'h00A2; B = 16'h00AE; #100;
A = 16'h00A2; B = 16'h00AF; #100;
A = 16'h00A2; B = 16'h00B0; #100;
A = 16'h00A2; B = 16'h00B1; #100;
A = 16'h00A2; B = 16'h00B2; #100;
A = 16'h00A2; B = 16'h00B3; #100;
A = 16'h00A2; B = 16'h00B4; #100;
A = 16'h00A2; B = 16'h00B5; #100;
A = 16'h00A2; B = 16'h00B6; #100;
A = 16'h00A2; B = 16'h00B7; #100;
A = 16'h00A2; B = 16'h00B8; #100;
A = 16'h00A2; B = 16'h00B9; #100;
A = 16'h00A2; B = 16'h00BA; #100;
A = 16'h00A2; B = 16'h00BB; #100;
A = 16'h00A2; B = 16'h00BC; #100;
A = 16'h00A2; B = 16'h00BD; #100;
A = 16'h00A2; B = 16'h00BE; #100;
A = 16'h00A2; B = 16'h00BF; #100;
A = 16'h00A2; B = 16'h00C0; #100;
A = 16'h00A2; B = 16'h00C1; #100;
A = 16'h00A2; B = 16'h00C2; #100;
A = 16'h00A2; B = 16'h00C3; #100;
A = 16'h00A2; B = 16'h00C4; #100;
A = 16'h00A2; B = 16'h00C5; #100;
A = 16'h00A2; B = 16'h00C6; #100;
A = 16'h00A2; B = 16'h00C7; #100;
A = 16'h00A2; B = 16'h00C8; #100;
A = 16'h00A2; B = 16'h00C9; #100;
A = 16'h00A2; B = 16'h00CA; #100;
A = 16'h00A2; B = 16'h00CB; #100;
A = 16'h00A2; B = 16'h00CC; #100;
A = 16'h00A2; B = 16'h00CD; #100;
A = 16'h00A2; B = 16'h00CE; #100;
A = 16'h00A2; B = 16'h00CF; #100;
A = 16'h00A2; B = 16'h00D0; #100;
A = 16'h00A2; B = 16'h00D1; #100;
A = 16'h00A2; B = 16'h00D2; #100;
A = 16'h00A2; B = 16'h00D3; #100;
A = 16'h00A2; B = 16'h00D4; #100;
A = 16'h00A2; B = 16'h00D5; #100;
A = 16'h00A2; B = 16'h00D6; #100;
A = 16'h00A2; B = 16'h00D7; #100;
A = 16'h00A2; B = 16'h00D8; #100;
A = 16'h00A2; B = 16'h00D9; #100;
A = 16'h00A2; B = 16'h00DA; #100;
A = 16'h00A2; B = 16'h00DB; #100;
A = 16'h00A2; B = 16'h00DC; #100;
A = 16'h00A2; B = 16'h00DD; #100;
A = 16'h00A2; B = 16'h00DE; #100;
A = 16'h00A2; B = 16'h00DF; #100;
A = 16'h00A2; B = 16'h00E0; #100;
A = 16'h00A2; B = 16'h00E1; #100;
A = 16'h00A2; B = 16'h00E2; #100;
A = 16'h00A2; B = 16'h00E3; #100;
A = 16'h00A2; B = 16'h00E4; #100;
A = 16'h00A2; B = 16'h00E5; #100;
A = 16'h00A2; B = 16'h00E6; #100;
A = 16'h00A2; B = 16'h00E7; #100;
A = 16'h00A2; B = 16'h00E8; #100;
A = 16'h00A2; B = 16'h00E9; #100;
A = 16'h00A2; B = 16'h00EA; #100;
A = 16'h00A2; B = 16'h00EB; #100;
A = 16'h00A2; B = 16'h00EC; #100;
A = 16'h00A2; B = 16'h00ED; #100;
A = 16'h00A2; B = 16'h00EE; #100;
A = 16'h00A2; B = 16'h00EF; #100;
A = 16'h00A2; B = 16'h00F0; #100;
A = 16'h00A2; B = 16'h00F1; #100;
A = 16'h00A2; B = 16'h00F2; #100;
A = 16'h00A2; B = 16'h00F3; #100;
A = 16'h00A2; B = 16'h00F4; #100;
A = 16'h00A2; B = 16'h00F5; #100;
A = 16'h00A2; B = 16'h00F6; #100;
A = 16'h00A2; B = 16'h00F7; #100;
A = 16'h00A2; B = 16'h00F8; #100;
A = 16'h00A2; B = 16'h00F9; #100;
A = 16'h00A2; B = 16'h00FA; #100;
A = 16'h00A2; B = 16'h00FB; #100;
A = 16'h00A2; B = 16'h00FC; #100;
A = 16'h00A2; B = 16'h00FD; #100;
A = 16'h00A2; B = 16'h00FE; #100;
A = 16'h00A2; B = 16'h00FF; #100;
A = 16'h00A3; B = 16'h000; #100;
A = 16'h00A3; B = 16'h001; #100;
A = 16'h00A3; B = 16'h002; #100;
A = 16'h00A3; B = 16'h003; #100;
A = 16'h00A3; B = 16'h004; #100;
A = 16'h00A3; B = 16'h005; #100;
A = 16'h00A3; B = 16'h006; #100;
A = 16'h00A3; B = 16'h007; #100;
A = 16'h00A3; B = 16'h008; #100;
A = 16'h00A3; B = 16'h009; #100;
A = 16'h00A3; B = 16'h00A; #100;
A = 16'h00A3; B = 16'h00B; #100;
A = 16'h00A3; B = 16'h00C; #100;
A = 16'h00A3; B = 16'h00D; #100;
A = 16'h00A3; B = 16'h00E; #100;
A = 16'h00A3; B = 16'h00F; #100;
A = 16'h00A3; B = 16'h0010; #100;
A = 16'h00A3; B = 16'h0011; #100;
A = 16'h00A3; B = 16'h0012; #100;
A = 16'h00A3; B = 16'h0013; #100;
A = 16'h00A3; B = 16'h0014; #100;
A = 16'h00A3; B = 16'h0015; #100;
A = 16'h00A3; B = 16'h0016; #100;
A = 16'h00A3; B = 16'h0017; #100;
A = 16'h00A3; B = 16'h0018; #100;
A = 16'h00A3; B = 16'h0019; #100;
A = 16'h00A3; B = 16'h001A; #100;
A = 16'h00A3; B = 16'h001B; #100;
A = 16'h00A3; B = 16'h001C; #100;
A = 16'h00A3; B = 16'h001D; #100;
A = 16'h00A3; B = 16'h001E; #100;
A = 16'h00A3; B = 16'h001F; #100;
A = 16'h00A3; B = 16'h0020; #100;
A = 16'h00A3; B = 16'h0021; #100;
A = 16'h00A3; B = 16'h0022; #100;
A = 16'h00A3; B = 16'h0023; #100;
A = 16'h00A3; B = 16'h0024; #100;
A = 16'h00A3; B = 16'h0025; #100;
A = 16'h00A3; B = 16'h0026; #100;
A = 16'h00A3; B = 16'h0027; #100;
A = 16'h00A3; B = 16'h0028; #100;
A = 16'h00A3; B = 16'h0029; #100;
A = 16'h00A3; B = 16'h002A; #100;
A = 16'h00A3; B = 16'h002B; #100;
A = 16'h00A3; B = 16'h002C; #100;
A = 16'h00A3; B = 16'h002D; #100;
A = 16'h00A3; B = 16'h002E; #100;
A = 16'h00A3; B = 16'h002F; #100;
A = 16'h00A3; B = 16'h0030; #100;
A = 16'h00A3; B = 16'h0031; #100;
A = 16'h00A3; B = 16'h0032; #100;
A = 16'h00A3; B = 16'h0033; #100;
A = 16'h00A3; B = 16'h0034; #100;
A = 16'h00A3; B = 16'h0035; #100;
A = 16'h00A3; B = 16'h0036; #100;
A = 16'h00A3; B = 16'h0037; #100;
A = 16'h00A3; B = 16'h0038; #100;
A = 16'h00A3; B = 16'h0039; #100;
A = 16'h00A3; B = 16'h003A; #100;
A = 16'h00A3; B = 16'h003B; #100;
A = 16'h00A3; B = 16'h003C; #100;
A = 16'h00A3; B = 16'h003D; #100;
A = 16'h00A3; B = 16'h003E; #100;
A = 16'h00A3; B = 16'h003F; #100;
A = 16'h00A3; B = 16'h0040; #100;
A = 16'h00A3; B = 16'h0041; #100;
A = 16'h00A3; B = 16'h0042; #100;
A = 16'h00A3; B = 16'h0043; #100;
A = 16'h00A3; B = 16'h0044; #100;
A = 16'h00A3; B = 16'h0045; #100;
A = 16'h00A3; B = 16'h0046; #100;
A = 16'h00A3; B = 16'h0047; #100;
A = 16'h00A3; B = 16'h0048; #100;
A = 16'h00A3; B = 16'h0049; #100;
A = 16'h00A3; B = 16'h004A; #100;
A = 16'h00A3; B = 16'h004B; #100;
A = 16'h00A3; B = 16'h004C; #100;
A = 16'h00A3; B = 16'h004D; #100;
A = 16'h00A3; B = 16'h004E; #100;
A = 16'h00A3; B = 16'h004F; #100;
A = 16'h00A3; B = 16'h0050; #100;
A = 16'h00A3; B = 16'h0051; #100;
A = 16'h00A3; B = 16'h0052; #100;
A = 16'h00A3; B = 16'h0053; #100;
A = 16'h00A3; B = 16'h0054; #100;
A = 16'h00A3; B = 16'h0055; #100;
A = 16'h00A3; B = 16'h0056; #100;
A = 16'h00A3; B = 16'h0057; #100;
A = 16'h00A3; B = 16'h0058; #100;
A = 16'h00A3; B = 16'h0059; #100;
A = 16'h00A3; B = 16'h005A; #100;
A = 16'h00A3; B = 16'h005B; #100;
A = 16'h00A3; B = 16'h005C; #100;
A = 16'h00A3; B = 16'h005D; #100;
A = 16'h00A3; B = 16'h005E; #100;
A = 16'h00A3; B = 16'h005F; #100;
A = 16'h00A3; B = 16'h0060; #100;
A = 16'h00A3; B = 16'h0061; #100;
A = 16'h00A3; B = 16'h0062; #100;
A = 16'h00A3; B = 16'h0063; #100;
A = 16'h00A3; B = 16'h0064; #100;
A = 16'h00A3; B = 16'h0065; #100;
A = 16'h00A3; B = 16'h0066; #100;
A = 16'h00A3; B = 16'h0067; #100;
A = 16'h00A3; B = 16'h0068; #100;
A = 16'h00A3; B = 16'h0069; #100;
A = 16'h00A3; B = 16'h006A; #100;
A = 16'h00A3; B = 16'h006B; #100;
A = 16'h00A3; B = 16'h006C; #100;
A = 16'h00A3; B = 16'h006D; #100;
A = 16'h00A3; B = 16'h006E; #100;
A = 16'h00A3; B = 16'h006F; #100;
A = 16'h00A3; B = 16'h0070; #100;
A = 16'h00A3; B = 16'h0071; #100;
A = 16'h00A3; B = 16'h0072; #100;
A = 16'h00A3; B = 16'h0073; #100;
A = 16'h00A3; B = 16'h0074; #100;
A = 16'h00A3; B = 16'h0075; #100;
A = 16'h00A3; B = 16'h0076; #100;
A = 16'h00A3; B = 16'h0077; #100;
A = 16'h00A3; B = 16'h0078; #100;
A = 16'h00A3; B = 16'h0079; #100;
A = 16'h00A3; B = 16'h007A; #100;
A = 16'h00A3; B = 16'h007B; #100;
A = 16'h00A3; B = 16'h007C; #100;
A = 16'h00A3; B = 16'h007D; #100;
A = 16'h00A3; B = 16'h007E; #100;
A = 16'h00A3; B = 16'h007F; #100;
A = 16'h00A3; B = 16'h0080; #100;
A = 16'h00A3; B = 16'h0081; #100;
A = 16'h00A3; B = 16'h0082; #100;
A = 16'h00A3; B = 16'h0083; #100;
A = 16'h00A3; B = 16'h0084; #100;
A = 16'h00A3; B = 16'h0085; #100;
A = 16'h00A3; B = 16'h0086; #100;
A = 16'h00A3; B = 16'h0087; #100;
A = 16'h00A3; B = 16'h0088; #100;
A = 16'h00A3; B = 16'h0089; #100;
A = 16'h00A3; B = 16'h008A; #100;
A = 16'h00A3; B = 16'h008B; #100;
A = 16'h00A3; B = 16'h008C; #100;
A = 16'h00A3; B = 16'h008D; #100;
A = 16'h00A3; B = 16'h008E; #100;
A = 16'h00A3; B = 16'h008F; #100;
A = 16'h00A3; B = 16'h0090; #100;
A = 16'h00A3; B = 16'h0091; #100;
A = 16'h00A3; B = 16'h0092; #100;
A = 16'h00A3; B = 16'h0093; #100;
A = 16'h00A3; B = 16'h0094; #100;
A = 16'h00A3; B = 16'h0095; #100;
A = 16'h00A3; B = 16'h0096; #100;
A = 16'h00A3; B = 16'h0097; #100;
A = 16'h00A3; B = 16'h0098; #100;
A = 16'h00A3; B = 16'h0099; #100;
A = 16'h00A3; B = 16'h009A; #100;
A = 16'h00A3; B = 16'h009B; #100;
A = 16'h00A3; B = 16'h009C; #100;
A = 16'h00A3; B = 16'h009D; #100;
A = 16'h00A3; B = 16'h009E; #100;
A = 16'h00A3; B = 16'h009F; #100;
A = 16'h00A3; B = 16'h00A0; #100;
A = 16'h00A3; B = 16'h00A1; #100;
A = 16'h00A3; B = 16'h00A2; #100;
A = 16'h00A3; B = 16'h00A3; #100;
A = 16'h00A3; B = 16'h00A4; #100;
A = 16'h00A3; B = 16'h00A5; #100;
A = 16'h00A3; B = 16'h00A6; #100;
A = 16'h00A3; B = 16'h00A7; #100;
A = 16'h00A3; B = 16'h00A8; #100;
A = 16'h00A3; B = 16'h00A9; #100;
A = 16'h00A3; B = 16'h00AA; #100;
A = 16'h00A3; B = 16'h00AB; #100;
A = 16'h00A3; B = 16'h00AC; #100;
A = 16'h00A3; B = 16'h00AD; #100;
A = 16'h00A3; B = 16'h00AE; #100;
A = 16'h00A3; B = 16'h00AF; #100;
A = 16'h00A3; B = 16'h00B0; #100;
A = 16'h00A3; B = 16'h00B1; #100;
A = 16'h00A3; B = 16'h00B2; #100;
A = 16'h00A3; B = 16'h00B3; #100;
A = 16'h00A3; B = 16'h00B4; #100;
A = 16'h00A3; B = 16'h00B5; #100;
A = 16'h00A3; B = 16'h00B6; #100;
A = 16'h00A3; B = 16'h00B7; #100;
A = 16'h00A3; B = 16'h00B8; #100;
A = 16'h00A3; B = 16'h00B9; #100;
A = 16'h00A3; B = 16'h00BA; #100;
A = 16'h00A3; B = 16'h00BB; #100;
A = 16'h00A3; B = 16'h00BC; #100;
A = 16'h00A3; B = 16'h00BD; #100;
A = 16'h00A3; B = 16'h00BE; #100;
A = 16'h00A3; B = 16'h00BF; #100;
A = 16'h00A3; B = 16'h00C0; #100;
A = 16'h00A3; B = 16'h00C1; #100;
A = 16'h00A3; B = 16'h00C2; #100;
A = 16'h00A3; B = 16'h00C3; #100;
A = 16'h00A3; B = 16'h00C4; #100;
A = 16'h00A3; B = 16'h00C5; #100;
A = 16'h00A3; B = 16'h00C6; #100;
A = 16'h00A3; B = 16'h00C7; #100;
A = 16'h00A3; B = 16'h00C8; #100;
A = 16'h00A3; B = 16'h00C9; #100;
A = 16'h00A3; B = 16'h00CA; #100;
A = 16'h00A3; B = 16'h00CB; #100;
A = 16'h00A3; B = 16'h00CC; #100;
A = 16'h00A3; B = 16'h00CD; #100;
A = 16'h00A3; B = 16'h00CE; #100;
A = 16'h00A3; B = 16'h00CF; #100;
A = 16'h00A3; B = 16'h00D0; #100;
A = 16'h00A3; B = 16'h00D1; #100;
A = 16'h00A3; B = 16'h00D2; #100;
A = 16'h00A3; B = 16'h00D3; #100;
A = 16'h00A3; B = 16'h00D4; #100;
A = 16'h00A3; B = 16'h00D5; #100;
A = 16'h00A3; B = 16'h00D6; #100;
A = 16'h00A3; B = 16'h00D7; #100;
A = 16'h00A3; B = 16'h00D8; #100;
A = 16'h00A3; B = 16'h00D9; #100;
A = 16'h00A3; B = 16'h00DA; #100;
A = 16'h00A3; B = 16'h00DB; #100;
A = 16'h00A3; B = 16'h00DC; #100;
A = 16'h00A3; B = 16'h00DD; #100;
A = 16'h00A3; B = 16'h00DE; #100;
A = 16'h00A3; B = 16'h00DF; #100;
A = 16'h00A3; B = 16'h00E0; #100;
A = 16'h00A3; B = 16'h00E1; #100;
A = 16'h00A3; B = 16'h00E2; #100;
A = 16'h00A3; B = 16'h00E3; #100;
A = 16'h00A3; B = 16'h00E4; #100;
A = 16'h00A3; B = 16'h00E5; #100;
A = 16'h00A3; B = 16'h00E6; #100;
A = 16'h00A3; B = 16'h00E7; #100;
A = 16'h00A3; B = 16'h00E8; #100;
A = 16'h00A3; B = 16'h00E9; #100;
A = 16'h00A3; B = 16'h00EA; #100;
A = 16'h00A3; B = 16'h00EB; #100;
A = 16'h00A3; B = 16'h00EC; #100;
A = 16'h00A3; B = 16'h00ED; #100;
A = 16'h00A3; B = 16'h00EE; #100;
A = 16'h00A3; B = 16'h00EF; #100;
A = 16'h00A3; B = 16'h00F0; #100;
A = 16'h00A3; B = 16'h00F1; #100;
A = 16'h00A3; B = 16'h00F2; #100;
A = 16'h00A3; B = 16'h00F3; #100;
A = 16'h00A3; B = 16'h00F4; #100;
A = 16'h00A3; B = 16'h00F5; #100;
A = 16'h00A3; B = 16'h00F6; #100;
A = 16'h00A3; B = 16'h00F7; #100;
A = 16'h00A3; B = 16'h00F8; #100;
A = 16'h00A3; B = 16'h00F9; #100;
A = 16'h00A3; B = 16'h00FA; #100;
A = 16'h00A3; B = 16'h00FB; #100;
A = 16'h00A3; B = 16'h00FC; #100;
A = 16'h00A3; B = 16'h00FD; #100;
A = 16'h00A3; B = 16'h00FE; #100;
A = 16'h00A3; B = 16'h00FF; #100;
A = 16'h00A4; B = 16'h000; #100;
A = 16'h00A4; B = 16'h001; #100;
A = 16'h00A4; B = 16'h002; #100;
A = 16'h00A4; B = 16'h003; #100;
A = 16'h00A4; B = 16'h004; #100;
A = 16'h00A4; B = 16'h005; #100;
A = 16'h00A4; B = 16'h006; #100;
A = 16'h00A4; B = 16'h007; #100;
A = 16'h00A4; B = 16'h008; #100;
A = 16'h00A4; B = 16'h009; #100;
A = 16'h00A4; B = 16'h00A; #100;
A = 16'h00A4; B = 16'h00B; #100;
A = 16'h00A4; B = 16'h00C; #100;
A = 16'h00A4; B = 16'h00D; #100;
A = 16'h00A4; B = 16'h00E; #100;
A = 16'h00A4; B = 16'h00F; #100;
A = 16'h00A4; B = 16'h0010; #100;
A = 16'h00A4; B = 16'h0011; #100;
A = 16'h00A4; B = 16'h0012; #100;
A = 16'h00A4; B = 16'h0013; #100;
A = 16'h00A4; B = 16'h0014; #100;
A = 16'h00A4; B = 16'h0015; #100;
A = 16'h00A4; B = 16'h0016; #100;
A = 16'h00A4; B = 16'h0017; #100;
A = 16'h00A4; B = 16'h0018; #100;
A = 16'h00A4; B = 16'h0019; #100;
A = 16'h00A4; B = 16'h001A; #100;
A = 16'h00A4; B = 16'h001B; #100;
A = 16'h00A4; B = 16'h001C; #100;
A = 16'h00A4; B = 16'h001D; #100;
A = 16'h00A4; B = 16'h001E; #100;
A = 16'h00A4; B = 16'h001F; #100;
A = 16'h00A4; B = 16'h0020; #100;
A = 16'h00A4; B = 16'h0021; #100;
A = 16'h00A4; B = 16'h0022; #100;
A = 16'h00A4; B = 16'h0023; #100;
A = 16'h00A4; B = 16'h0024; #100;
A = 16'h00A4; B = 16'h0025; #100;
A = 16'h00A4; B = 16'h0026; #100;
A = 16'h00A4; B = 16'h0027; #100;
A = 16'h00A4; B = 16'h0028; #100;
A = 16'h00A4; B = 16'h0029; #100;
A = 16'h00A4; B = 16'h002A; #100;
A = 16'h00A4; B = 16'h002B; #100;
A = 16'h00A4; B = 16'h002C; #100;
A = 16'h00A4; B = 16'h002D; #100;
A = 16'h00A4; B = 16'h002E; #100;
A = 16'h00A4; B = 16'h002F; #100;
A = 16'h00A4; B = 16'h0030; #100;
A = 16'h00A4; B = 16'h0031; #100;
A = 16'h00A4; B = 16'h0032; #100;
A = 16'h00A4; B = 16'h0033; #100;
A = 16'h00A4; B = 16'h0034; #100;
A = 16'h00A4; B = 16'h0035; #100;
A = 16'h00A4; B = 16'h0036; #100;
A = 16'h00A4; B = 16'h0037; #100;
A = 16'h00A4; B = 16'h0038; #100;
A = 16'h00A4; B = 16'h0039; #100;
A = 16'h00A4; B = 16'h003A; #100;
A = 16'h00A4; B = 16'h003B; #100;
A = 16'h00A4; B = 16'h003C; #100;
A = 16'h00A4; B = 16'h003D; #100;
A = 16'h00A4; B = 16'h003E; #100;
A = 16'h00A4; B = 16'h003F; #100;
A = 16'h00A4; B = 16'h0040; #100;
A = 16'h00A4; B = 16'h0041; #100;
A = 16'h00A4; B = 16'h0042; #100;
A = 16'h00A4; B = 16'h0043; #100;
A = 16'h00A4; B = 16'h0044; #100;
A = 16'h00A4; B = 16'h0045; #100;
A = 16'h00A4; B = 16'h0046; #100;
A = 16'h00A4; B = 16'h0047; #100;
A = 16'h00A4; B = 16'h0048; #100;
A = 16'h00A4; B = 16'h0049; #100;
A = 16'h00A4; B = 16'h004A; #100;
A = 16'h00A4; B = 16'h004B; #100;
A = 16'h00A4; B = 16'h004C; #100;
A = 16'h00A4; B = 16'h004D; #100;
A = 16'h00A4; B = 16'h004E; #100;
A = 16'h00A4; B = 16'h004F; #100;
A = 16'h00A4; B = 16'h0050; #100;
A = 16'h00A4; B = 16'h0051; #100;
A = 16'h00A4; B = 16'h0052; #100;
A = 16'h00A4; B = 16'h0053; #100;
A = 16'h00A4; B = 16'h0054; #100;
A = 16'h00A4; B = 16'h0055; #100;
A = 16'h00A4; B = 16'h0056; #100;
A = 16'h00A4; B = 16'h0057; #100;
A = 16'h00A4; B = 16'h0058; #100;
A = 16'h00A4; B = 16'h0059; #100;
A = 16'h00A4; B = 16'h005A; #100;
A = 16'h00A4; B = 16'h005B; #100;
A = 16'h00A4; B = 16'h005C; #100;
A = 16'h00A4; B = 16'h005D; #100;
A = 16'h00A4; B = 16'h005E; #100;
A = 16'h00A4; B = 16'h005F; #100;
A = 16'h00A4; B = 16'h0060; #100;
A = 16'h00A4; B = 16'h0061; #100;
A = 16'h00A4; B = 16'h0062; #100;
A = 16'h00A4; B = 16'h0063; #100;
A = 16'h00A4; B = 16'h0064; #100;
A = 16'h00A4; B = 16'h0065; #100;
A = 16'h00A4; B = 16'h0066; #100;
A = 16'h00A4; B = 16'h0067; #100;
A = 16'h00A4; B = 16'h0068; #100;
A = 16'h00A4; B = 16'h0069; #100;
A = 16'h00A4; B = 16'h006A; #100;
A = 16'h00A4; B = 16'h006B; #100;
A = 16'h00A4; B = 16'h006C; #100;
A = 16'h00A4; B = 16'h006D; #100;
A = 16'h00A4; B = 16'h006E; #100;
A = 16'h00A4; B = 16'h006F; #100;
A = 16'h00A4; B = 16'h0070; #100;
A = 16'h00A4; B = 16'h0071; #100;
A = 16'h00A4; B = 16'h0072; #100;
A = 16'h00A4; B = 16'h0073; #100;
A = 16'h00A4; B = 16'h0074; #100;
A = 16'h00A4; B = 16'h0075; #100;
A = 16'h00A4; B = 16'h0076; #100;
A = 16'h00A4; B = 16'h0077; #100;
A = 16'h00A4; B = 16'h0078; #100;
A = 16'h00A4; B = 16'h0079; #100;
A = 16'h00A4; B = 16'h007A; #100;
A = 16'h00A4; B = 16'h007B; #100;
A = 16'h00A4; B = 16'h007C; #100;
A = 16'h00A4; B = 16'h007D; #100;
A = 16'h00A4; B = 16'h007E; #100;
A = 16'h00A4; B = 16'h007F; #100;
A = 16'h00A4; B = 16'h0080; #100;
A = 16'h00A4; B = 16'h0081; #100;
A = 16'h00A4; B = 16'h0082; #100;
A = 16'h00A4; B = 16'h0083; #100;
A = 16'h00A4; B = 16'h0084; #100;
A = 16'h00A4; B = 16'h0085; #100;
A = 16'h00A4; B = 16'h0086; #100;
A = 16'h00A4; B = 16'h0087; #100;
A = 16'h00A4; B = 16'h0088; #100;
A = 16'h00A4; B = 16'h0089; #100;
A = 16'h00A4; B = 16'h008A; #100;
A = 16'h00A4; B = 16'h008B; #100;
A = 16'h00A4; B = 16'h008C; #100;
A = 16'h00A4; B = 16'h008D; #100;
A = 16'h00A4; B = 16'h008E; #100;
A = 16'h00A4; B = 16'h008F; #100;
A = 16'h00A4; B = 16'h0090; #100;
A = 16'h00A4; B = 16'h0091; #100;
A = 16'h00A4; B = 16'h0092; #100;
A = 16'h00A4; B = 16'h0093; #100;
A = 16'h00A4; B = 16'h0094; #100;
A = 16'h00A4; B = 16'h0095; #100;
A = 16'h00A4; B = 16'h0096; #100;
A = 16'h00A4; B = 16'h0097; #100;
A = 16'h00A4; B = 16'h0098; #100;
A = 16'h00A4; B = 16'h0099; #100;
A = 16'h00A4; B = 16'h009A; #100;
A = 16'h00A4; B = 16'h009B; #100;
A = 16'h00A4; B = 16'h009C; #100;
A = 16'h00A4; B = 16'h009D; #100;
A = 16'h00A4; B = 16'h009E; #100;
A = 16'h00A4; B = 16'h009F; #100;
A = 16'h00A4; B = 16'h00A0; #100;
A = 16'h00A4; B = 16'h00A1; #100;
A = 16'h00A4; B = 16'h00A2; #100;
A = 16'h00A4; B = 16'h00A3; #100;
A = 16'h00A4; B = 16'h00A4; #100;
A = 16'h00A4; B = 16'h00A5; #100;
A = 16'h00A4; B = 16'h00A6; #100;
A = 16'h00A4; B = 16'h00A7; #100;
A = 16'h00A4; B = 16'h00A8; #100;
A = 16'h00A4; B = 16'h00A9; #100;
A = 16'h00A4; B = 16'h00AA; #100;
A = 16'h00A4; B = 16'h00AB; #100;
A = 16'h00A4; B = 16'h00AC; #100;
A = 16'h00A4; B = 16'h00AD; #100;
A = 16'h00A4; B = 16'h00AE; #100;
A = 16'h00A4; B = 16'h00AF; #100;
A = 16'h00A4; B = 16'h00B0; #100;
A = 16'h00A4; B = 16'h00B1; #100;
A = 16'h00A4; B = 16'h00B2; #100;
A = 16'h00A4; B = 16'h00B3; #100;
A = 16'h00A4; B = 16'h00B4; #100;
A = 16'h00A4; B = 16'h00B5; #100;
A = 16'h00A4; B = 16'h00B6; #100;
A = 16'h00A4; B = 16'h00B7; #100;
A = 16'h00A4; B = 16'h00B8; #100;
A = 16'h00A4; B = 16'h00B9; #100;
A = 16'h00A4; B = 16'h00BA; #100;
A = 16'h00A4; B = 16'h00BB; #100;
A = 16'h00A4; B = 16'h00BC; #100;
A = 16'h00A4; B = 16'h00BD; #100;
A = 16'h00A4; B = 16'h00BE; #100;
A = 16'h00A4; B = 16'h00BF; #100;
A = 16'h00A4; B = 16'h00C0; #100;
A = 16'h00A4; B = 16'h00C1; #100;
A = 16'h00A4; B = 16'h00C2; #100;
A = 16'h00A4; B = 16'h00C3; #100;
A = 16'h00A4; B = 16'h00C4; #100;
A = 16'h00A4; B = 16'h00C5; #100;
A = 16'h00A4; B = 16'h00C6; #100;
A = 16'h00A4; B = 16'h00C7; #100;
A = 16'h00A4; B = 16'h00C8; #100;
A = 16'h00A4; B = 16'h00C9; #100;
A = 16'h00A4; B = 16'h00CA; #100;
A = 16'h00A4; B = 16'h00CB; #100;
A = 16'h00A4; B = 16'h00CC; #100;
A = 16'h00A4; B = 16'h00CD; #100;
A = 16'h00A4; B = 16'h00CE; #100;
A = 16'h00A4; B = 16'h00CF; #100;
A = 16'h00A4; B = 16'h00D0; #100;
A = 16'h00A4; B = 16'h00D1; #100;
A = 16'h00A4; B = 16'h00D2; #100;
A = 16'h00A4; B = 16'h00D3; #100;
A = 16'h00A4; B = 16'h00D4; #100;
A = 16'h00A4; B = 16'h00D5; #100;
A = 16'h00A4; B = 16'h00D6; #100;
A = 16'h00A4; B = 16'h00D7; #100;
A = 16'h00A4; B = 16'h00D8; #100;
A = 16'h00A4; B = 16'h00D9; #100;
A = 16'h00A4; B = 16'h00DA; #100;
A = 16'h00A4; B = 16'h00DB; #100;
A = 16'h00A4; B = 16'h00DC; #100;
A = 16'h00A4; B = 16'h00DD; #100;
A = 16'h00A4; B = 16'h00DE; #100;
A = 16'h00A4; B = 16'h00DF; #100;
A = 16'h00A4; B = 16'h00E0; #100;
A = 16'h00A4; B = 16'h00E1; #100;
A = 16'h00A4; B = 16'h00E2; #100;
A = 16'h00A4; B = 16'h00E3; #100;
A = 16'h00A4; B = 16'h00E4; #100;
A = 16'h00A4; B = 16'h00E5; #100;
A = 16'h00A4; B = 16'h00E6; #100;
A = 16'h00A4; B = 16'h00E7; #100;
A = 16'h00A4; B = 16'h00E8; #100;
A = 16'h00A4; B = 16'h00E9; #100;
A = 16'h00A4; B = 16'h00EA; #100;
A = 16'h00A4; B = 16'h00EB; #100;
A = 16'h00A4; B = 16'h00EC; #100;
A = 16'h00A4; B = 16'h00ED; #100;
A = 16'h00A4; B = 16'h00EE; #100;
A = 16'h00A4; B = 16'h00EF; #100;
A = 16'h00A4; B = 16'h00F0; #100;
A = 16'h00A4; B = 16'h00F1; #100;
A = 16'h00A4; B = 16'h00F2; #100;
A = 16'h00A4; B = 16'h00F3; #100;
A = 16'h00A4; B = 16'h00F4; #100;
A = 16'h00A4; B = 16'h00F5; #100;
A = 16'h00A4; B = 16'h00F6; #100;
A = 16'h00A4; B = 16'h00F7; #100;
A = 16'h00A4; B = 16'h00F8; #100;
A = 16'h00A4; B = 16'h00F9; #100;
A = 16'h00A4; B = 16'h00FA; #100;
A = 16'h00A4; B = 16'h00FB; #100;
A = 16'h00A4; B = 16'h00FC; #100;
A = 16'h00A4; B = 16'h00FD; #100;
A = 16'h00A4; B = 16'h00FE; #100;
A = 16'h00A4; B = 16'h00FF; #100;
A = 16'h00A5; B = 16'h000; #100;
A = 16'h00A5; B = 16'h001; #100;
A = 16'h00A5; B = 16'h002; #100;
A = 16'h00A5; B = 16'h003; #100;
A = 16'h00A5; B = 16'h004; #100;
A = 16'h00A5; B = 16'h005; #100;
A = 16'h00A5; B = 16'h006; #100;
A = 16'h00A5; B = 16'h007; #100;
A = 16'h00A5; B = 16'h008; #100;
A = 16'h00A5; B = 16'h009; #100;
A = 16'h00A5; B = 16'h00A; #100;
A = 16'h00A5; B = 16'h00B; #100;
A = 16'h00A5; B = 16'h00C; #100;
A = 16'h00A5; B = 16'h00D; #100;
A = 16'h00A5; B = 16'h00E; #100;
A = 16'h00A5; B = 16'h00F; #100;
A = 16'h00A5; B = 16'h0010; #100;
A = 16'h00A5; B = 16'h0011; #100;
A = 16'h00A5; B = 16'h0012; #100;
A = 16'h00A5; B = 16'h0013; #100;
A = 16'h00A5; B = 16'h0014; #100;
A = 16'h00A5; B = 16'h0015; #100;
A = 16'h00A5; B = 16'h0016; #100;
A = 16'h00A5; B = 16'h0017; #100;
A = 16'h00A5; B = 16'h0018; #100;
A = 16'h00A5; B = 16'h0019; #100;
A = 16'h00A5; B = 16'h001A; #100;
A = 16'h00A5; B = 16'h001B; #100;
A = 16'h00A5; B = 16'h001C; #100;
A = 16'h00A5; B = 16'h001D; #100;
A = 16'h00A5; B = 16'h001E; #100;
A = 16'h00A5; B = 16'h001F; #100;
A = 16'h00A5; B = 16'h0020; #100;
A = 16'h00A5; B = 16'h0021; #100;
A = 16'h00A5; B = 16'h0022; #100;
A = 16'h00A5; B = 16'h0023; #100;
A = 16'h00A5; B = 16'h0024; #100;
A = 16'h00A5; B = 16'h0025; #100;
A = 16'h00A5; B = 16'h0026; #100;
A = 16'h00A5; B = 16'h0027; #100;
A = 16'h00A5; B = 16'h0028; #100;
A = 16'h00A5; B = 16'h0029; #100;
A = 16'h00A5; B = 16'h002A; #100;
A = 16'h00A5; B = 16'h002B; #100;
A = 16'h00A5; B = 16'h002C; #100;
A = 16'h00A5; B = 16'h002D; #100;
A = 16'h00A5; B = 16'h002E; #100;
A = 16'h00A5; B = 16'h002F; #100;
A = 16'h00A5; B = 16'h0030; #100;
A = 16'h00A5; B = 16'h0031; #100;
A = 16'h00A5; B = 16'h0032; #100;
A = 16'h00A5; B = 16'h0033; #100;
A = 16'h00A5; B = 16'h0034; #100;
A = 16'h00A5; B = 16'h0035; #100;
A = 16'h00A5; B = 16'h0036; #100;
A = 16'h00A5; B = 16'h0037; #100;
A = 16'h00A5; B = 16'h0038; #100;
A = 16'h00A5; B = 16'h0039; #100;
A = 16'h00A5; B = 16'h003A; #100;
A = 16'h00A5; B = 16'h003B; #100;
A = 16'h00A5; B = 16'h003C; #100;
A = 16'h00A5; B = 16'h003D; #100;
A = 16'h00A5; B = 16'h003E; #100;
A = 16'h00A5; B = 16'h003F; #100;
A = 16'h00A5; B = 16'h0040; #100;
A = 16'h00A5; B = 16'h0041; #100;
A = 16'h00A5; B = 16'h0042; #100;
A = 16'h00A5; B = 16'h0043; #100;
A = 16'h00A5; B = 16'h0044; #100;
A = 16'h00A5; B = 16'h0045; #100;
A = 16'h00A5; B = 16'h0046; #100;
A = 16'h00A5; B = 16'h0047; #100;
A = 16'h00A5; B = 16'h0048; #100;
A = 16'h00A5; B = 16'h0049; #100;
A = 16'h00A5; B = 16'h004A; #100;
A = 16'h00A5; B = 16'h004B; #100;
A = 16'h00A5; B = 16'h004C; #100;
A = 16'h00A5; B = 16'h004D; #100;
A = 16'h00A5; B = 16'h004E; #100;
A = 16'h00A5; B = 16'h004F; #100;
A = 16'h00A5; B = 16'h0050; #100;
A = 16'h00A5; B = 16'h0051; #100;
A = 16'h00A5; B = 16'h0052; #100;
A = 16'h00A5; B = 16'h0053; #100;
A = 16'h00A5; B = 16'h0054; #100;
A = 16'h00A5; B = 16'h0055; #100;
A = 16'h00A5; B = 16'h0056; #100;
A = 16'h00A5; B = 16'h0057; #100;
A = 16'h00A5; B = 16'h0058; #100;
A = 16'h00A5; B = 16'h0059; #100;
A = 16'h00A5; B = 16'h005A; #100;
A = 16'h00A5; B = 16'h005B; #100;
A = 16'h00A5; B = 16'h005C; #100;
A = 16'h00A5; B = 16'h005D; #100;
A = 16'h00A5; B = 16'h005E; #100;
A = 16'h00A5; B = 16'h005F; #100;
A = 16'h00A5; B = 16'h0060; #100;
A = 16'h00A5; B = 16'h0061; #100;
A = 16'h00A5; B = 16'h0062; #100;
A = 16'h00A5; B = 16'h0063; #100;
A = 16'h00A5; B = 16'h0064; #100;
A = 16'h00A5; B = 16'h0065; #100;
A = 16'h00A5; B = 16'h0066; #100;
A = 16'h00A5; B = 16'h0067; #100;
A = 16'h00A5; B = 16'h0068; #100;
A = 16'h00A5; B = 16'h0069; #100;
A = 16'h00A5; B = 16'h006A; #100;
A = 16'h00A5; B = 16'h006B; #100;
A = 16'h00A5; B = 16'h006C; #100;
A = 16'h00A5; B = 16'h006D; #100;
A = 16'h00A5; B = 16'h006E; #100;
A = 16'h00A5; B = 16'h006F; #100;
A = 16'h00A5; B = 16'h0070; #100;
A = 16'h00A5; B = 16'h0071; #100;
A = 16'h00A5; B = 16'h0072; #100;
A = 16'h00A5; B = 16'h0073; #100;
A = 16'h00A5; B = 16'h0074; #100;
A = 16'h00A5; B = 16'h0075; #100;
A = 16'h00A5; B = 16'h0076; #100;
A = 16'h00A5; B = 16'h0077; #100;
A = 16'h00A5; B = 16'h0078; #100;
A = 16'h00A5; B = 16'h0079; #100;
A = 16'h00A5; B = 16'h007A; #100;
A = 16'h00A5; B = 16'h007B; #100;
A = 16'h00A5; B = 16'h007C; #100;
A = 16'h00A5; B = 16'h007D; #100;
A = 16'h00A5; B = 16'h007E; #100;
A = 16'h00A5; B = 16'h007F; #100;
A = 16'h00A5; B = 16'h0080; #100;
A = 16'h00A5; B = 16'h0081; #100;
A = 16'h00A5; B = 16'h0082; #100;
A = 16'h00A5; B = 16'h0083; #100;
A = 16'h00A5; B = 16'h0084; #100;
A = 16'h00A5; B = 16'h0085; #100;
A = 16'h00A5; B = 16'h0086; #100;
A = 16'h00A5; B = 16'h0087; #100;
A = 16'h00A5; B = 16'h0088; #100;
A = 16'h00A5; B = 16'h0089; #100;
A = 16'h00A5; B = 16'h008A; #100;
A = 16'h00A5; B = 16'h008B; #100;
A = 16'h00A5; B = 16'h008C; #100;
A = 16'h00A5; B = 16'h008D; #100;
A = 16'h00A5; B = 16'h008E; #100;
A = 16'h00A5; B = 16'h008F; #100;
A = 16'h00A5; B = 16'h0090; #100;
A = 16'h00A5; B = 16'h0091; #100;
A = 16'h00A5; B = 16'h0092; #100;
A = 16'h00A5; B = 16'h0093; #100;
A = 16'h00A5; B = 16'h0094; #100;
A = 16'h00A5; B = 16'h0095; #100;
A = 16'h00A5; B = 16'h0096; #100;
A = 16'h00A5; B = 16'h0097; #100;
A = 16'h00A5; B = 16'h0098; #100;
A = 16'h00A5; B = 16'h0099; #100;
A = 16'h00A5; B = 16'h009A; #100;
A = 16'h00A5; B = 16'h009B; #100;
A = 16'h00A5; B = 16'h009C; #100;
A = 16'h00A5; B = 16'h009D; #100;
A = 16'h00A5; B = 16'h009E; #100;
A = 16'h00A5; B = 16'h009F; #100;
A = 16'h00A5; B = 16'h00A0; #100;
A = 16'h00A5; B = 16'h00A1; #100;
A = 16'h00A5; B = 16'h00A2; #100;
A = 16'h00A5; B = 16'h00A3; #100;
A = 16'h00A5; B = 16'h00A4; #100;
A = 16'h00A5; B = 16'h00A5; #100;
A = 16'h00A5; B = 16'h00A6; #100;
A = 16'h00A5; B = 16'h00A7; #100;
A = 16'h00A5; B = 16'h00A8; #100;
A = 16'h00A5; B = 16'h00A9; #100;
A = 16'h00A5; B = 16'h00AA; #100;
A = 16'h00A5; B = 16'h00AB; #100;
A = 16'h00A5; B = 16'h00AC; #100;
A = 16'h00A5; B = 16'h00AD; #100;
A = 16'h00A5; B = 16'h00AE; #100;
A = 16'h00A5; B = 16'h00AF; #100;
A = 16'h00A5; B = 16'h00B0; #100;
A = 16'h00A5; B = 16'h00B1; #100;
A = 16'h00A5; B = 16'h00B2; #100;
A = 16'h00A5; B = 16'h00B3; #100;
A = 16'h00A5; B = 16'h00B4; #100;
A = 16'h00A5; B = 16'h00B5; #100;
A = 16'h00A5; B = 16'h00B6; #100;
A = 16'h00A5; B = 16'h00B7; #100;
A = 16'h00A5; B = 16'h00B8; #100;
A = 16'h00A5; B = 16'h00B9; #100;
A = 16'h00A5; B = 16'h00BA; #100;
A = 16'h00A5; B = 16'h00BB; #100;
A = 16'h00A5; B = 16'h00BC; #100;
A = 16'h00A5; B = 16'h00BD; #100;
A = 16'h00A5; B = 16'h00BE; #100;
A = 16'h00A5; B = 16'h00BF; #100;
A = 16'h00A5; B = 16'h00C0; #100;
A = 16'h00A5; B = 16'h00C1; #100;
A = 16'h00A5; B = 16'h00C2; #100;
A = 16'h00A5; B = 16'h00C3; #100;
A = 16'h00A5; B = 16'h00C4; #100;
A = 16'h00A5; B = 16'h00C5; #100;
A = 16'h00A5; B = 16'h00C6; #100;
A = 16'h00A5; B = 16'h00C7; #100;
A = 16'h00A5; B = 16'h00C8; #100;
A = 16'h00A5; B = 16'h00C9; #100;
A = 16'h00A5; B = 16'h00CA; #100;
A = 16'h00A5; B = 16'h00CB; #100;
A = 16'h00A5; B = 16'h00CC; #100;
A = 16'h00A5; B = 16'h00CD; #100;
A = 16'h00A5; B = 16'h00CE; #100;
A = 16'h00A5; B = 16'h00CF; #100;
A = 16'h00A5; B = 16'h00D0; #100;
A = 16'h00A5; B = 16'h00D1; #100;
A = 16'h00A5; B = 16'h00D2; #100;
A = 16'h00A5; B = 16'h00D3; #100;
A = 16'h00A5; B = 16'h00D4; #100;
A = 16'h00A5; B = 16'h00D5; #100;
A = 16'h00A5; B = 16'h00D6; #100;
A = 16'h00A5; B = 16'h00D7; #100;
A = 16'h00A5; B = 16'h00D8; #100;
A = 16'h00A5; B = 16'h00D9; #100;
A = 16'h00A5; B = 16'h00DA; #100;
A = 16'h00A5; B = 16'h00DB; #100;
A = 16'h00A5; B = 16'h00DC; #100;
A = 16'h00A5; B = 16'h00DD; #100;
A = 16'h00A5; B = 16'h00DE; #100;
A = 16'h00A5; B = 16'h00DF; #100;
A = 16'h00A5; B = 16'h00E0; #100;
A = 16'h00A5; B = 16'h00E1; #100;
A = 16'h00A5; B = 16'h00E2; #100;
A = 16'h00A5; B = 16'h00E3; #100;
A = 16'h00A5; B = 16'h00E4; #100;
A = 16'h00A5; B = 16'h00E5; #100;
A = 16'h00A5; B = 16'h00E6; #100;
A = 16'h00A5; B = 16'h00E7; #100;
A = 16'h00A5; B = 16'h00E8; #100;
A = 16'h00A5; B = 16'h00E9; #100;
A = 16'h00A5; B = 16'h00EA; #100;
A = 16'h00A5; B = 16'h00EB; #100;
A = 16'h00A5; B = 16'h00EC; #100;
A = 16'h00A5; B = 16'h00ED; #100;
A = 16'h00A5; B = 16'h00EE; #100;
A = 16'h00A5; B = 16'h00EF; #100;
A = 16'h00A5; B = 16'h00F0; #100;
A = 16'h00A5; B = 16'h00F1; #100;
A = 16'h00A5; B = 16'h00F2; #100;
A = 16'h00A5; B = 16'h00F3; #100;
A = 16'h00A5; B = 16'h00F4; #100;
A = 16'h00A5; B = 16'h00F5; #100;
A = 16'h00A5; B = 16'h00F6; #100;
A = 16'h00A5; B = 16'h00F7; #100;
A = 16'h00A5; B = 16'h00F8; #100;
A = 16'h00A5; B = 16'h00F9; #100;
A = 16'h00A5; B = 16'h00FA; #100;
A = 16'h00A5; B = 16'h00FB; #100;
A = 16'h00A5; B = 16'h00FC; #100;
A = 16'h00A5; B = 16'h00FD; #100;
A = 16'h00A5; B = 16'h00FE; #100;
A = 16'h00A5; B = 16'h00FF; #100;
A = 16'h00A6; B = 16'h000; #100;
A = 16'h00A6; B = 16'h001; #100;
A = 16'h00A6; B = 16'h002; #100;
A = 16'h00A6; B = 16'h003; #100;
A = 16'h00A6; B = 16'h004; #100;
A = 16'h00A6; B = 16'h005; #100;
A = 16'h00A6; B = 16'h006; #100;
A = 16'h00A6; B = 16'h007; #100;
A = 16'h00A6; B = 16'h008; #100;
A = 16'h00A6; B = 16'h009; #100;
A = 16'h00A6; B = 16'h00A; #100;
A = 16'h00A6; B = 16'h00B; #100;
A = 16'h00A6; B = 16'h00C; #100;
A = 16'h00A6; B = 16'h00D; #100;
A = 16'h00A6; B = 16'h00E; #100;
A = 16'h00A6; B = 16'h00F; #100;
A = 16'h00A6; B = 16'h0010; #100;
A = 16'h00A6; B = 16'h0011; #100;
A = 16'h00A6; B = 16'h0012; #100;
A = 16'h00A6; B = 16'h0013; #100;
A = 16'h00A6; B = 16'h0014; #100;
A = 16'h00A6; B = 16'h0015; #100;
A = 16'h00A6; B = 16'h0016; #100;
A = 16'h00A6; B = 16'h0017; #100;
A = 16'h00A6; B = 16'h0018; #100;
A = 16'h00A6; B = 16'h0019; #100;
A = 16'h00A6; B = 16'h001A; #100;
A = 16'h00A6; B = 16'h001B; #100;
A = 16'h00A6; B = 16'h001C; #100;
A = 16'h00A6; B = 16'h001D; #100;
A = 16'h00A6; B = 16'h001E; #100;
A = 16'h00A6; B = 16'h001F; #100;
A = 16'h00A6; B = 16'h0020; #100;
A = 16'h00A6; B = 16'h0021; #100;
A = 16'h00A6; B = 16'h0022; #100;
A = 16'h00A6; B = 16'h0023; #100;
A = 16'h00A6; B = 16'h0024; #100;
A = 16'h00A6; B = 16'h0025; #100;
A = 16'h00A6; B = 16'h0026; #100;
A = 16'h00A6; B = 16'h0027; #100;
A = 16'h00A6; B = 16'h0028; #100;
A = 16'h00A6; B = 16'h0029; #100;
A = 16'h00A6; B = 16'h002A; #100;
A = 16'h00A6; B = 16'h002B; #100;
A = 16'h00A6; B = 16'h002C; #100;
A = 16'h00A6; B = 16'h002D; #100;
A = 16'h00A6; B = 16'h002E; #100;
A = 16'h00A6; B = 16'h002F; #100;
A = 16'h00A6; B = 16'h0030; #100;
A = 16'h00A6; B = 16'h0031; #100;
A = 16'h00A6; B = 16'h0032; #100;
A = 16'h00A6; B = 16'h0033; #100;
A = 16'h00A6; B = 16'h0034; #100;
A = 16'h00A6; B = 16'h0035; #100;
A = 16'h00A6; B = 16'h0036; #100;
A = 16'h00A6; B = 16'h0037; #100;
A = 16'h00A6; B = 16'h0038; #100;
A = 16'h00A6; B = 16'h0039; #100;
A = 16'h00A6; B = 16'h003A; #100;
A = 16'h00A6; B = 16'h003B; #100;
A = 16'h00A6; B = 16'h003C; #100;
A = 16'h00A6; B = 16'h003D; #100;
A = 16'h00A6; B = 16'h003E; #100;
A = 16'h00A6; B = 16'h003F; #100;
A = 16'h00A6; B = 16'h0040; #100;
A = 16'h00A6; B = 16'h0041; #100;
A = 16'h00A6; B = 16'h0042; #100;
A = 16'h00A6; B = 16'h0043; #100;
A = 16'h00A6; B = 16'h0044; #100;
A = 16'h00A6; B = 16'h0045; #100;
A = 16'h00A6; B = 16'h0046; #100;
A = 16'h00A6; B = 16'h0047; #100;
A = 16'h00A6; B = 16'h0048; #100;
A = 16'h00A6; B = 16'h0049; #100;
A = 16'h00A6; B = 16'h004A; #100;
A = 16'h00A6; B = 16'h004B; #100;
A = 16'h00A6; B = 16'h004C; #100;
A = 16'h00A6; B = 16'h004D; #100;
A = 16'h00A6; B = 16'h004E; #100;
A = 16'h00A6; B = 16'h004F; #100;
A = 16'h00A6; B = 16'h0050; #100;
A = 16'h00A6; B = 16'h0051; #100;
A = 16'h00A6; B = 16'h0052; #100;
A = 16'h00A6; B = 16'h0053; #100;
A = 16'h00A6; B = 16'h0054; #100;
A = 16'h00A6; B = 16'h0055; #100;
A = 16'h00A6; B = 16'h0056; #100;
A = 16'h00A6; B = 16'h0057; #100;
A = 16'h00A6; B = 16'h0058; #100;
A = 16'h00A6; B = 16'h0059; #100;
A = 16'h00A6; B = 16'h005A; #100;
A = 16'h00A6; B = 16'h005B; #100;
A = 16'h00A6; B = 16'h005C; #100;
A = 16'h00A6; B = 16'h005D; #100;
A = 16'h00A6; B = 16'h005E; #100;
A = 16'h00A6; B = 16'h005F; #100;
A = 16'h00A6; B = 16'h0060; #100;
A = 16'h00A6; B = 16'h0061; #100;
A = 16'h00A6; B = 16'h0062; #100;
A = 16'h00A6; B = 16'h0063; #100;
A = 16'h00A6; B = 16'h0064; #100;
A = 16'h00A6; B = 16'h0065; #100;
A = 16'h00A6; B = 16'h0066; #100;
A = 16'h00A6; B = 16'h0067; #100;
A = 16'h00A6; B = 16'h0068; #100;
A = 16'h00A6; B = 16'h0069; #100;
A = 16'h00A6; B = 16'h006A; #100;
A = 16'h00A6; B = 16'h006B; #100;
A = 16'h00A6; B = 16'h006C; #100;
A = 16'h00A6; B = 16'h006D; #100;
A = 16'h00A6; B = 16'h006E; #100;
A = 16'h00A6; B = 16'h006F; #100;
A = 16'h00A6; B = 16'h0070; #100;
A = 16'h00A6; B = 16'h0071; #100;
A = 16'h00A6; B = 16'h0072; #100;
A = 16'h00A6; B = 16'h0073; #100;
A = 16'h00A6; B = 16'h0074; #100;
A = 16'h00A6; B = 16'h0075; #100;
A = 16'h00A6; B = 16'h0076; #100;
A = 16'h00A6; B = 16'h0077; #100;
A = 16'h00A6; B = 16'h0078; #100;
A = 16'h00A6; B = 16'h0079; #100;
A = 16'h00A6; B = 16'h007A; #100;
A = 16'h00A6; B = 16'h007B; #100;
A = 16'h00A6; B = 16'h007C; #100;
A = 16'h00A6; B = 16'h007D; #100;
A = 16'h00A6; B = 16'h007E; #100;
A = 16'h00A6; B = 16'h007F; #100;
A = 16'h00A6; B = 16'h0080; #100;
A = 16'h00A6; B = 16'h0081; #100;
A = 16'h00A6; B = 16'h0082; #100;
A = 16'h00A6; B = 16'h0083; #100;
A = 16'h00A6; B = 16'h0084; #100;
A = 16'h00A6; B = 16'h0085; #100;
A = 16'h00A6; B = 16'h0086; #100;
A = 16'h00A6; B = 16'h0087; #100;
A = 16'h00A6; B = 16'h0088; #100;
A = 16'h00A6; B = 16'h0089; #100;
A = 16'h00A6; B = 16'h008A; #100;
A = 16'h00A6; B = 16'h008B; #100;
A = 16'h00A6; B = 16'h008C; #100;
A = 16'h00A6; B = 16'h008D; #100;
A = 16'h00A6; B = 16'h008E; #100;
A = 16'h00A6; B = 16'h008F; #100;
A = 16'h00A6; B = 16'h0090; #100;
A = 16'h00A6; B = 16'h0091; #100;
A = 16'h00A6; B = 16'h0092; #100;
A = 16'h00A6; B = 16'h0093; #100;
A = 16'h00A6; B = 16'h0094; #100;
A = 16'h00A6; B = 16'h0095; #100;
A = 16'h00A6; B = 16'h0096; #100;
A = 16'h00A6; B = 16'h0097; #100;
A = 16'h00A6; B = 16'h0098; #100;
A = 16'h00A6; B = 16'h0099; #100;
A = 16'h00A6; B = 16'h009A; #100;
A = 16'h00A6; B = 16'h009B; #100;
A = 16'h00A6; B = 16'h009C; #100;
A = 16'h00A6; B = 16'h009D; #100;
A = 16'h00A6; B = 16'h009E; #100;
A = 16'h00A6; B = 16'h009F; #100;
A = 16'h00A6; B = 16'h00A0; #100;
A = 16'h00A6; B = 16'h00A1; #100;
A = 16'h00A6; B = 16'h00A2; #100;
A = 16'h00A6; B = 16'h00A3; #100;
A = 16'h00A6; B = 16'h00A4; #100;
A = 16'h00A6; B = 16'h00A5; #100;
A = 16'h00A6; B = 16'h00A6; #100;
A = 16'h00A6; B = 16'h00A7; #100;
A = 16'h00A6; B = 16'h00A8; #100;
A = 16'h00A6; B = 16'h00A9; #100;
A = 16'h00A6; B = 16'h00AA; #100;
A = 16'h00A6; B = 16'h00AB; #100;
A = 16'h00A6; B = 16'h00AC; #100;
A = 16'h00A6; B = 16'h00AD; #100;
A = 16'h00A6; B = 16'h00AE; #100;
A = 16'h00A6; B = 16'h00AF; #100;
A = 16'h00A6; B = 16'h00B0; #100;
A = 16'h00A6; B = 16'h00B1; #100;
A = 16'h00A6; B = 16'h00B2; #100;
A = 16'h00A6; B = 16'h00B3; #100;
A = 16'h00A6; B = 16'h00B4; #100;
A = 16'h00A6; B = 16'h00B5; #100;
A = 16'h00A6; B = 16'h00B6; #100;
A = 16'h00A6; B = 16'h00B7; #100;
A = 16'h00A6; B = 16'h00B8; #100;
A = 16'h00A6; B = 16'h00B9; #100;
A = 16'h00A6; B = 16'h00BA; #100;
A = 16'h00A6; B = 16'h00BB; #100;
A = 16'h00A6; B = 16'h00BC; #100;
A = 16'h00A6; B = 16'h00BD; #100;
A = 16'h00A6; B = 16'h00BE; #100;
A = 16'h00A6; B = 16'h00BF; #100;
A = 16'h00A6; B = 16'h00C0; #100;
A = 16'h00A6; B = 16'h00C1; #100;
A = 16'h00A6; B = 16'h00C2; #100;
A = 16'h00A6; B = 16'h00C3; #100;
A = 16'h00A6; B = 16'h00C4; #100;
A = 16'h00A6; B = 16'h00C5; #100;
A = 16'h00A6; B = 16'h00C6; #100;
A = 16'h00A6; B = 16'h00C7; #100;
A = 16'h00A6; B = 16'h00C8; #100;
A = 16'h00A6; B = 16'h00C9; #100;
A = 16'h00A6; B = 16'h00CA; #100;
A = 16'h00A6; B = 16'h00CB; #100;
A = 16'h00A6; B = 16'h00CC; #100;
A = 16'h00A6; B = 16'h00CD; #100;
A = 16'h00A6; B = 16'h00CE; #100;
A = 16'h00A6; B = 16'h00CF; #100;
A = 16'h00A6; B = 16'h00D0; #100;
A = 16'h00A6; B = 16'h00D1; #100;
A = 16'h00A6; B = 16'h00D2; #100;
A = 16'h00A6; B = 16'h00D3; #100;
A = 16'h00A6; B = 16'h00D4; #100;
A = 16'h00A6; B = 16'h00D5; #100;
A = 16'h00A6; B = 16'h00D6; #100;
A = 16'h00A6; B = 16'h00D7; #100;
A = 16'h00A6; B = 16'h00D8; #100;
A = 16'h00A6; B = 16'h00D9; #100;
A = 16'h00A6; B = 16'h00DA; #100;
A = 16'h00A6; B = 16'h00DB; #100;
A = 16'h00A6; B = 16'h00DC; #100;
A = 16'h00A6; B = 16'h00DD; #100;
A = 16'h00A6; B = 16'h00DE; #100;
A = 16'h00A6; B = 16'h00DF; #100;
A = 16'h00A6; B = 16'h00E0; #100;
A = 16'h00A6; B = 16'h00E1; #100;
A = 16'h00A6; B = 16'h00E2; #100;
A = 16'h00A6; B = 16'h00E3; #100;
A = 16'h00A6; B = 16'h00E4; #100;
A = 16'h00A6; B = 16'h00E5; #100;
A = 16'h00A6; B = 16'h00E6; #100;
A = 16'h00A6; B = 16'h00E7; #100;
A = 16'h00A6; B = 16'h00E8; #100;
A = 16'h00A6; B = 16'h00E9; #100;
A = 16'h00A6; B = 16'h00EA; #100;
A = 16'h00A6; B = 16'h00EB; #100;
A = 16'h00A6; B = 16'h00EC; #100;
A = 16'h00A6; B = 16'h00ED; #100;
A = 16'h00A6; B = 16'h00EE; #100;
A = 16'h00A6; B = 16'h00EF; #100;
A = 16'h00A6; B = 16'h00F0; #100;
A = 16'h00A6; B = 16'h00F1; #100;
A = 16'h00A6; B = 16'h00F2; #100;
A = 16'h00A6; B = 16'h00F3; #100;
A = 16'h00A6; B = 16'h00F4; #100;
A = 16'h00A6; B = 16'h00F5; #100;
A = 16'h00A6; B = 16'h00F6; #100;
A = 16'h00A6; B = 16'h00F7; #100;
A = 16'h00A6; B = 16'h00F8; #100;
A = 16'h00A6; B = 16'h00F9; #100;
A = 16'h00A6; B = 16'h00FA; #100;
A = 16'h00A6; B = 16'h00FB; #100;
A = 16'h00A6; B = 16'h00FC; #100;
A = 16'h00A6; B = 16'h00FD; #100;
A = 16'h00A6; B = 16'h00FE; #100;
A = 16'h00A6; B = 16'h00FF; #100;
A = 16'h00A7; B = 16'h000; #100;
A = 16'h00A7; B = 16'h001; #100;
A = 16'h00A7; B = 16'h002; #100;
A = 16'h00A7; B = 16'h003; #100;
A = 16'h00A7; B = 16'h004; #100;
A = 16'h00A7; B = 16'h005; #100;
A = 16'h00A7; B = 16'h006; #100;
A = 16'h00A7; B = 16'h007; #100;
A = 16'h00A7; B = 16'h008; #100;
A = 16'h00A7; B = 16'h009; #100;
A = 16'h00A7; B = 16'h00A; #100;
A = 16'h00A7; B = 16'h00B; #100;
A = 16'h00A7; B = 16'h00C; #100;
A = 16'h00A7; B = 16'h00D; #100;
A = 16'h00A7; B = 16'h00E; #100;
A = 16'h00A7; B = 16'h00F; #100;
A = 16'h00A7; B = 16'h0010; #100;
A = 16'h00A7; B = 16'h0011; #100;
A = 16'h00A7; B = 16'h0012; #100;
A = 16'h00A7; B = 16'h0013; #100;
A = 16'h00A7; B = 16'h0014; #100;
A = 16'h00A7; B = 16'h0015; #100;
A = 16'h00A7; B = 16'h0016; #100;
A = 16'h00A7; B = 16'h0017; #100;
A = 16'h00A7; B = 16'h0018; #100;
A = 16'h00A7; B = 16'h0019; #100;
A = 16'h00A7; B = 16'h001A; #100;
A = 16'h00A7; B = 16'h001B; #100;
A = 16'h00A7; B = 16'h001C; #100;
A = 16'h00A7; B = 16'h001D; #100;
A = 16'h00A7; B = 16'h001E; #100;
A = 16'h00A7; B = 16'h001F; #100;
A = 16'h00A7; B = 16'h0020; #100;
A = 16'h00A7; B = 16'h0021; #100;
A = 16'h00A7; B = 16'h0022; #100;
A = 16'h00A7; B = 16'h0023; #100;
A = 16'h00A7; B = 16'h0024; #100;
A = 16'h00A7; B = 16'h0025; #100;
A = 16'h00A7; B = 16'h0026; #100;
A = 16'h00A7; B = 16'h0027; #100;
A = 16'h00A7; B = 16'h0028; #100;
A = 16'h00A7; B = 16'h0029; #100;
A = 16'h00A7; B = 16'h002A; #100;
A = 16'h00A7; B = 16'h002B; #100;
A = 16'h00A7; B = 16'h002C; #100;
A = 16'h00A7; B = 16'h002D; #100;
A = 16'h00A7; B = 16'h002E; #100;
A = 16'h00A7; B = 16'h002F; #100;
A = 16'h00A7; B = 16'h0030; #100;
A = 16'h00A7; B = 16'h0031; #100;
A = 16'h00A7; B = 16'h0032; #100;
A = 16'h00A7; B = 16'h0033; #100;
A = 16'h00A7; B = 16'h0034; #100;
A = 16'h00A7; B = 16'h0035; #100;
A = 16'h00A7; B = 16'h0036; #100;
A = 16'h00A7; B = 16'h0037; #100;
A = 16'h00A7; B = 16'h0038; #100;
A = 16'h00A7; B = 16'h0039; #100;
A = 16'h00A7; B = 16'h003A; #100;
A = 16'h00A7; B = 16'h003B; #100;
A = 16'h00A7; B = 16'h003C; #100;
A = 16'h00A7; B = 16'h003D; #100;
A = 16'h00A7; B = 16'h003E; #100;
A = 16'h00A7; B = 16'h003F; #100;
A = 16'h00A7; B = 16'h0040; #100;
A = 16'h00A7; B = 16'h0041; #100;
A = 16'h00A7; B = 16'h0042; #100;
A = 16'h00A7; B = 16'h0043; #100;
A = 16'h00A7; B = 16'h0044; #100;
A = 16'h00A7; B = 16'h0045; #100;
A = 16'h00A7; B = 16'h0046; #100;
A = 16'h00A7; B = 16'h0047; #100;
A = 16'h00A7; B = 16'h0048; #100;
A = 16'h00A7; B = 16'h0049; #100;
A = 16'h00A7; B = 16'h004A; #100;
A = 16'h00A7; B = 16'h004B; #100;
A = 16'h00A7; B = 16'h004C; #100;
A = 16'h00A7; B = 16'h004D; #100;
A = 16'h00A7; B = 16'h004E; #100;
A = 16'h00A7; B = 16'h004F; #100;
A = 16'h00A7; B = 16'h0050; #100;
A = 16'h00A7; B = 16'h0051; #100;
A = 16'h00A7; B = 16'h0052; #100;
A = 16'h00A7; B = 16'h0053; #100;
A = 16'h00A7; B = 16'h0054; #100;
A = 16'h00A7; B = 16'h0055; #100;
A = 16'h00A7; B = 16'h0056; #100;
A = 16'h00A7; B = 16'h0057; #100;
A = 16'h00A7; B = 16'h0058; #100;
A = 16'h00A7; B = 16'h0059; #100;
A = 16'h00A7; B = 16'h005A; #100;
A = 16'h00A7; B = 16'h005B; #100;
A = 16'h00A7; B = 16'h005C; #100;
A = 16'h00A7; B = 16'h005D; #100;
A = 16'h00A7; B = 16'h005E; #100;
A = 16'h00A7; B = 16'h005F; #100;
A = 16'h00A7; B = 16'h0060; #100;
A = 16'h00A7; B = 16'h0061; #100;
A = 16'h00A7; B = 16'h0062; #100;
A = 16'h00A7; B = 16'h0063; #100;
A = 16'h00A7; B = 16'h0064; #100;
A = 16'h00A7; B = 16'h0065; #100;
A = 16'h00A7; B = 16'h0066; #100;
A = 16'h00A7; B = 16'h0067; #100;
A = 16'h00A7; B = 16'h0068; #100;
A = 16'h00A7; B = 16'h0069; #100;
A = 16'h00A7; B = 16'h006A; #100;
A = 16'h00A7; B = 16'h006B; #100;
A = 16'h00A7; B = 16'h006C; #100;
A = 16'h00A7; B = 16'h006D; #100;
A = 16'h00A7; B = 16'h006E; #100;
A = 16'h00A7; B = 16'h006F; #100;
A = 16'h00A7; B = 16'h0070; #100;
A = 16'h00A7; B = 16'h0071; #100;
A = 16'h00A7; B = 16'h0072; #100;
A = 16'h00A7; B = 16'h0073; #100;
A = 16'h00A7; B = 16'h0074; #100;
A = 16'h00A7; B = 16'h0075; #100;
A = 16'h00A7; B = 16'h0076; #100;
A = 16'h00A7; B = 16'h0077; #100;
A = 16'h00A7; B = 16'h0078; #100;
A = 16'h00A7; B = 16'h0079; #100;
A = 16'h00A7; B = 16'h007A; #100;
A = 16'h00A7; B = 16'h007B; #100;
A = 16'h00A7; B = 16'h007C; #100;
A = 16'h00A7; B = 16'h007D; #100;
A = 16'h00A7; B = 16'h007E; #100;
A = 16'h00A7; B = 16'h007F; #100;
A = 16'h00A7; B = 16'h0080; #100;
A = 16'h00A7; B = 16'h0081; #100;
A = 16'h00A7; B = 16'h0082; #100;
A = 16'h00A7; B = 16'h0083; #100;
A = 16'h00A7; B = 16'h0084; #100;
A = 16'h00A7; B = 16'h0085; #100;
A = 16'h00A7; B = 16'h0086; #100;
A = 16'h00A7; B = 16'h0087; #100;
A = 16'h00A7; B = 16'h0088; #100;
A = 16'h00A7; B = 16'h0089; #100;
A = 16'h00A7; B = 16'h008A; #100;
A = 16'h00A7; B = 16'h008B; #100;
A = 16'h00A7; B = 16'h008C; #100;
A = 16'h00A7; B = 16'h008D; #100;
A = 16'h00A7; B = 16'h008E; #100;
A = 16'h00A7; B = 16'h008F; #100;
A = 16'h00A7; B = 16'h0090; #100;
A = 16'h00A7; B = 16'h0091; #100;
A = 16'h00A7; B = 16'h0092; #100;
A = 16'h00A7; B = 16'h0093; #100;
A = 16'h00A7; B = 16'h0094; #100;
A = 16'h00A7; B = 16'h0095; #100;
A = 16'h00A7; B = 16'h0096; #100;
A = 16'h00A7; B = 16'h0097; #100;
A = 16'h00A7; B = 16'h0098; #100;
A = 16'h00A7; B = 16'h0099; #100;
A = 16'h00A7; B = 16'h009A; #100;
A = 16'h00A7; B = 16'h009B; #100;
A = 16'h00A7; B = 16'h009C; #100;
A = 16'h00A7; B = 16'h009D; #100;
A = 16'h00A7; B = 16'h009E; #100;
A = 16'h00A7; B = 16'h009F; #100;
A = 16'h00A7; B = 16'h00A0; #100;
A = 16'h00A7; B = 16'h00A1; #100;
A = 16'h00A7; B = 16'h00A2; #100;
A = 16'h00A7; B = 16'h00A3; #100;
A = 16'h00A7; B = 16'h00A4; #100;
A = 16'h00A7; B = 16'h00A5; #100;
A = 16'h00A7; B = 16'h00A6; #100;
A = 16'h00A7; B = 16'h00A7; #100;
A = 16'h00A7; B = 16'h00A8; #100;
A = 16'h00A7; B = 16'h00A9; #100;
A = 16'h00A7; B = 16'h00AA; #100;
A = 16'h00A7; B = 16'h00AB; #100;
A = 16'h00A7; B = 16'h00AC; #100;
A = 16'h00A7; B = 16'h00AD; #100;
A = 16'h00A7; B = 16'h00AE; #100;
A = 16'h00A7; B = 16'h00AF; #100;
A = 16'h00A7; B = 16'h00B0; #100;
A = 16'h00A7; B = 16'h00B1; #100;
A = 16'h00A7; B = 16'h00B2; #100;
A = 16'h00A7; B = 16'h00B3; #100;
A = 16'h00A7; B = 16'h00B4; #100;
A = 16'h00A7; B = 16'h00B5; #100;
A = 16'h00A7; B = 16'h00B6; #100;
A = 16'h00A7; B = 16'h00B7; #100;
A = 16'h00A7; B = 16'h00B8; #100;
A = 16'h00A7; B = 16'h00B9; #100;
A = 16'h00A7; B = 16'h00BA; #100;
A = 16'h00A7; B = 16'h00BB; #100;
A = 16'h00A7; B = 16'h00BC; #100;
A = 16'h00A7; B = 16'h00BD; #100;
A = 16'h00A7; B = 16'h00BE; #100;
A = 16'h00A7; B = 16'h00BF; #100;
A = 16'h00A7; B = 16'h00C0; #100;
A = 16'h00A7; B = 16'h00C1; #100;
A = 16'h00A7; B = 16'h00C2; #100;
A = 16'h00A7; B = 16'h00C3; #100;
A = 16'h00A7; B = 16'h00C4; #100;
A = 16'h00A7; B = 16'h00C5; #100;
A = 16'h00A7; B = 16'h00C6; #100;
A = 16'h00A7; B = 16'h00C7; #100;
A = 16'h00A7; B = 16'h00C8; #100;
A = 16'h00A7; B = 16'h00C9; #100;
A = 16'h00A7; B = 16'h00CA; #100;
A = 16'h00A7; B = 16'h00CB; #100;
A = 16'h00A7; B = 16'h00CC; #100;
A = 16'h00A7; B = 16'h00CD; #100;
A = 16'h00A7; B = 16'h00CE; #100;
A = 16'h00A7; B = 16'h00CF; #100;
A = 16'h00A7; B = 16'h00D0; #100;
A = 16'h00A7; B = 16'h00D1; #100;
A = 16'h00A7; B = 16'h00D2; #100;
A = 16'h00A7; B = 16'h00D3; #100;
A = 16'h00A7; B = 16'h00D4; #100;
A = 16'h00A7; B = 16'h00D5; #100;
A = 16'h00A7; B = 16'h00D6; #100;
A = 16'h00A7; B = 16'h00D7; #100;
A = 16'h00A7; B = 16'h00D8; #100;
A = 16'h00A7; B = 16'h00D9; #100;
A = 16'h00A7; B = 16'h00DA; #100;
A = 16'h00A7; B = 16'h00DB; #100;
A = 16'h00A7; B = 16'h00DC; #100;
A = 16'h00A7; B = 16'h00DD; #100;
A = 16'h00A7; B = 16'h00DE; #100;
A = 16'h00A7; B = 16'h00DF; #100;
A = 16'h00A7; B = 16'h00E0; #100;
A = 16'h00A7; B = 16'h00E1; #100;
A = 16'h00A7; B = 16'h00E2; #100;
A = 16'h00A7; B = 16'h00E3; #100;
A = 16'h00A7; B = 16'h00E4; #100;
A = 16'h00A7; B = 16'h00E5; #100;
A = 16'h00A7; B = 16'h00E6; #100;
A = 16'h00A7; B = 16'h00E7; #100;
A = 16'h00A7; B = 16'h00E8; #100;
A = 16'h00A7; B = 16'h00E9; #100;
A = 16'h00A7; B = 16'h00EA; #100;
A = 16'h00A7; B = 16'h00EB; #100;
A = 16'h00A7; B = 16'h00EC; #100;
A = 16'h00A7; B = 16'h00ED; #100;
A = 16'h00A7; B = 16'h00EE; #100;
A = 16'h00A7; B = 16'h00EF; #100;
A = 16'h00A7; B = 16'h00F0; #100;
A = 16'h00A7; B = 16'h00F1; #100;
A = 16'h00A7; B = 16'h00F2; #100;
A = 16'h00A7; B = 16'h00F3; #100;
A = 16'h00A7; B = 16'h00F4; #100;
A = 16'h00A7; B = 16'h00F5; #100;
A = 16'h00A7; B = 16'h00F6; #100;
A = 16'h00A7; B = 16'h00F7; #100;
A = 16'h00A7; B = 16'h00F8; #100;
A = 16'h00A7; B = 16'h00F9; #100;
A = 16'h00A7; B = 16'h00FA; #100;
A = 16'h00A7; B = 16'h00FB; #100;
A = 16'h00A7; B = 16'h00FC; #100;
A = 16'h00A7; B = 16'h00FD; #100;
A = 16'h00A7; B = 16'h00FE; #100;
A = 16'h00A7; B = 16'h00FF; #100;
A = 16'h00A8; B = 16'h000; #100;
A = 16'h00A8; B = 16'h001; #100;
A = 16'h00A8; B = 16'h002; #100;
A = 16'h00A8; B = 16'h003; #100;
A = 16'h00A8; B = 16'h004; #100;
A = 16'h00A8; B = 16'h005; #100;
A = 16'h00A8; B = 16'h006; #100;
A = 16'h00A8; B = 16'h007; #100;
A = 16'h00A8; B = 16'h008; #100;
A = 16'h00A8; B = 16'h009; #100;
A = 16'h00A8; B = 16'h00A; #100;
A = 16'h00A8; B = 16'h00B; #100;
A = 16'h00A8; B = 16'h00C; #100;
A = 16'h00A8; B = 16'h00D; #100;
A = 16'h00A8; B = 16'h00E; #100;
A = 16'h00A8; B = 16'h00F; #100;
A = 16'h00A8; B = 16'h0010; #100;
A = 16'h00A8; B = 16'h0011; #100;
A = 16'h00A8; B = 16'h0012; #100;
A = 16'h00A8; B = 16'h0013; #100;
A = 16'h00A8; B = 16'h0014; #100;
A = 16'h00A8; B = 16'h0015; #100;
A = 16'h00A8; B = 16'h0016; #100;
A = 16'h00A8; B = 16'h0017; #100;
A = 16'h00A8; B = 16'h0018; #100;
A = 16'h00A8; B = 16'h0019; #100;
A = 16'h00A8; B = 16'h001A; #100;
A = 16'h00A8; B = 16'h001B; #100;
A = 16'h00A8; B = 16'h001C; #100;
A = 16'h00A8; B = 16'h001D; #100;
A = 16'h00A8; B = 16'h001E; #100;
A = 16'h00A8; B = 16'h001F; #100;
A = 16'h00A8; B = 16'h0020; #100;
A = 16'h00A8; B = 16'h0021; #100;
A = 16'h00A8; B = 16'h0022; #100;
A = 16'h00A8; B = 16'h0023; #100;
A = 16'h00A8; B = 16'h0024; #100;
A = 16'h00A8; B = 16'h0025; #100;
A = 16'h00A8; B = 16'h0026; #100;
A = 16'h00A8; B = 16'h0027; #100;
A = 16'h00A8; B = 16'h0028; #100;
A = 16'h00A8; B = 16'h0029; #100;
A = 16'h00A8; B = 16'h002A; #100;
A = 16'h00A8; B = 16'h002B; #100;
A = 16'h00A8; B = 16'h002C; #100;
A = 16'h00A8; B = 16'h002D; #100;
A = 16'h00A8; B = 16'h002E; #100;
A = 16'h00A8; B = 16'h002F; #100;
A = 16'h00A8; B = 16'h0030; #100;
A = 16'h00A8; B = 16'h0031; #100;
A = 16'h00A8; B = 16'h0032; #100;
A = 16'h00A8; B = 16'h0033; #100;
A = 16'h00A8; B = 16'h0034; #100;
A = 16'h00A8; B = 16'h0035; #100;
A = 16'h00A8; B = 16'h0036; #100;
A = 16'h00A8; B = 16'h0037; #100;
A = 16'h00A8; B = 16'h0038; #100;
A = 16'h00A8; B = 16'h0039; #100;
A = 16'h00A8; B = 16'h003A; #100;
A = 16'h00A8; B = 16'h003B; #100;
A = 16'h00A8; B = 16'h003C; #100;
A = 16'h00A8; B = 16'h003D; #100;
A = 16'h00A8; B = 16'h003E; #100;
A = 16'h00A8; B = 16'h003F; #100;
A = 16'h00A8; B = 16'h0040; #100;
A = 16'h00A8; B = 16'h0041; #100;
A = 16'h00A8; B = 16'h0042; #100;
A = 16'h00A8; B = 16'h0043; #100;
A = 16'h00A8; B = 16'h0044; #100;
A = 16'h00A8; B = 16'h0045; #100;
A = 16'h00A8; B = 16'h0046; #100;
A = 16'h00A8; B = 16'h0047; #100;
A = 16'h00A8; B = 16'h0048; #100;
A = 16'h00A8; B = 16'h0049; #100;
A = 16'h00A8; B = 16'h004A; #100;
A = 16'h00A8; B = 16'h004B; #100;
A = 16'h00A8; B = 16'h004C; #100;
A = 16'h00A8; B = 16'h004D; #100;
A = 16'h00A8; B = 16'h004E; #100;
A = 16'h00A8; B = 16'h004F; #100;
A = 16'h00A8; B = 16'h0050; #100;
A = 16'h00A8; B = 16'h0051; #100;
A = 16'h00A8; B = 16'h0052; #100;
A = 16'h00A8; B = 16'h0053; #100;
A = 16'h00A8; B = 16'h0054; #100;
A = 16'h00A8; B = 16'h0055; #100;
A = 16'h00A8; B = 16'h0056; #100;
A = 16'h00A8; B = 16'h0057; #100;
A = 16'h00A8; B = 16'h0058; #100;
A = 16'h00A8; B = 16'h0059; #100;
A = 16'h00A8; B = 16'h005A; #100;
A = 16'h00A8; B = 16'h005B; #100;
A = 16'h00A8; B = 16'h005C; #100;
A = 16'h00A8; B = 16'h005D; #100;
A = 16'h00A8; B = 16'h005E; #100;
A = 16'h00A8; B = 16'h005F; #100;
A = 16'h00A8; B = 16'h0060; #100;
A = 16'h00A8; B = 16'h0061; #100;
A = 16'h00A8; B = 16'h0062; #100;
A = 16'h00A8; B = 16'h0063; #100;
A = 16'h00A8; B = 16'h0064; #100;
A = 16'h00A8; B = 16'h0065; #100;
A = 16'h00A8; B = 16'h0066; #100;
A = 16'h00A8; B = 16'h0067; #100;
A = 16'h00A8; B = 16'h0068; #100;
A = 16'h00A8; B = 16'h0069; #100;
A = 16'h00A8; B = 16'h006A; #100;
A = 16'h00A8; B = 16'h006B; #100;
A = 16'h00A8; B = 16'h006C; #100;
A = 16'h00A8; B = 16'h006D; #100;
A = 16'h00A8; B = 16'h006E; #100;
A = 16'h00A8; B = 16'h006F; #100;
A = 16'h00A8; B = 16'h0070; #100;
A = 16'h00A8; B = 16'h0071; #100;
A = 16'h00A8; B = 16'h0072; #100;
A = 16'h00A8; B = 16'h0073; #100;
A = 16'h00A8; B = 16'h0074; #100;
A = 16'h00A8; B = 16'h0075; #100;
A = 16'h00A8; B = 16'h0076; #100;
A = 16'h00A8; B = 16'h0077; #100;
A = 16'h00A8; B = 16'h0078; #100;
A = 16'h00A8; B = 16'h0079; #100;
A = 16'h00A8; B = 16'h007A; #100;
A = 16'h00A8; B = 16'h007B; #100;
A = 16'h00A8; B = 16'h007C; #100;
A = 16'h00A8; B = 16'h007D; #100;
A = 16'h00A8; B = 16'h007E; #100;
A = 16'h00A8; B = 16'h007F; #100;
A = 16'h00A8; B = 16'h0080; #100;
A = 16'h00A8; B = 16'h0081; #100;
A = 16'h00A8; B = 16'h0082; #100;
A = 16'h00A8; B = 16'h0083; #100;
A = 16'h00A8; B = 16'h0084; #100;
A = 16'h00A8; B = 16'h0085; #100;
A = 16'h00A8; B = 16'h0086; #100;
A = 16'h00A8; B = 16'h0087; #100;
A = 16'h00A8; B = 16'h0088; #100;
A = 16'h00A8; B = 16'h0089; #100;
A = 16'h00A8; B = 16'h008A; #100;
A = 16'h00A8; B = 16'h008B; #100;
A = 16'h00A8; B = 16'h008C; #100;
A = 16'h00A8; B = 16'h008D; #100;
A = 16'h00A8; B = 16'h008E; #100;
A = 16'h00A8; B = 16'h008F; #100;
A = 16'h00A8; B = 16'h0090; #100;
A = 16'h00A8; B = 16'h0091; #100;
A = 16'h00A8; B = 16'h0092; #100;
A = 16'h00A8; B = 16'h0093; #100;
A = 16'h00A8; B = 16'h0094; #100;
A = 16'h00A8; B = 16'h0095; #100;
A = 16'h00A8; B = 16'h0096; #100;
A = 16'h00A8; B = 16'h0097; #100;
A = 16'h00A8; B = 16'h0098; #100;
A = 16'h00A8; B = 16'h0099; #100;
A = 16'h00A8; B = 16'h009A; #100;
A = 16'h00A8; B = 16'h009B; #100;
A = 16'h00A8; B = 16'h009C; #100;
A = 16'h00A8; B = 16'h009D; #100;
A = 16'h00A8; B = 16'h009E; #100;
A = 16'h00A8; B = 16'h009F; #100;
A = 16'h00A8; B = 16'h00A0; #100;
A = 16'h00A8; B = 16'h00A1; #100;
A = 16'h00A8; B = 16'h00A2; #100;
A = 16'h00A8; B = 16'h00A3; #100;
A = 16'h00A8; B = 16'h00A4; #100;
A = 16'h00A8; B = 16'h00A5; #100;
A = 16'h00A8; B = 16'h00A6; #100;
A = 16'h00A8; B = 16'h00A7; #100;
A = 16'h00A8; B = 16'h00A8; #100;
A = 16'h00A8; B = 16'h00A9; #100;
A = 16'h00A8; B = 16'h00AA; #100;
A = 16'h00A8; B = 16'h00AB; #100;
A = 16'h00A8; B = 16'h00AC; #100;
A = 16'h00A8; B = 16'h00AD; #100;
A = 16'h00A8; B = 16'h00AE; #100;
A = 16'h00A8; B = 16'h00AF; #100;
A = 16'h00A8; B = 16'h00B0; #100;
A = 16'h00A8; B = 16'h00B1; #100;
A = 16'h00A8; B = 16'h00B2; #100;
A = 16'h00A8; B = 16'h00B3; #100;
A = 16'h00A8; B = 16'h00B4; #100;
A = 16'h00A8; B = 16'h00B5; #100;
A = 16'h00A8; B = 16'h00B6; #100;
A = 16'h00A8; B = 16'h00B7; #100;
A = 16'h00A8; B = 16'h00B8; #100;
A = 16'h00A8; B = 16'h00B9; #100;
A = 16'h00A8; B = 16'h00BA; #100;
A = 16'h00A8; B = 16'h00BB; #100;
A = 16'h00A8; B = 16'h00BC; #100;
A = 16'h00A8; B = 16'h00BD; #100;
A = 16'h00A8; B = 16'h00BE; #100;
A = 16'h00A8; B = 16'h00BF; #100;
A = 16'h00A8; B = 16'h00C0; #100;
A = 16'h00A8; B = 16'h00C1; #100;
A = 16'h00A8; B = 16'h00C2; #100;
A = 16'h00A8; B = 16'h00C3; #100;
A = 16'h00A8; B = 16'h00C4; #100;
A = 16'h00A8; B = 16'h00C5; #100;
A = 16'h00A8; B = 16'h00C6; #100;
A = 16'h00A8; B = 16'h00C7; #100;
A = 16'h00A8; B = 16'h00C8; #100;
A = 16'h00A8; B = 16'h00C9; #100;
A = 16'h00A8; B = 16'h00CA; #100;
A = 16'h00A8; B = 16'h00CB; #100;
A = 16'h00A8; B = 16'h00CC; #100;
A = 16'h00A8; B = 16'h00CD; #100;
A = 16'h00A8; B = 16'h00CE; #100;
A = 16'h00A8; B = 16'h00CF; #100;
A = 16'h00A8; B = 16'h00D0; #100;
A = 16'h00A8; B = 16'h00D1; #100;
A = 16'h00A8; B = 16'h00D2; #100;
A = 16'h00A8; B = 16'h00D3; #100;
A = 16'h00A8; B = 16'h00D4; #100;
A = 16'h00A8; B = 16'h00D5; #100;
A = 16'h00A8; B = 16'h00D6; #100;
A = 16'h00A8; B = 16'h00D7; #100;
A = 16'h00A8; B = 16'h00D8; #100;
A = 16'h00A8; B = 16'h00D9; #100;
A = 16'h00A8; B = 16'h00DA; #100;
A = 16'h00A8; B = 16'h00DB; #100;
A = 16'h00A8; B = 16'h00DC; #100;
A = 16'h00A8; B = 16'h00DD; #100;
A = 16'h00A8; B = 16'h00DE; #100;
A = 16'h00A8; B = 16'h00DF; #100;
A = 16'h00A8; B = 16'h00E0; #100;
A = 16'h00A8; B = 16'h00E1; #100;
A = 16'h00A8; B = 16'h00E2; #100;
A = 16'h00A8; B = 16'h00E3; #100;
A = 16'h00A8; B = 16'h00E4; #100;
A = 16'h00A8; B = 16'h00E5; #100;
A = 16'h00A8; B = 16'h00E6; #100;
A = 16'h00A8; B = 16'h00E7; #100;
A = 16'h00A8; B = 16'h00E8; #100;
A = 16'h00A8; B = 16'h00E9; #100;
A = 16'h00A8; B = 16'h00EA; #100;
A = 16'h00A8; B = 16'h00EB; #100;
A = 16'h00A8; B = 16'h00EC; #100;
A = 16'h00A8; B = 16'h00ED; #100;
A = 16'h00A8; B = 16'h00EE; #100;
A = 16'h00A8; B = 16'h00EF; #100;
A = 16'h00A8; B = 16'h00F0; #100;
A = 16'h00A8; B = 16'h00F1; #100;
A = 16'h00A8; B = 16'h00F2; #100;
A = 16'h00A8; B = 16'h00F3; #100;
A = 16'h00A8; B = 16'h00F4; #100;
A = 16'h00A8; B = 16'h00F5; #100;
A = 16'h00A8; B = 16'h00F6; #100;
A = 16'h00A8; B = 16'h00F7; #100;
A = 16'h00A8; B = 16'h00F8; #100;
A = 16'h00A8; B = 16'h00F9; #100;
A = 16'h00A8; B = 16'h00FA; #100;
A = 16'h00A8; B = 16'h00FB; #100;
A = 16'h00A8; B = 16'h00FC; #100;
A = 16'h00A8; B = 16'h00FD; #100;
A = 16'h00A8; B = 16'h00FE; #100;
A = 16'h00A8; B = 16'h00FF; #100;
A = 16'h00A9; B = 16'h000; #100;
A = 16'h00A9; B = 16'h001; #100;
A = 16'h00A9; B = 16'h002; #100;
A = 16'h00A9; B = 16'h003; #100;
A = 16'h00A9; B = 16'h004; #100;
A = 16'h00A9; B = 16'h005; #100;
A = 16'h00A9; B = 16'h006; #100;
A = 16'h00A9; B = 16'h007; #100;
A = 16'h00A9; B = 16'h008; #100;
A = 16'h00A9; B = 16'h009; #100;
A = 16'h00A9; B = 16'h00A; #100;
A = 16'h00A9; B = 16'h00B; #100;
A = 16'h00A9; B = 16'h00C; #100;
A = 16'h00A9; B = 16'h00D; #100;
A = 16'h00A9; B = 16'h00E; #100;
A = 16'h00A9; B = 16'h00F; #100;
A = 16'h00A9; B = 16'h0010; #100;
A = 16'h00A9; B = 16'h0011; #100;
A = 16'h00A9; B = 16'h0012; #100;
A = 16'h00A9; B = 16'h0013; #100;
A = 16'h00A9; B = 16'h0014; #100;
A = 16'h00A9; B = 16'h0015; #100;
A = 16'h00A9; B = 16'h0016; #100;
A = 16'h00A9; B = 16'h0017; #100;
A = 16'h00A9; B = 16'h0018; #100;
A = 16'h00A9; B = 16'h0019; #100;
A = 16'h00A9; B = 16'h001A; #100;
A = 16'h00A9; B = 16'h001B; #100;
A = 16'h00A9; B = 16'h001C; #100;
A = 16'h00A9; B = 16'h001D; #100;
A = 16'h00A9; B = 16'h001E; #100;
A = 16'h00A9; B = 16'h001F; #100;
A = 16'h00A9; B = 16'h0020; #100;
A = 16'h00A9; B = 16'h0021; #100;
A = 16'h00A9; B = 16'h0022; #100;
A = 16'h00A9; B = 16'h0023; #100;
A = 16'h00A9; B = 16'h0024; #100;
A = 16'h00A9; B = 16'h0025; #100;
A = 16'h00A9; B = 16'h0026; #100;
A = 16'h00A9; B = 16'h0027; #100;
A = 16'h00A9; B = 16'h0028; #100;
A = 16'h00A9; B = 16'h0029; #100;
A = 16'h00A9; B = 16'h002A; #100;
A = 16'h00A9; B = 16'h002B; #100;
A = 16'h00A9; B = 16'h002C; #100;
A = 16'h00A9; B = 16'h002D; #100;
A = 16'h00A9; B = 16'h002E; #100;
A = 16'h00A9; B = 16'h002F; #100;
A = 16'h00A9; B = 16'h0030; #100;
A = 16'h00A9; B = 16'h0031; #100;
A = 16'h00A9; B = 16'h0032; #100;
A = 16'h00A9; B = 16'h0033; #100;
A = 16'h00A9; B = 16'h0034; #100;
A = 16'h00A9; B = 16'h0035; #100;
A = 16'h00A9; B = 16'h0036; #100;
A = 16'h00A9; B = 16'h0037; #100;
A = 16'h00A9; B = 16'h0038; #100;
A = 16'h00A9; B = 16'h0039; #100;
A = 16'h00A9; B = 16'h003A; #100;
A = 16'h00A9; B = 16'h003B; #100;
A = 16'h00A9; B = 16'h003C; #100;
A = 16'h00A9; B = 16'h003D; #100;
A = 16'h00A9; B = 16'h003E; #100;
A = 16'h00A9; B = 16'h003F; #100;
A = 16'h00A9; B = 16'h0040; #100;
A = 16'h00A9; B = 16'h0041; #100;
A = 16'h00A9; B = 16'h0042; #100;
A = 16'h00A9; B = 16'h0043; #100;
A = 16'h00A9; B = 16'h0044; #100;
A = 16'h00A9; B = 16'h0045; #100;
A = 16'h00A9; B = 16'h0046; #100;
A = 16'h00A9; B = 16'h0047; #100;
A = 16'h00A9; B = 16'h0048; #100;
A = 16'h00A9; B = 16'h0049; #100;
A = 16'h00A9; B = 16'h004A; #100;
A = 16'h00A9; B = 16'h004B; #100;
A = 16'h00A9; B = 16'h004C; #100;
A = 16'h00A9; B = 16'h004D; #100;
A = 16'h00A9; B = 16'h004E; #100;
A = 16'h00A9; B = 16'h004F; #100;
A = 16'h00A9; B = 16'h0050; #100;
A = 16'h00A9; B = 16'h0051; #100;
A = 16'h00A9; B = 16'h0052; #100;
A = 16'h00A9; B = 16'h0053; #100;
A = 16'h00A9; B = 16'h0054; #100;
A = 16'h00A9; B = 16'h0055; #100;
A = 16'h00A9; B = 16'h0056; #100;
A = 16'h00A9; B = 16'h0057; #100;
A = 16'h00A9; B = 16'h0058; #100;
A = 16'h00A9; B = 16'h0059; #100;
A = 16'h00A9; B = 16'h005A; #100;
A = 16'h00A9; B = 16'h005B; #100;
A = 16'h00A9; B = 16'h005C; #100;
A = 16'h00A9; B = 16'h005D; #100;
A = 16'h00A9; B = 16'h005E; #100;
A = 16'h00A9; B = 16'h005F; #100;
A = 16'h00A9; B = 16'h0060; #100;
A = 16'h00A9; B = 16'h0061; #100;
A = 16'h00A9; B = 16'h0062; #100;
A = 16'h00A9; B = 16'h0063; #100;
A = 16'h00A9; B = 16'h0064; #100;
A = 16'h00A9; B = 16'h0065; #100;
A = 16'h00A9; B = 16'h0066; #100;
A = 16'h00A9; B = 16'h0067; #100;
A = 16'h00A9; B = 16'h0068; #100;
A = 16'h00A9; B = 16'h0069; #100;
A = 16'h00A9; B = 16'h006A; #100;
A = 16'h00A9; B = 16'h006B; #100;
A = 16'h00A9; B = 16'h006C; #100;
A = 16'h00A9; B = 16'h006D; #100;
A = 16'h00A9; B = 16'h006E; #100;
A = 16'h00A9; B = 16'h006F; #100;
A = 16'h00A9; B = 16'h0070; #100;
A = 16'h00A9; B = 16'h0071; #100;
A = 16'h00A9; B = 16'h0072; #100;
A = 16'h00A9; B = 16'h0073; #100;
A = 16'h00A9; B = 16'h0074; #100;
A = 16'h00A9; B = 16'h0075; #100;
A = 16'h00A9; B = 16'h0076; #100;
A = 16'h00A9; B = 16'h0077; #100;
A = 16'h00A9; B = 16'h0078; #100;
A = 16'h00A9; B = 16'h0079; #100;
A = 16'h00A9; B = 16'h007A; #100;
A = 16'h00A9; B = 16'h007B; #100;
A = 16'h00A9; B = 16'h007C; #100;
A = 16'h00A9; B = 16'h007D; #100;
A = 16'h00A9; B = 16'h007E; #100;
A = 16'h00A9; B = 16'h007F; #100;
A = 16'h00A9; B = 16'h0080; #100;
A = 16'h00A9; B = 16'h0081; #100;
A = 16'h00A9; B = 16'h0082; #100;
A = 16'h00A9; B = 16'h0083; #100;
A = 16'h00A9; B = 16'h0084; #100;
A = 16'h00A9; B = 16'h0085; #100;
A = 16'h00A9; B = 16'h0086; #100;
A = 16'h00A9; B = 16'h0087; #100;
A = 16'h00A9; B = 16'h0088; #100;
A = 16'h00A9; B = 16'h0089; #100;
A = 16'h00A9; B = 16'h008A; #100;
A = 16'h00A9; B = 16'h008B; #100;
A = 16'h00A9; B = 16'h008C; #100;
A = 16'h00A9; B = 16'h008D; #100;
A = 16'h00A9; B = 16'h008E; #100;
A = 16'h00A9; B = 16'h008F; #100;
A = 16'h00A9; B = 16'h0090; #100;
A = 16'h00A9; B = 16'h0091; #100;
A = 16'h00A9; B = 16'h0092; #100;
A = 16'h00A9; B = 16'h0093; #100;
A = 16'h00A9; B = 16'h0094; #100;
A = 16'h00A9; B = 16'h0095; #100;
A = 16'h00A9; B = 16'h0096; #100;
A = 16'h00A9; B = 16'h0097; #100;
A = 16'h00A9; B = 16'h0098; #100;
A = 16'h00A9; B = 16'h0099; #100;
A = 16'h00A9; B = 16'h009A; #100;
A = 16'h00A9; B = 16'h009B; #100;
A = 16'h00A9; B = 16'h009C; #100;
A = 16'h00A9; B = 16'h009D; #100;
A = 16'h00A9; B = 16'h009E; #100;
A = 16'h00A9; B = 16'h009F; #100;
A = 16'h00A9; B = 16'h00A0; #100;
A = 16'h00A9; B = 16'h00A1; #100;
A = 16'h00A9; B = 16'h00A2; #100;
A = 16'h00A9; B = 16'h00A3; #100;
A = 16'h00A9; B = 16'h00A4; #100;
A = 16'h00A9; B = 16'h00A5; #100;
A = 16'h00A9; B = 16'h00A6; #100;
A = 16'h00A9; B = 16'h00A7; #100;
A = 16'h00A9; B = 16'h00A8; #100;
A = 16'h00A9; B = 16'h00A9; #100;
A = 16'h00A9; B = 16'h00AA; #100;
A = 16'h00A9; B = 16'h00AB; #100;
A = 16'h00A9; B = 16'h00AC; #100;
A = 16'h00A9; B = 16'h00AD; #100;
A = 16'h00A9; B = 16'h00AE; #100;
A = 16'h00A9; B = 16'h00AF; #100;
A = 16'h00A9; B = 16'h00B0; #100;
A = 16'h00A9; B = 16'h00B1; #100;
A = 16'h00A9; B = 16'h00B2; #100;
A = 16'h00A9; B = 16'h00B3; #100;
A = 16'h00A9; B = 16'h00B4; #100;
A = 16'h00A9; B = 16'h00B5; #100;
A = 16'h00A9; B = 16'h00B6; #100;
A = 16'h00A9; B = 16'h00B7; #100;
A = 16'h00A9; B = 16'h00B8; #100;
A = 16'h00A9; B = 16'h00B9; #100;
A = 16'h00A9; B = 16'h00BA; #100;
A = 16'h00A9; B = 16'h00BB; #100;
A = 16'h00A9; B = 16'h00BC; #100;
A = 16'h00A9; B = 16'h00BD; #100;
A = 16'h00A9; B = 16'h00BE; #100;
A = 16'h00A9; B = 16'h00BF; #100;
A = 16'h00A9; B = 16'h00C0; #100;
A = 16'h00A9; B = 16'h00C1; #100;
A = 16'h00A9; B = 16'h00C2; #100;
A = 16'h00A9; B = 16'h00C3; #100;
A = 16'h00A9; B = 16'h00C4; #100;
A = 16'h00A9; B = 16'h00C5; #100;
A = 16'h00A9; B = 16'h00C6; #100;
A = 16'h00A9; B = 16'h00C7; #100;
A = 16'h00A9; B = 16'h00C8; #100;
A = 16'h00A9; B = 16'h00C9; #100;
A = 16'h00A9; B = 16'h00CA; #100;
A = 16'h00A9; B = 16'h00CB; #100;
A = 16'h00A9; B = 16'h00CC; #100;
A = 16'h00A9; B = 16'h00CD; #100;
A = 16'h00A9; B = 16'h00CE; #100;
A = 16'h00A9; B = 16'h00CF; #100;
A = 16'h00A9; B = 16'h00D0; #100;
A = 16'h00A9; B = 16'h00D1; #100;
A = 16'h00A9; B = 16'h00D2; #100;
A = 16'h00A9; B = 16'h00D3; #100;
A = 16'h00A9; B = 16'h00D4; #100;
A = 16'h00A9; B = 16'h00D5; #100;
A = 16'h00A9; B = 16'h00D6; #100;
A = 16'h00A9; B = 16'h00D7; #100;
A = 16'h00A9; B = 16'h00D8; #100;
A = 16'h00A9; B = 16'h00D9; #100;
A = 16'h00A9; B = 16'h00DA; #100;
A = 16'h00A9; B = 16'h00DB; #100;
A = 16'h00A9; B = 16'h00DC; #100;
A = 16'h00A9; B = 16'h00DD; #100;
A = 16'h00A9; B = 16'h00DE; #100;
A = 16'h00A9; B = 16'h00DF; #100;
A = 16'h00A9; B = 16'h00E0; #100;
A = 16'h00A9; B = 16'h00E1; #100;
A = 16'h00A9; B = 16'h00E2; #100;
A = 16'h00A9; B = 16'h00E3; #100;
A = 16'h00A9; B = 16'h00E4; #100;
A = 16'h00A9; B = 16'h00E5; #100;
A = 16'h00A9; B = 16'h00E6; #100;
A = 16'h00A9; B = 16'h00E7; #100;
A = 16'h00A9; B = 16'h00E8; #100;
A = 16'h00A9; B = 16'h00E9; #100;
A = 16'h00A9; B = 16'h00EA; #100;
A = 16'h00A9; B = 16'h00EB; #100;
A = 16'h00A9; B = 16'h00EC; #100;
A = 16'h00A9; B = 16'h00ED; #100;
A = 16'h00A9; B = 16'h00EE; #100;
A = 16'h00A9; B = 16'h00EF; #100;
A = 16'h00A9; B = 16'h00F0; #100;
A = 16'h00A9; B = 16'h00F1; #100;
A = 16'h00A9; B = 16'h00F2; #100;
A = 16'h00A9; B = 16'h00F3; #100;
A = 16'h00A9; B = 16'h00F4; #100;
A = 16'h00A9; B = 16'h00F5; #100;
A = 16'h00A9; B = 16'h00F6; #100;
A = 16'h00A9; B = 16'h00F7; #100;
A = 16'h00A9; B = 16'h00F8; #100;
A = 16'h00A9; B = 16'h00F9; #100;
A = 16'h00A9; B = 16'h00FA; #100;
A = 16'h00A9; B = 16'h00FB; #100;
A = 16'h00A9; B = 16'h00FC; #100;
A = 16'h00A9; B = 16'h00FD; #100;
A = 16'h00A9; B = 16'h00FE; #100;
A = 16'h00A9; B = 16'h00FF; #100;
A = 16'h00AA; B = 16'h000; #100;
A = 16'h00AA; B = 16'h001; #100;
A = 16'h00AA; B = 16'h002; #100;
A = 16'h00AA; B = 16'h003; #100;
A = 16'h00AA; B = 16'h004; #100;
A = 16'h00AA; B = 16'h005; #100;
A = 16'h00AA; B = 16'h006; #100;
A = 16'h00AA; B = 16'h007; #100;
A = 16'h00AA; B = 16'h008; #100;
A = 16'h00AA; B = 16'h009; #100;
A = 16'h00AA; B = 16'h00A; #100;
A = 16'h00AA; B = 16'h00B; #100;
A = 16'h00AA; B = 16'h00C; #100;
A = 16'h00AA; B = 16'h00D; #100;
A = 16'h00AA; B = 16'h00E; #100;
A = 16'h00AA; B = 16'h00F; #100;
A = 16'h00AA; B = 16'h0010; #100;
A = 16'h00AA; B = 16'h0011; #100;
A = 16'h00AA; B = 16'h0012; #100;
A = 16'h00AA; B = 16'h0013; #100;
A = 16'h00AA; B = 16'h0014; #100;
A = 16'h00AA; B = 16'h0015; #100;
A = 16'h00AA; B = 16'h0016; #100;
A = 16'h00AA; B = 16'h0017; #100;
A = 16'h00AA; B = 16'h0018; #100;
A = 16'h00AA; B = 16'h0019; #100;
A = 16'h00AA; B = 16'h001A; #100;
A = 16'h00AA; B = 16'h001B; #100;
A = 16'h00AA; B = 16'h001C; #100;
A = 16'h00AA; B = 16'h001D; #100;
A = 16'h00AA; B = 16'h001E; #100;
A = 16'h00AA; B = 16'h001F; #100;
A = 16'h00AA; B = 16'h0020; #100;
A = 16'h00AA; B = 16'h0021; #100;
A = 16'h00AA; B = 16'h0022; #100;
A = 16'h00AA; B = 16'h0023; #100;
A = 16'h00AA; B = 16'h0024; #100;
A = 16'h00AA; B = 16'h0025; #100;
A = 16'h00AA; B = 16'h0026; #100;
A = 16'h00AA; B = 16'h0027; #100;
A = 16'h00AA; B = 16'h0028; #100;
A = 16'h00AA; B = 16'h0029; #100;
A = 16'h00AA; B = 16'h002A; #100;
A = 16'h00AA; B = 16'h002B; #100;
A = 16'h00AA; B = 16'h002C; #100;
A = 16'h00AA; B = 16'h002D; #100;
A = 16'h00AA; B = 16'h002E; #100;
A = 16'h00AA; B = 16'h002F; #100;
A = 16'h00AA; B = 16'h0030; #100;
A = 16'h00AA; B = 16'h0031; #100;
A = 16'h00AA; B = 16'h0032; #100;
A = 16'h00AA; B = 16'h0033; #100;
A = 16'h00AA; B = 16'h0034; #100;
A = 16'h00AA; B = 16'h0035; #100;
A = 16'h00AA; B = 16'h0036; #100;
A = 16'h00AA; B = 16'h0037; #100;
A = 16'h00AA; B = 16'h0038; #100;
A = 16'h00AA; B = 16'h0039; #100;
A = 16'h00AA; B = 16'h003A; #100;
A = 16'h00AA; B = 16'h003B; #100;
A = 16'h00AA; B = 16'h003C; #100;
A = 16'h00AA; B = 16'h003D; #100;
A = 16'h00AA; B = 16'h003E; #100;
A = 16'h00AA; B = 16'h003F; #100;
A = 16'h00AA; B = 16'h0040; #100;
A = 16'h00AA; B = 16'h0041; #100;
A = 16'h00AA; B = 16'h0042; #100;
A = 16'h00AA; B = 16'h0043; #100;
A = 16'h00AA; B = 16'h0044; #100;
A = 16'h00AA; B = 16'h0045; #100;
A = 16'h00AA; B = 16'h0046; #100;
A = 16'h00AA; B = 16'h0047; #100;
A = 16'h00AA; B = 16'h0048; #100;
A = 16'h00AA; B = 16'h0049; #100;
A = 16'h00AA; B = 16'h004A; #100;
A = 16'h00AA; B = 16'h004B; #100;
A = 16'h00AA; B = 16'h004C; #100;
A = 16'h00AA; B = 16'h004D; #100;
A = 16'h00AA; B = 16'h004E; #100;
A = 16'h00AA; B = 16'h004F; #100;
A = 16'h00AA; B = 16'h0050; #100;
A = 16'h00AA; B = 16'h0051; #100;
A = 16'h00AA; B = 16'h0052; #100;
A = 16'h00AA; B = 16'h0053; #100;
A = 16'h00AA; B = 16'h0054; #100;
A = 16'h00AA; B = 16'h0055; #100;
A = 16'h00AA; B = 16'h0056; #100;
A = 16'h00AA; B = 16'h0057; #100;
A = 16'h00AA; B = 16'h0058; #100;
A = 16'h00AA; B = 16'h0059; #100;
A = 16'h00AA; B = 16'h005A; #100;
A = 16'h00AA; B = 16'h005B; #100;
A = 16'h00AA; B = 16'h005C; #100;
A = 16'h00AA; B = 16'h005D; #100;
A = 16'h00AA; B = 16'h005E; #100;
A = 16'h00AA; B = 16'h005F; #100;
A = 16'h00AA; B = 16'h0060; #100;
A = 16'h00AA; B = 16'h0061; #100;
A = 16'h00AA; B = 16'h0062; #100;
A = 16'h00AA; B = 16'h0063; #100;
A = 16'h00AA; B = 16'h0064; #100;
A = 16'h00AA; B = 16'h0065; #100;
A = 16'h00AA; B = 16'h0066; #100;
A = 16'h00AA; B = 16'h0067; #100;
A = 16'h00AA; B = 16'h0068; #100;
A = 16'h00AA; B = 16'h0069; #100;
A = 16'h00AA; B = 16'h006A; #100;
A = 16'h00AA; B = 16'h006B; #100;
A = 16'h00AA; B = 16'h006C; #100;
A = 16'h00AA; B = 16'h006D; #100;
A = 16'h00AA; B = 16'h006E; #100;
A = 16'h00AA; B = 16'h006F; #100;
A = 16'h00AA; B = 16'h0070; #100;
A = 16'h00AA; B = 16'h0071; #100;
A = 16'h00AA; B = 16'h0072; #100;
A = 16'h00AA; B = 16'h0073; #100;
A = 16'h00AA; B = 16'h0074; #100;
A = 16'h00AA; B = 16'h0075; #100;
A = 16'h00AA; B = 16'h0076; #100;
A = 16'h00AA; B = 16'h0077; #100;
A = 16'h00AA; B = 16'h0078; #100;
A = 16'h00AA; B = 16'h0079; #100;
A = 16'h00AA; B = 16'h007A; #100;
A = 16'h00AA; B = 16'h007B; #100;
A = 16'h00AA; B = 16'h007C; #100;
A = 16'h00AA; B = 16'h007D; #100;
A = 16'h00AA; B = 16'h007E; #100;
A = 16'h00AA; B = 16'h007F; #100;
A = 16'h00AA; B = 16'h0080; #100;
A = 16'h00AA; B = 16'h0081; #100;
A = 16'h00AA; B = 16'h0082; #100;
A = 16'h00AA; B = 16'h0083; #100;
A = 16'h00AA; B = 16'h0084; #100;
A = 16'h00AA; B = 16'h0085; #100;
A = 16'h00AA; B = 16'h0086; #100;
A = 16'h00AA; B = 16'h0087; #100;
A = 16'h00AA; B = 16'h0088; #100;
A = 16'h00AA; B = 16'h0089; #100;
A = 16'h00AA; B = 16'h008A; #100;
A = 16'h00AA; B = 16'h008B; #100;
A = 16'h00AA; B = 16'h008C; #100;
A = 16'h00AA; B = 16'h008D; #100;
A = 16'h00AA; B = 16'h008E; #100;
A = 16'h00AA; B = 16'h008F; #100;
A = 16'h00AA; B = 16'h0090; #100;
A = 16'h00AA; B = 16'h0091; #100;
A = 16'h00AA; B = 16'h0092; #100;
A = 16'h00AA; B = 16'h0093; #100;
A = 16'h00AA; B = 16'h0094; #100;
A = 16'h00AA; B = 16'h0095; #100;
A = 16'h00AA; B = 16'h0096; #100;
A = 16'h00AA; B = 16'h0097; #100;
A = 16'h00AA; B = 16'h0098; #100;
A = 16'h00AA; B = 16'h0099; #100;
A = 16'h00AA; B = 16'h009A; #100;
A = 16'h00AA; B = 16'h009B; #100;
A = 16'h00AA; B = 16'h009C; #100;
A = 16'h00AA; B = 16'h009D; #100;
A = 16'h00AA; B = 16'h009E; #100;
A = 16'h00AA; B = 16'h009F; #100;
A = 16'h00AA; B = 16'h00A0; #100;
A = 16'h00AA; B = 16'h00A1; #100;
A = 16'h00AA; B = 16'h00A2; #100;
A = 16'h00AA; B = 16'h00A3; #100;
A = 16'h00AA; B = 16'h00A4; #100;
A = 16'h00AA; B = 16'h00A5; #100;
A = 16'h00AA; B = 16'h00A6; #100;
A = 16'h00AA; B = 16'h00A7; #100;
A = 16'h00AA; B = 16'h00A8; #100;
A = 16'h00AA; B = 16'h00A9; #100;
A = 16'h00AA; B = 16'h00AA; #100;
A = 16'h00AA; B = 16'h00AB; #100;
A = 16'h00AA; B = 16'h00AC; #100;
A = 16'h00AA; B = 16'h00AD; #100;
A = 16'h00AA; B = 16'h00AE; #100;
A = 16'h00AA; B = 16'h00AF; #100;
A = 16'h00AA; B = 16'h00B0; #100;
A = 16'h00AA; B = 16'h00B1; #100;
A = 16'h00AA; B = 16'h00B2; #100;
A = 16'h00AA; B = 16'h00B3; #100;
A = 16'h00AA; B = 16'h00B4; #100;
A = 16'h00AA; B = 16'h00B5; #100;
A = 16'h00AA; B = 16'h00B6; #100;
A = 16'h00AA; B = 16'h00B7; #100;
A = 16'h00AA; B = 16'h00B8; #100;
A = 16'h00AA; B = 16'h00B9; #100;
A = 16'h00AA; B = 16'h00BA; #100;
A = 16'h00AA; B = 16'h00BB; #100;
A = 16'h00AA; B = 16'h00BC; #100;
A = 16'h00AA; B = 16'h00BD; #100;
A = 16'h00AA; B = 16'h00BE; #100;
A = 16'h00AA; B = 16'h00BF; #100;
A = 16'h00AA; B = 16'h00C0; #100;
A = 16'h00AA; B = 16'h00C1; #100;
A = 16'h00AA; B = 16'h00C2; #100;
A = 16'h00AA; B = 16'h00C3; #100;
A = 16'h00AA; B = 16'h00C4; #100;
A = 16'h00AA; B = 16'h00C5; #100;
A = 16'h00AA; B = 16'h00C6; #100;
A = 16'h00AA; B = 16'h00C7; #100;
A = 16'h00AA; B = 16'h00C8; #100;
A = 16'h00AA; B = 16'h00C9; #100;
A = 16'h00AA; B = 16'h00CA; #100;
A = 16'h00AA; B = 16'h00CB; #100;
A = 16'h00AA; B = 16'h00CC; #100;
A = 16'h00AA; B = 16'h00CD; #100;
A = 16'h00AA; B = 16'h00CE; #100;
A = 16'h00AA; B = 16'h00CF; #100;
A = 16'h00AA; B = 16'h00D0; #100;
A = 16'h00AA; B = 16'h00D1; #100;
A = 16'h00AA; B = 16'h00D2; #100;
A = 16'h00AA; B = 16'h00D3; #100;
A = 16'h00AA; B = 16'h00D4; #100;
A = 16'h00AA; B = 16'h00D5; #100;
A = 16'h00AA; B = 16'h00D6; #100;
A = 16'h00AA; B = 16'h00D7; #100;
A = 16'h00AA; B = 16'h00D8; #100;
A = 16'h00AA; B = 16'h00D9; #100;
A = 16'h00AA; B = 16'h00DA; #100;
A = 16'h00AA; B = 16'h00DB; #100;
A = 16'h00AA; B = 16'h00DC; #100;
A = 16'h00AA; B = 16'h00DD; #100;
A = 16'h00AA; B = 16'h00DE; #100;
A = 16'h00AA; B = 16'h00DF; #100;
A = 16'h00AA; B = 16'h00E0; #100;
A = 16'h00AA; B = 16'h00E1; #100;
A = 16'h00AA; B = 16'h00E2; #100;
A = 16'h00AA; B = 16'h00E3; #100;
A = 16'h00AA; B = 16'h00E4; #100;
A = 16'h00AA; B = 16'h00E5; #100;
A = 16'h00AA; B = 16'h00E6; #100;
A = 16'h00AA; B = 16'h00E7; #100;
A = 16'h00AA; B = 16'h00E8; #100;
A = 16'h00AA; B = 16'h00E9; #100;
A = 16'h00AA; B = 16'h00EA; #100;
A = 16'h00AA; B = 16'h00EB; #100;
A = 16'h00AA; B = 16'h00EC; #100;
A = 16'h00AA; B = 16'h00ED; #100;
A = 16'h00AA; B = 16'h00EE; #100;
A = 16'h00AA; B = 16'h00EF; #100;
A = 16'h00AA; B = 16'h00F0; #100;
A = 16'h00AA; B = 16'h00F1; #100;
A = 16'h00AA; B = 16'h00F2; #100;
A = 16'h00AA; B = 16'h00F3; #100;
A = 16'h00AA; B = 16'h00F4; #100;
A = 16'h00AA; B = 16'h00F5; #100;
A = 16'h00AA; B = 16'h00F6; #100;
A = 16'h00AA; B = 16'h00F7; #100;
A = 16'h00AA; B = 16'h00F8; #100;
A = 16'h00AA; B = 16'h00F9; #100;
A = 16'h00AA; B = 16'h00FA; #100;
A = 16'h00AA; B = 16'h00FB; #100;
A = 16'h00AA; B = 16'h00FC; #100;
A = 16'h00AA; B = 16'h00FD; #100;
A = 16'h00AA; B = 16'h00FE; #100;
A = 16'h00AA; B = 16'h00FF; #100;
A = 16'h00AB; B = 16'h000; #100;
A = 16'h00AB; B = 16'h001; #100;
A = 16'h00AB; B = 16'h002; #100;
A = 16'h00AB; B = 16'h003; #100;
A = 16'h00AB; B = 16'h004; #100;
A = 16'h00AB; B = 16'h005; #100;
A = 16'h00AB; B = 16'h006; #100;
A = 16'h00AB; B = 16'h007; #100;
A = 16'h00AB; B = 16'h008; #100;
A = 16'h00AB; B = 16'h009; #100;
A = 16'h00AB; B = 16'h00A; #100;
A = 16'h00AB; B = 16'h00B; #100;
A = 16'h00AB; B = 16'h00C; #100;
A = 16'h00AB; B = 16'h00D; #100;
A = 16'h00AB; B = 16'h00E; #100;
A = 16'h00AB; B = 16'h00F; #100;
A = 16'h00AB; B = 16'h0010; #100;
A = 16'h00AB; B = 16'h0011; #100;
A = 16'h00AB; B = 16'h0012; #100;
A = 16'h00AB; B = 16'h0013; #100;
A = 16'h00AB; B = 16'h0014; #100;
A = 16'h00AB; B = 16'h0015; #100;
A = 16'h00AB; B = 16'h0016; #100;
A = 16'h00AB; B = 16'h0017; #100;
A = 16'h00AB; B = 16'h0018; #100;
A = 16'h00AB; B = 16'h0019; #100;
A = 16'h00AB; B = 16'h001A; #100;
A = 16'h00AB; B = 16'h001B; #100;
A = 16'h00AB; B = 16'h001C; #100;
A = 16'h00AB; B = 16'h001D; #100;
A = 16'h00AB; B = 16'h001E; #100;
A = 16'h00AB; B = 16'h001F; #100;
A = 16'h00AB; B = 16'h0020; #100;
A = 16'h00AB; B = 16'h0021; #100;
A = 16'h00AB; B = 16'h0022; #100;
A = 16'h00AB; B = 16'h0023; #100;
A = 16'h00AB; B = 16'h0024; #100;
A = 16'h00AB; B = 16'h0025; #100;
A = 16'h00AB; B = 16'h0026; #100;
A = 16'h00AB; B = 16'h0027; #100;
A = 16'h00AB; B = 16'h0028; #100;
A = 16'h00AB; B = 16'h0029; #100;
A = 16'h00AB; B = 16'h002A; #100;
A = 16'h00AB; B = 16'h002B; #100;
A = 16'h00AB; B = 16'h002C; #100;
A = 16'h00AB; B = 16'h002D; #100;
A = 16'h00AB; B = 16'h002E; #100;
A = 16'h00AB; B = 16'h002F; #100;
A = 16'h00AB; B = 16'h0030; #100;
A = 16'h00AB; B = 16'h0031; #100;
A = 16'h00AB; B = 16'h0032; #100;
A = 16'h00AB; B = 16'h0033; #100;
A = 16'h00AB; B = 16'h0034; #100;
A = 16'h00AB; B = 16'h0035; #100;
A = 16'h00AB; B = 16'h0036; #100;
A = 16'h00AB; B = 16'h0037; #100;
A = 16'h00AB; B = 16'h0038; #100;
A = 16'h00AB; B = 16'h0039; #100;
A = 16'h00AB; B = 16'h003A; #100;
A = 16'h00AB; B = 16'h003B; #100;
A = 16'h00AB; B = 16'h003C; #100;
A = 16'h00AB; B = 16'h003D; #100;
A = 16'h00AB; B = 16'h003E; #100;
A = 16'h00AB; B = 16'h003F; #100;
A = 16'h00AB; B = 16'h0040; #100;
A = 16'h00AB; B = 16'h0041; #100;
A = 16'h00AB; B = 16'h0042; #100;
A = 16'h00AB; B = 16'h0043; #100;
A = 16'h00AB; B = 16'h0044; #100;
A = 16'h00AB; B = 16'h0045; #100;
A = 16'h00AB; B = 16'h0046; #100;
A = 16'h00AB; B = 16'h0047; #100;
A = 16'h00AB; B = 16'h0048; #100;
A = 16'h00AB; B = 16'h0049; #100;
A = 16'h00AB; B = 16'h004A; #100;
A = 16'h00AB; B = 16'h004B; #100;
A = 16'h00AB; B = 16'h004C; #100;
A = 16'h00AB; B = 16'h004D; #100;
A = 16'h00AB; B = 16'h004E; #100;
A = 16'h00AB; B = 16'h004F; #100;
A = 16'h00AB; B = 16'h0050; #100;
A = 16'h00AB; B = 16'h0051; #100;
A = 16'h00AB; B = 16'h0052; #100;
A = 16'h00AB; B = 16'h0053; #100;
A = 16'h00AB; B = 16'h0054; #100;
A = 16'h00AB; B = 16'h0055; #100;
A = 16'h00AB; B = 16'h0056; #100;
A = 16'h00AB; B = 16'h0057; #100;
A = 16'h00AB; B = 16'h0058; #100;
A = 16'h00AB; B = 16'h0059; #100;
A = 16'h00AB; B = 16'h005A; #100;
A = 16'h00AB; B = 16'h005B; #100;
A = 16'h00AB; B = 16'h005C; #100;
A = 16'h00AB; B = 16'h005D; #100;
A = 16'h00AB; B = 16'h005E; #100;
A = 16'h00AB; B = 16'h005F; #100;
A = 16'h00AB; B = 16'h0060; #100;
A = 16'h00AB; B = 16'h0061; #100;
A = 16'h00AB; B = 16'h0062; #100;
A = 16'h00AB; B = 16'h0063; #100;
A = 16'h00AB; B = 16'h0064; #100;
A = 16'h00AB; B = 16'h0065; #100;
A = 16'h00AB; B = 16'h0066; #100;
A = 16'h00AB; B = 16'h0067; #100;
A = 16'h00AB; B = 16'h0068; #100;
A = 16'h00AB; B = 16'h0069; #100;
A = 16'h00AB; B = 16'h006A; #100;
A = 16'h00AB; B = 16'h006B; #100;
A = 16'h00AB; B = 16'h006C; #100;
A = 16'h00AB; B = 16'h006D; #100;
A = 16'h00AB; B = 16'h006E; #100;
A = 16'h00AB; B = 16'h006F; #100;
A = 16'h00AB; B = 16'h0070; #100;
A = 16'h00AB; B = 16'h0071; #100;
A = 16'h00AB; B = 16'h0072; #100;
A = 16'h00AB; B = 16'h0073; #100;
A = 16'h00AB; B = 16'h0074; #100;
A = 16'h00AB; B = 16'h0075; #100;
A = 16'h00AB; B = 16'h0076; #100;
A = 16'h00AB; B = 16'h0077; #100;
A = 16'h00AB; B = 16'h0078; #100;
A = 16'h00AB; B = 16'h0079; #100;
A = 16'h00AB; B = 16'h007A; #100;
A = 16'h00AB; B = 16'h007B; #100;
A = 16'h00AB; B = 16'h007C; #100;
A = 16'h00AB; B = 16'h007D; #100;
A = 16'h00AB; B = 16'h007E; #100;
A = 16'h00AB; B = 16'h007F; #100;
A = 16'h00AB; B = 16'h0080; #100;
A = 16'h00AB; B = 16'h0081; #100;
A = 16'h00AB; B = 16'h0082; #100;
A = 16'h00AB; B = 16'h0083; #100;
A = 16'h00AB; B = 16'h0084; #100;
A = 16'h00AB; B = 16'h0085; #100;
A = 16'h00AB; B = 16'h0086; #100;
A = 16'h00AB; B = 16'h0087; #100;
A = 16'h00AB; B = 16'h0088; #100;
A = 16'h00AB; B = 16'h0089; #100;
A = 16'h00AB; B = 16'h008A; #100;
A = 16'h00AB; B = 16'h008B; #100;
A = 16'h00AB; B = 16'h008C; #100;
A = 16'h00AB; B = 16'h008D; #100;
A = 16'h00AB; B = 16'h008E; #100;
A = 16'h00AB; B = 16'h008F; #100;
A = 16'h00AB; B = 16'h0090; #100;
A = 16'h00AB; B = 16'h0091; #100;
A = 16'h00AB; B = 16'h0092; #100;
A = 16'h00AB; B = 16'h0093; #100;
A = 16'h00AB; B = 16'h0094; #100;
A = 16'h00AB; B = 16'h0095; #100;
A = 16'h00AB; B = 16'h0096; #100;
A = 16'h00AB; B = 16'h0097; #100;
A = 16'h00AB; B = 16'h0098; #100;
A = 16'h00AB; B = 16'h0099; #100;
A = 16'h00AB; B = 16'h009A; #100;
A = 16'h00AB; B = 16'h009B; #100;
A = 16'h00AB; B = 16'h009C; #100;
A = 16'h00AB; B = 16'h009D; #100;
A = 16'h00AB; B = 16'h009E; #100;
A = 16'h00AB; B = 16'h009F; #100;
A = 16'h00AB; B = 16'h00A0; #100;
A = 16'h00AB; B = 16'h00A1; #100;
A = 16'h00AB; B = 16'h00A2; #100;
A = 16'h00AB; B = 16'h00A3; #100;
A = 16'h00AB; B = 16'h00A4; #100;
A = 16'h00AB; B = 16'h00A5; #100;
A = 16'h00AB; B = 16'h00A6; #100;
A = 16'h00AB; B = 16'h00A7; #100;
A = 16'h00AB; B = 16'h00A8; #100;
A = 16'h00AB; B = 16'h00A9; #100;
A = 16'h00AB; B = 16'h00AA; #100;
A = 16'h00AB; B = 16'h00AB; #100;
A = 16'h00AB; B = 16'h00AC; #100;
A = 16'h00AB; B = 16'h00AD; #100;
A = 16'h00AB; B = 16'h00AE; #100;
A = 16'h00AB; B = 16'h00AF; #100;
A = 16'h00AB; B = 16'h00B0; #100;
A = 16'h00AB; B = 16'h00B1; #100;
A = 16'h00AB; B = 16'h00B2; #100;
A = 16'h00AB; B = 16'h00B3; #100;
A = 16'h00AB; B = 16'h00B4; #100;
A = 16'h00AB; B = 16'h00B5; #100;
A = 16'h00AB; B = 16'h00B6; #100;
A = 16'h00AB; B = 16'h00B7; #100;
A = 16'h00AB; B = 16'h00B8; #100;
A = 16'h00AB; B = 16'h00B9; #100;
A = 16'h00AB; B = 16'h00BA; #100;
A = 16'h00AB; B = 16'h00BB; #100;
A = 16'h00AB; B = 16'h00BC; #100;
A = 16'h00AB; B = 16'h00BD; #100;
A = 16'h00AB; B = 16'h00BE; #100;
A = 16'h00AB; B = 16'h00BF; #100;
A = 16'h00AB; B = 16'h00C0; #100;
A = 16'h00AB; B = 16'h00C1; #100;
A = 16'h00AB; B = 16'h00C2; #100;
A = 16'h00AB; B = 16'h00C3; #100;
A = 16'h00AB; B = 16'h00C4; #100;
A = 16'h00AB; B = 16'h00C5; #100;
A = 16'h00AB; B = 16'h00C6; #100;
A = 16'h00AB; B = 16'h00C7; #100;
A = 16'h00AB; B = 16'h00C8; #100;
A = 16'h00AB; B = 16'h00C9; #100;
A = 16'h00AB; B = 16'h00CA; #100;
A = 16'h00AB; B = 16'h00CB; #100;
A = 16'h00AB; B = 16'h00CC; #100;
A = 16'h00AB; B = 16'h00CD; #100;
A = 16'h00AB; B = 16'h00CE; #100;
A = 16'h00AB; B = 16'h00CF; #100;
A = 16'h00AB; B = 16'h00D0; #100;
A = 16'h00AB; B = 16'h00D1; #100;
A = 16'h00AB; B = 16'h00D2; #100;
A = 16'h00AB; B = 16'h00D3; #100;
A = 16'h00AB; B = 16'h00D4; #100;
A = 16'h00AB; B = 16'h00D5; #100;
A = 16'h00AB; B = 16'h00D6; #100;
A = 16'h00AB; B = 16'h00D7; #100;
A = 16'h00AB; B = 16'h00D8; #100;
A = 16'h00AB; B = 16'h00D9; #100;
A = 16'h00AB; B = 16'h00DA; #100;
A = 16'h00AB; B = 16'h00DB; #100;
A = 16'h00AB; B = 16'h00DC; #100;
A = 16'h00AB; B = 16'h00DD; #100;
A = 16'h00AB; B = 16'h00DE; #100;
A = 16'h00AB; B = 16'h00DF; #100;
A = 16'h00AB; B = 16'h00E0; #100;
A = 16'h00AB; B = 16'h00E1; #100;
A = 16'h00AB; B = 16'h00E2; #100;
A = 16'h00AB; B = 16'h00E3; #100;
A = 16'h00AB; B = 16'h00E4; #100;
A = 16'h00AB; B = 16'h00E5; #100;
A = 16'h00AB; B = 16'h00E6; #100;
A = 16'h00AB; B = 16'h00E7; #100;
A = 16'h00AB; B = 16'h00E8; #100;
A = 16'h00AB; B = 16'h00E9; #100;
A = 16'h00AB; B = 16'h00EA; #100;
A = 16'h00AB; B = 16'h00EB; #100;
A = 16'h00AB; B = 16'h00EC; #100;
A = 16'h00AB; B = 16'h00ED; #100;
A = 16'h00AB; B = 16'h00EE; #100;
A = 16'h00AB; B = 16'h00EF; #100;
A = 16'h00AB; B = 16'h00F0; #100;
A = 16'h00AB; B = 16'h00F1; #100;
A = 16'h00AB; B = 16'h00F2; #100;
A = 16'h00AB; B = 16'h00F3; #100;
A = 16'h00AB; B = 16'h00F4; #100;
A = 16'h00AB; B = 16'h00F5; #100;
A = 16'h00AB; B = 16'h00F6; #100;
A = 16'h00AB; B = 16'h00F7; #100;
A = 16'h00AB; B = 16'h00F8; #100;
A = 16'h00AB; B = 16'h00F9; #100;
A = 16'h00AB; B = 16'h00FA; #100;
A = 16'h00AB; B = 16'h00FB; #100;
A = 16'h00AB; B = 16'h00FC; #100;
A = 16'h00AB; B = 16'h00FD; #100;
A = 16'h00AB; B = 16'h00FE; #100;
A = 16'h00AB; B = 16'h00FF; #100;
A = 16'h00AC; B = 16'h000; #100;
A = 16'h00AC; B = 16'h001; #100;
A = 16'h00AC; B = 16'h002; #100;
A = 16'h00AC; B = 16'h003; #100;
A = 16'h00AC; B = 16'h004; #100;
A = 16'h00AC; B = 16'h005; #100;
A = 16'h00AC; B = 16'h006; #100;
A = 16'h00AC; B = 16'h007; #100;
A = 16'h00AC; B = 16'h008; #100;
A = 16'h00AC; B = 16'h009; #100;
A = 16'h00AC; B = 16'h00A; #100;
A = 16'h00AC; B = 16'h00B; #100;
A = 16'h00AC; B = 16'h00C; #100;
A = 16'h00AC; B = 16'h00D; #100;
A = 16'h00AC; B = 16'h00E; #100;
A = 16'h00AC; B = 16'h00F; #100;
A = 16'h00AC; B = 16'h0010; #100;
A = 16'h00AC; B = 16'h0011; #100;
A = 16'h00AC; B = 16'h0012; #100;
A = 16'h00AC; B = 16'h0013; #100;
A = 16'h00AC; B = 16'h0014; #100;
A = 16'h00AC; B = 16'h0015; #100;
A = 16'h00AC; B = 16'h0016; #100;
A = 16'h00AC; B = 16'h0017; #100;
A = 16'h00AC; B = 16'h0018; #100;
A = 16'h00AC; B = 16'h0019; #100;
A = 16'h00AC; B = 16'h001A; #100;
A = 16'h00AC; B = 16'h001B; #100;
A = 16'h00AC; B = 16'h001C; #100;
A = 16'h00AC; B = 16'h001D; #100;
A = 16'h00AC; B = 16'h001E; #100;
A = 16'h00AC; B = 16'h001F; #100;
A = 16'h00AC; B = 16'h0020; #100;
A = 16'h00AC; B = 16'h0021; #100;
A = 16'h00AC; B = 16'h0022; #100;
A = 16'h00AC; B = 16'h0023; #100;
A = 16'h00AC; B = 16'h0024; #100;
A = 16'h00AC; B = 16'h0025; #100;
A = 16'h00AC; B = 16'h0026; #100;
A = 16'h00AC; B = 16'h0027; #100;
A = 16'h00AC; B = 16'h0028; #100;
A = 16'h00AC; B = 16'h0029; #100;
A = 16'h00AC; B = 16'h002A; #100;
A = 16'h00AC; B = 16'h002B; #100;
A = 16'h00AC; B = 16'h002C; #100;
A = 16'h00AC; B = 16'h002D; #100;
A = 16'h00AC; B = 16'h002E; #100;
A = 16'h00AC; B = 16'h002F; #100;
A = 16'h00AC; B = 16'h0030; #100;
A = 16'h00AC; B = 16'h0031; #100;
A = 16'h00AC; B = 16'h0032; #100;
A = 16'h00AC; B = 16'h0033; #100;
A = 16'h00AC; B = 16'h0034; #100;
A = 16'h00AC; B = 16'h0035; #100;
A = 16'h00AC; B = 16'h0036; #100;
A = 16'h00AC; B = 16'h0037; #100;
A = 16'h00AC; B = 16'h0038; #100;
A = 16'h00AC; B = 16'h0039; #100;
A = 16'h00AC; B = 16'h003A; #100;
A = 16'h00AC; B = 16'h003B; #100;
A = 16'h00AC; B = 16'h003C; #100;
A = 16'h00AC; B = 16'h003D; #100;
A = 16'h00AC; B = 16'h003E; #100;
A = 16'h00AC; B = 16'h003F; #100;
A = 16'h00AC; B = 16'h0040; #100;
A = 16'h00AC; B = 16'h0041; #100;
A = 16'h00AC; B = 16'h0042; #100;
A = 16'h00AC; B = 16'h0043; #100;
A = 16'h00AC; B = 16'h0044; #100;
A = 16'h00AC; B = 16'h0045; #100;
A = 16'h00AC; B = 16'h0046; #100;
A = 16'h00AC; B = 16'h0047; #100;
A = 16'h00AC; B = 16'h0048; #100;
A = 16'h00AC; B = 16'h0049; #100;
A = 16'h00AC; B = 16'h004A; #100;
A = 16'h00AC; B = 16'h004B; #100;
A = 16'h00AC; B = 16'h004C; #100;
A = 16'h00AC; B = 16'h004D; #100;
A = 16'h00AC; B = 16'h004E; #100;
A = 16'h00AC; B = 16'h004F; #100;
A = 16'h00AC; B = 16'h0050; #100;
A = 16'h00AC; B = 16'h0051; #100;
A = 16'h00AC; B = 16'h0052; #100;
A = 16'h00AC; B = 16'h0053; #100;
A = 16'h00AC; B = 16'h0054; #100;
A = 16'h00AC; B = 16'h0055; #100;
A = 16'h00AC; B = 16'h0056; #100;
A = 16'h00AC; B = 16'h0057; #100;
A = 16'h00AC; B = 16'h0058; #100;
A = 16'h00AC; B = 16'h0059; #100;
A = 16'h00AC; B = 16'h005A; #100;
A = 16'h00AC; B = 16'h005B; #100;
A = 16'h00AC; B = 16'h005C; #100;
A = 16'h00AC; B = 16'h005D; #100;
A = 16'h00AC; B = 16'h005E; #100;
A = 16'h00AC; B = 16'h005F; #100;
A = 16'h00AC; B = 16'h0060; #100;
A = 16'h00AC; B = 16'h0061; #100;
A = 16'h00AC; B = 16'h0062; #100;
A = 16'h00AC; B = 16'h0063; #100;
A = 16'h00AC; B = 16'h0064; #100;
A = 16'h00AC; B = 16'h0065; #100;
A = 16'h00AC; B = 16'h0066; #100;
A = 16'h00AC; B = 16'h0067; #100;
A = 16'h00AC; B = 16'h0068; #100;
A = 16'h00AC; B = 16'h0069; #100;
A = 16'h00AC; B = 16'h006A; #100;
A = 16'h00AC; B = 16'h006B; #100;
A = 16'h00AC; B = 16'h006C; #100;
A = 16'h00AC; B = 16'h006D; #100;
A = 16'h00AC; B = 16'h006E; #100;
A = 16'h00AC; B = 16'h006F; #100;
A = 16'h00AC; B = 16'h0070; #100;
A = 16'h00AC; B = 16'h0071; #100;
A = 16'h00AC; B = 16'h0072; #100;
A = 16'h00AC; B = 16'h0073; #100;
A = 16'h00AC; B = 16'h0074; #100;
A = 16'h00AC; B = 16'h0075; #100;
A = 16'h00AC; B = 16'h0076; #100;
A = 16'h00AC; B = 16'h0077; #100;
A = 16'h00AC; B = 16'h0078; #100;
A = 16'h00AC; B = 16'h0079; #100;
A = 16'h00AC; B = 16'h007A; #100;
A = 16'h00AC; B = 16'h007B; #100;
A = 16'h00AC; B = 16'h007C; #100;
A = 16'h00AC; B = 16'h007D; #100;
A = 16'h00AC; B = 16'h007E; #100;
A = 16'h00AC; B = 16'h007F; #100;
A = 16'h00AC; B = 16'h0080; #100;
A = 16'h00AC; B = 16'h0081; #100;
A = 16'h00AC; B = 16'h0082; #100;
A = 16'h00AC; B = 16'h0083; #100;
A = 16'h00AC; B = 16'h0084; #100;
A = 16'h00AC; B = 16'h0085; #100;
A = 16'h00AC; B = 16'h0086; #100;
A = 16'h00AC; B = 16'h0087; #100;
A = 16'h00AC; B = 16'h0088; #100;
A = 16'h00AC; B = 16'h0089; #100;
A = 16'h00AC; B = 16'h008A; #100;
A = 16'h00AC; B = 16'h008B; #100;
A = 16'h00AC; B = 16'h008C; #100;
A = 16'h00AC; B = 16'h008D; #100;
A = 16'h00AC; B = 16'h008E; #100;
A = 16'h00AC; B = 16'h008F; #100;
A = 16'h00AC; B = 16'h0090; #100;
A = 16'h00AC; B = 16'h0091; #100;
A = 16'h00AC; B = 16'h0092; #100;
A = 16'h00AC; B = 16'h0093; #100;
A = 16'h00AC; B = 16'h0094; #100;
A = 16'h00AC; B = 16'h0095; #100;
A = 16'h00AC; B = 16'h0096; #100;
A = 16'h00AC; B = 16'h0097; #100;
A = 16'h00AC; B = 16'h0098; #100;
A = 16'h00AC; B = 16'h0099; #100;
A = 16'h00AC; B = 16'h009A; #100;
A = 16'h00AC; B = 16'h009B; #100;
A = 16'h00AC; B = 16'h009C; #100;
A = 16'h00AC; B = 16'h009D; #100;
A = 16'h00AC; B = 16'h009E; #100;
A = 16'h00AC; B = 16'h009F; #100;
A = 16'h00AC; B = 16'h00A0; #100;
A = 16'h00AC; B = 16'h00A1; #100;
A = 16'h00AC; B = 16'h00A2; #100;
A = 16'h00AC; B = 16'h00A3; #100;
A = 16'h00AC; B = 16'h00A4; #100;
A = 16'h00AC; B = 16'h00A5; #100;
A = 16'h00AC; B = 16'h00A6; #100;
A = 16'h00AC; B = 16'h00A7; #100;
A = 16'h00AC; B = 16'h00A8; #100;
A = 16'h00AC; B = 16'h00A9; #100;
A = 16'h00AC; B = 16'h00AA; #100;
A = 16'h00AC; B = 16'h00AB; #100;
A = 16'h00AC; B = 16'h00AC; #100;
A = 16'h00AC; B = 16'h00AD; #100;
A = 16'h00AC; B = 16'h00AE; #100;
A = 16'h00AC; B = 16'h00AF; #100;
A = 16'h00AC; B = 16'h00B0; #100;
A = 16'h00AC; B = 16'h00B1; #100;
A = 16'h00AC; B = 16'h00B2; #100;
A = 16'h00AC; B = 16'h00B3; #100;
A = 16'h00AC; B = 16'h00B4; #100;
A = 16'h00AC; B = 16'h00B5; #100;
A = 16'h00AC; B = 16'h00B6; #100;
A = 16'h00AC; B = 16'h00B7; #100;
A = 16'h00AC; B = 16'h00B8; #100;
A = 16'h00AC; B = 16'h00B9; #100;
A = 16'h00AC; B = 16'h00BA; #100;
A = 16'h00AC; B = 16'h00BB; #100;
A = 16'h00AC; B = 16'h00BC; #100;
A = 16'h00AC; B = 16'h00BD; #100;
A = 16'h00AC; B = 16'h00BE; #100;
A = 16'h00AC; B = 16'h00BF; #100;
A = 16'h00AC; B = 16'h00C0; #100;
A = 16'h00AC; B = 16'h00C1; #100;
A = 16'h00AC; B = 16'h00C2; #100;
A = 16'h00AC; B = 16'h00C3; #100;
A = 16'h00AC; B = 16'h00C4; #100;
A = 16'h00AC; B = 16'h00C5; #100;
A = 16'h00AC; B = 16'h00C6; #100;
A = 16'h00AC; B = 16'h00C7; #100;
A = 16'h00AC; B = 16'h00C8; #100;
A = 16'h00AC; B = 16'h00C9; #100;
A = 16'h00AC; B = 16'h00CA; #100;
A = 16'h00AC; B = 16'h00CB; #100;
A = 16'h00AC; B = 16'h00CC; #100;
A = 16'h00AC; B = 16'h00CD; #100;
A = 16'h00AC; B = 16'h00CE; #100;
A = 16'h00AC; B = 16'h00CF; #100;
A = 16'h00AC; B = 16'h00D0; #100;
A = 16'h00AC; B = 16'h00D1; #100;
A = 16'h00AC; B = 16'h00D2; #100;
A = 16'h00AC; B = 16'h00D3; #100;
A = 16'h00AC; B = 16'h00D4; #100;
A = 16'h00AC; B = 16'h00D5; #100;
A = 16'h00AC; B = 16'h00D6; #100;
A = 16'h00AC; B = 16'h00D7; #100;
A = 16'h00AC; B = 16'h00D8; #100;
A = 16'h00AC; B = 16'h00D9; #100;
A = 16'h00AC; B = 16'h00DA; #100;
A = 16'h00AC; B = 16'h00DB; #100;
A = 16'h00AC; B = 16'h00DC; #100;
A = 16'h00AC; B = 16'h00DD; #100;
A = 16'h00AC; B = 16'h00DE; #100;
A = 16'h00AC; B = 16'h00DF; #100;
A = 16'h00AC; B = 16'h00E0; #100;
A = 16'h00AC; B = 16'h00E1; #100;
A = 16'h00AC; B = 16'h00E2; #100;
A = 16'h00AC; B = 16'h00E3; #100;
A = 16'h00AC; B = 16'h00E4; #100;
A = 16'h00AC; B = 16'h00E5; #100;
A = 16'h00AC; B = 16'h00E6; #100;
A = 16'h00AC; B = 16'h00E7; #100;
A = 16'h00AC; B = 16'h00E8; #100;
A = 16'h00AC; B = 16'h00E9; #100;
A = 16'h00AC; B = 16'h00EA; #100;
A = 16'h00AC; B = 16'h00EB; #100;
A = 16'h00AC; B = 16'h00EC; #100;
A = 16'h00AC; B = 16'h00ED; #100;
A = 16'h00AC; B = 16'h00EE; #100;
A = 16'h00AC; B = 16'h00EF; #100;
A = 16'h00AC; B = 16'h00F0; #100;
A = 16'h00AC; B = 16'h00F1; #100;
A = 16'h00AC; B = 16'h00F2; #100;
A = 16'h00AC; B = 16'h00F3; #100;
A = 16'h00AC; B = 16'h00F4; #100;
A = 16'h00AC; B = 16'h00F5; #100;
A = 16'h00AC; B = 16'h00F6; #100;
A = 16'h00AC; B = 16'h00F7; #100;
A = 16'h00AC; B = 16'h00F8; #100;
A = 16'h00AC; B = 16'h00F9; #100;
A = 16'h00AC; B = 16'h00FA; #100;
A = 16'h00AC; B = 16'h00FB; #100;
A = 16'h00AC; B = 16'h00FC; #100;
A = 16'h00AC; B = 16'h00FD; #100;
A = 16'h00AC; B = 16'h00FE; #100;
A = 16'h00AC; B = 16'h00FF; #100;
A = 16'h00AD; B = 16'h000; #100;
A = 16'h00AD; B = 16'h001; #100;
A = 16'h00AD; B = 16'h002; #100;
A = 16'h00AD; B = 16'h003; #100;
A = 16'h00AD; B = 16'h004; #100;
A = 16'h00AD; B = 16'h005; #100;
A = 16'h00AD; B = 16'h006; #100;
A = 16'h00AD; B = 16'h007; #100;
A = 16'h00AD; B = 16'h008; #100;
A = 16'h00AD; B = 16'h009; #100;
A = 16'h00AD; B = 16'h00A; #100;
A = 16'h00AD; B = 16'h00B; #100;
A = 16'h00AD; B = 16'h00C; #100;
A = 16'h00AD; B = 16'h00D; #100;
A = 16'h00AD; B = 16'h00E; #100;
A = 16'h00AD; B = 16'h00F; #100;
A = 16'h00AD; B = 16'h0010; #100;
A = 16'h00AD; B = 16'h0011; #100;
A = 16'h00AD; B = 16'h0012; #100;
A = 16'h00AD; B = 16'h0013; #100;
A = 16'h00AD; B = 16'h0014; #100;
A = 16'h00AD; B = 16'h0015; #100;
A = 16'h00AD; B = 16'h0016; #100;
A = 16'h00AD; B = 16'h0017; #100;
A = 16'h00AD; B = 16'h0018; #100;
A = 16'h00AD; B = 16'h0019; #100;
A = 16'h00AD; B = 16'h001A; #100;
A = 16'h00AD; B = 16'h001B; #100;
A = 16'h00AD; B = 16'h001C; #100;
A = 16'h00AD; B = 16'h001D; #100;
A = 16'h00AD; B = 16'h001E; #100;
A = 16'h00AD; B = 16'h001F; #100;
A = 16'h00AD; B = 16'h0020; #100;
A = 16'h00AD; B = 16'h0021; #100;
A = 16'h00AD; B = 16'h0022; #100;
A = 16'h00AD; B = 16'h0023; #100;
A = 16'h00AD; B = 16'h0024; #100;
A = 16'h00AD; B = 16'h0025; #100;
A = 16'h00AD; B = 16'h0026; #100;
A = 16'h00AD; B = 16'h0027; #100;
A = 16'h00AD; B = 16'h0028; #100;
A = 16'h00AD; B = 16'h0029; #100;
A = 16'h00AD; B = 16'h002A; #100;
A = 16'h00AD; B = 16'h002B; #100;
A = 16'h00AD; B = 16'h002C; #100;
A = 16'h00AD; B = 16'h002D; #100;
A = 16'h00AD; B = 16'h002E; #100;
A = 16'h00AD; B = 16'h002F; #100;
A = 16'h00AD; B = 16'h0030; #100;
A = 16'h00AD; B = 16'h0031; #100;
A = 16'h00AD; B = 16'h0032; #100;
A = 16'h00AD; B = 16'h0033; #100;
A = 16'h00AD; B = 16'h0034; #100;
A = 16'h00AD; B = 16'h0035; #100;
A = 16'h00AD; B = 16'h0036; #100;
A = 16'h00AD; B = 16'h0037; #100;
A = 16'h00AD; B = 16'h0038; #100;
A = 16'h00AD; B = 16'h0039; #100;
A = 16'h00AD; B = 16'h003A; #100;
A = 16'h00AD; B = 16'h003B; #100;
A = 16'h00AD; B = 16'h003C; #100;
A = 16'h00AD; B = 16'h003D; #100;
A = 16'h00AD; B = 16'h003E; #100;
A = 16'h00AD; B = 16'h003F; #100;
A = 16'h00AD; B = 16'h0040; #100;
A = 16'h00AD; B = 16'h0041; #100;
A = 16'h00AD; B = 16'h0042; #100;
A = 16'h00AD; B = 16'h0043; #100;
A = 16'h00AD; B = 16'h0044; #100;
A = 16'h00AD; B = 16'h0045; #100;
A = 16'h00AD; B = 16'h0046; #100;
A = 16'h00AD; B = 16'h0047; #100;
A = 16'h00AD; B = 16'h0048; #100;
A = 16'h00AD; B = 16'h0049; #100;
A = 16'h00AD; B = 16'h004A; #100;
A = 16'h00AD; B = 16'h004B; #100;
A = 16'h00AD; B = 16'h004C; #100;
A = 16'h00AD; B = 16'h004D; #100;
A = 16'h00AD; B = 16'h004E; #100;
A = 16'h00AD; B = 16'h004F; #100;
A = 16'h00AD; B = 16'h0050; #100;
A = 16'h00AD; B = 16'h0051; #100;
A = 16'h00AD; B = 16'h0052; #100;
A = 16'h00AD; B = 16'h0053; #100;
A = 16'h00AD; B = 16'h0054; #100;
A = 16'h00AD; B = 16'h0055; #100;
A = 16'h00AD; B = 16'h0056; #100;
A = 16'h00AD; B = 16'h0057; #100;
A = 16'h00AD; B = 16'h0058; #100;
A = 16'h00AD; B = 16'h0059; #100;
A = 16'h00AD; B = 16'h005A; #100;
A = 16'h00AD; B = 16'h005B; #100;
A = 16'h00AD; B = 16'h005C; #100;
A = 16'h00AD; B = 16'h005D; #100;
A = 16'h00AD; B = 16'h005E; #100;
A = 16'h00AD; B = 16'h005F; #100;
A = 16'h00AD; B = 16'h0060; #100;
A = 16'h00AD; B = 16'h0061; #100;
A = 16'h00AD; B = 16'h0062; #100;
A = 16'h00AD; B = 16'h0063; #100;
A = 16'h00AD; B = 16'h0064; #100;
A = 16'h00AD; B = 16'h0065; #100;
A = 16'h00AD; B = 16'h0066; #100;
A = 16'h00AD; B = 16'h0067; #100;
A = 16'h00AD; B = 16'h0068; #100;
A = 16'h00AD; B = 16'h0069; #100;
A = 16'h00AD; B = 16'h006A; #100;
A = 16'h00AD; B = 16'h006B; #100;
A = 16'h00AD; B = 16'h006C; #100;
A = 16'h00AD; B = 16'h006D; #100;
A = 16'h00AD; B = 16'h006E; #100;
A = 16'h00AD; B = 16'h006F; #100;
A = 16'h00AD; B = 16'h0070; #100;
A = 16'h00AD; B = 16'h0071; #100;
A = 16'h00AD; B = 16'h0072; #100;
A = 16'h00AD; B = 16'h0073; #100;
A = 16'h00AD; B = 16'h0074; #100;
A = 16'h00AD; B = 16'h0075; #100;
A = 16'h00AD; B = 16'h0076; #100;
A = 16'h00AD; B = 16'h0077; #100;
A = 16'h00AD; B = 16'h0078; #100;
A = 16'h00AD; B = 16'h0079; #100;
A = 16'h00AD; B = 16'h007A; #100;
A = 16'h00AD; B = 16'h007B; #100;
A = 16'h00AD; B = 16'h007C; #100;
A = 16'h00AD; B = 16'h007D; #100;
A = 16'h00AD; B = 16'h007E; #100;
A = 16'h00AD; B = 16'h007F; #100;
A = 16'h00AD; B = 16'h0080; #100;
A = 16'h00AD; B = 16'h0081; #100;
A = 16'h00AD; B = 16'h0082; #100;
A = 16'h00AD; B = 16'h0083; #100;
A = 16'h00AD; B = 16'h0084; #100;
A = 16'h00AD; B = 16'h0085; #100;
A = 16'h00AD; B = 16'h0086; #100;
A = 16'h00AD; B = 16'h0087; #100;
A = 16'h00AD; B = 16'h0088; #100;
A = 16'h00AD; B = 16'h0089; #100;
A = 16'h00AD; B = 16'h008A; #100;
A = 16'h00AD; B = 16'h008B; #100;
A = 16'h00AD; B = 16'h008C; #100;
A = 16'h00AD; B = 16'h008D; #100;
A = 16'h00AD; B = 16'h008E; #100;
A = 16'h00AD; B = 16'h008F; #100;
A = 16'h00AD; B = 16'h0090; #100;
A = 16'h00AD; B = 16'h0091; #100;
A = 16'h00AD; B = 16'h0092; #100;
A = 16'h00AD; B = 16'h0093; #100;
A = 16'h00AD; B = 16'h0094; #100;
A = 16'h00AD; B = 16'h0095; #100;
A = 16'h00AD; B = 16'h0096; #100;
A = 16'h00AD; B = 16'h0097; #100;
A = 16'h00AD; B = 16'h0098; #100;
A = 16'h00AD; B = 16'h0099; #100;
A = 16'h00AD; B = 16'h009A; #100;
A = 16'h00AD; B = 16'h009B; #100;
A = 16'h00AD; B = 16'h009C; #100;
A = 16'h00AD; B = 16'h009D; #100;
A = 16'h00AD; B = 16'h009E; #100;
A = 16'h00AD; B = 16'h009F; #100;
A = 16'h00AD; B = 16'h00A0; #100;
A = 16'h00AD; B = 16'h00A1; #100;
A = 16'h00AD; B = 16'h00A2; #100;
A = 16'h00AD; B = 16'h00A3; #100;
A = 16'h00AD; B = 16'h00A4; #100;
A = 16'h00AD; B = 16'h00A5; #100;
A = 16'h00AD; B = 16'h00A6; #100;
A = 16'h00AD; B = 16'h00A7; #100;
A = 16'h00AD; B = 16'h00A8; #100;
A = 16'h00AD; B = 16'h00A9; #100;
A = 16'h00AD; B = 16'h00AA; #100;
A = 16'h00AD; B = 16'h00AB; #100;
A = 16'h00AD; B = 16'h00AC; #100;
A = 16'h00AD; B = 16'h00AD; #100;
A = 16'h00AD; B = 16'h00AE; #100;
A = 16'h00AD; B = 16'h00AF; #100;
A = 16'h00AD; B = 16'h00B0; #100;
A = 16'h00AD; B = 16'h00B1; #100;
A = 16'h00AD; B = 16'h00B2; #100;
A = 16'h00AD; B = 16'h00B3; #100;
A = 16'h00AD; B = 16'h00B4; #100;
A = 16'h00AD; B = 16'h00B5; #100;
A = 16'h00AD; B = 16'h00B6; #100;
A = 16'h00AD; B = 16'h00B7; #100;
A = 16'h00AD; B = 16'h00B8; #100;
A = 16'h00AD; B = 16'h00B9; #100;
A = 16'h00AD; B = 16'h00BA; #100;
A = 16'h00AD; B = 16'h00BB; #100;
A = 16'h00AD; B = 16'h00BC; #100;
A = 16'h00AD; B = 16'h00BD; #100;
A = 16'h00AD; B = 16'h00BE; #100;
A = 16'h00AD; B = 16'h00BF; #100;
A = 16'h00AD; B = 16'h00C0; #100;
A = 16'h00AD; B = 16'h00C1; #100;
A = 16'h00AD; B = 16'h00C2; #100;
A = 16'h00AD; B = 16'h00C3; #100;
A = 16'h00AD; B = 16'h00C4; #100;
A = 16'h00AD; B = 16'h00C5; #100;
A = 16'h00AD; B = 16'h00C6; #100;
A = 16'h00AD; B = 16'h00C7; #100;
A = 16'h00AD; B = 16'h00C8; #100;
A = 16'h00AD; B = 16'h00C9; #100;
A = 16'h00AD; B = 16'h00CA; #100;
A = 16'h00AD; B = 16'h00CB; #100;
A = 16'h00AD; B = 16'h00CC; #100;
A = 16'h00AD; B = 16'h00CD; #100;
A = 16'h00AD; B = 16'h00CE; #100;
A = 16'h00AD; B = 16'h00CF; #100;
A = 16'h00AD; B = 16'h00D0; #100;
A = 16'h00AD; B = 16'h00D1; #100;
A = 16'h00AD; B = 16'h00D2; #100;
A = 16'h00AD; B = 16'h00D3; #100;
A = 16'h00AD; B = 16'h00D4; #100;
A = 16'h00AD; B = 16'h00D5; #100;
A = 16'h00AD; B = 16'h00D6; #100;
A = 16'h00AD; B = 16'h00D7; #100;
A = 16'h00AD; B = 16'h00D8; #100;
A = 16'h00AD; B = 16'h00D9; #100;
A = 16'h00AD; B = 16'h00DA; #100;
A = 16'h00AD; B = 16'h00DB; #100;
A = 16'h00AD; B = 16'h00DC; #100;
A = 16'h00AD; B = 16'h00DD; #100;
A = 16'h00AD; B = 16'h00DE; #100;
A = 16'h00AD; B = 16'h00DF; #100;
A = 16'h00AD; B = 16'h00E0; #100;
A = 16'h00AD; B = 16'h00E1; #100;
A = 16'h00AD; B = 16'h00E2; #100;
A = 16'h00AD; B = 16'h00E3; #100;
A = 16'h00AD; B = 16'h00E4; #100;
A = 16'h00AD; B = 16'h00E5; #100;
A = 16'h00AD; B = 16'h00E6; #100;
A = 16'h00AD; B = 16'h00E7; #100;
A = 16'h00AD; B = 16'h00E8; #100;
A = 16'h00AD; B = 16'h00E9; #100;
A = 16'h00AD; B = 16'h00EA; #100;
A = 16'h00AD; B = 16'h00EB; #100;
A = 16'h00AD; B = 16'h00EC; #100;
A = 16'h00AD; B = 16'h00ED; #100;
A = 16'h00AD; B = 16'h00EE; #100;
A = 16'h00AD; B = 16'h00EF; #100;
A = 16'h00AD; B = 16'h00F0; #100;
A = 16'h00AD; B = 16'h00F1; #100;
A = 16'h00AD; B = 16'h00F2; #100;
A = 16'h00AD; B = 16'h00F3; #100;
A = 16'h00AD; B = 16'h00F4; #100;
A = 16'h00AD; B = 16'h00F5; #100;
A = 16'h00AD; B = 16'h00F6; #100;
A = 16'h00AD; B = 16'h00F7; #100;
A = 16'h00AD; B = 16'h00F8; #100;
A = 16'h00AD; B = 16'h00F9; #100;
A = 16'h00AD; B = 16'h00FA; #100;
A = 16'h00AD; B = 16'h00FB; #100;
A = 16'h00AD; B = 16'h00FC; #100;
A = 16'h00AD; B = 16'h00FD; #100;
A = 16'h00AD; B = 16'h00FE; #100;
A = 16'h00AD; B = 16'h00FF; #100;
A = 16'h00AE; B = 16'h000; #100;
A = 16'h00AE; B = 16'h001; #100;
A = 16'h00AE; B = 16'h002; #100;
A = 16'h00AE; B = 16'h003; #100;
A = 16'h00AE; B = 16'h004; #100;
A = 16'h00AE; B = 16'h005; #100;
A = 16'h00AE; B = 16'h006; #100;
A = 16'h00AE; B = 16'h007; #100;
A = 16'h00AE; B = 16'h008; #100;
A = 16'h00AE; B = 16'h009; #100;
A = 16'h00AE; B = 16'h00A; #100;
A = 16'h00AE; B = 16'h00B; #100;
A = 16'h00AE; B = 16'h00C; #100;
A = 16'h00AE; B = 16'h00D; #100;
A = 16'h00AE; B = 16'h00E; #100;
A = 16'h00AE; B = 16'h00F; #100;
A = 16'h00AE; B = 16'h0010; #100;
A = 16'h00AE; B = 16'h0011; #100;
A = 16'h00AE; B = 16'h0012; #100;
A = 16'h00AE; B = 16'h0013; #100;
A = 16'h00AE; B = 16'h0014; #100;
A = 16'h00AE; B = 16'h0015; #100;
A = 16'h00AE; B = 16'h0016; #100;
A = 16'h00AE; B = 16'h0017; #100;
A = 16'h00AE; B = 16'h0018; #100;
A = 16'h00AE; B = 16'h0019; #100;
A = 16'h00AE; B = 16'h001A; #100;
A = 16'h00AE; B = 16'h001B; #100;
A = 16'h00AE; B = 16'h001C; #100;
A = 16'h00AE; B = 16'h001D; #100;
A = 16'h00AE; B = 16'h001E; #100;
A = 16'h00AE; B = 16'h001F; #100;
A = 16'h00AE; B = 16'h0020; #100;
A = 16'h00AE; B = 16'h0021; #100;
A = 16'h00AE; B = 16'h0022; #100;
A = 16'h00AE; B = 16'h0023; #100;
A = 16'h00AE; B = 16'h0024; #100;
A = 16'h00AE; B = 16'h0025; #100;
A = 16'h00AE; B = 16'h0026; #100;
A = 16'h00AE; B = 16'h0027; #100;
A = 16'h00AE; B = 16'h0028; #100;
A = 16'h00AE; B = 16'h0029; #100;
A = 16'h00AE; B = 16'h002A; #100;
A = 16'h00AE; B = 16'h002B; #100;
A = 16'h00AE; B = 16'h002C; #100;
A = 16'h00AE; B = 16'h002D; #100;
A = 16'h00AE; B = 16'h002E; #100;
A = 16'h00AE; B = 16'h002F; #100;
A = 16'h00AE; B = 16'h0030; #100;
A = 16'h00AE; B = 16'h0031; #100;
A = 16'h00AE; B = 16'h0032; #100;
A = 16'h00AE; B = 16'h0033; #100;
A = 16'h00AE; B = 16'h0034; #100;
A = 16'h00AE; B = 16'h0035; #100;
A = 16'h00AE; B = 16'h0036; #100;
A = 16'h00AE; B = 16'h0037; #100;
A = 16'h00AE; B = 16'h0038; #100;
A = 16'h00AE; B = 16'h0039; #100;
A = 16'h00AE; B = 16'h003A; #100;
A = 16'h00AE; B = 16'h003B; #100;
A = 16'h00AE; B = 16'h003C; #100;
A = 16'h00AE; B = 16'h003D; #100;
A = 16'h00AE; B = 16'h003E; #100;
A = 16'h00AE; B = 16'h003F; #100;
A = 16'h00AE; B = 16'h0040; #100;
A = 16'h00AE; B = 16'h0041; #100;
A = 16'h00AE; B = 16'h0042; #100;
A = 16'h00AE; B = 16'h0043; #100;
A = 16'h00AE; B = 16'h0044; #100;
A = 16'h00AE; B = 16'h0045; #100;
A = 16'h00AE; B = 16'h0046; #100;
A = 16'h00AE; B = 16'h0047; #100;
A = 16'h00AE; B = 16'h0048; #100;
A = 16'h00AE; B = 16'h0049; #100;
A = 16'h00AE; B = 16'h004A; #100;
A = 16'h00AE; B = 16'h004B; #100;
A = 16'h00AE; B = 16'h004C; #100;
A = 16'h00AE; B = 16'h004D; #100;
A = 16'h00AE; B = 16'h004E; #100;
A = 16'h00AE; B = 16'h004F; #100;
A = 16'h00AE; B = 16'h0050; #100;
A = 16'h00AE; B = 16'h0051; #100;
A = 16'h00AE; B = 16'h0052; #100;
A = 16'h00AE; B = 16'h0053; #100;
A = 16'h00AE; B = 16'h0054; #100;
A = 16'h00AE; B = 16'h0055; #100;
A = 16'h00AE; B = 16'h0056; #100;
A = 16'h00AE; B = 16'h0057; #100;
A = 16'h00AE; B = 16'h0058; #100;
A = 16'h00AE; B = 16'h0059; #100;
A = 16'h00AE; B = 16'h005A; #100;
A = 16'h00AE; B = 16'h005B; #100;
A = 16'h00AE; B = 16'h005C; #100;
A = 16'h00AE; B = 16'h005D; #100;
A = 16'h00AE; B = 16'h005E; #100;
A = 16'h00AE; B = 16'h005F; #100;
A = 16'h00AE; B = 16'h0060; #100;
A = 16'h00AE; B = 16'h0061; #100;
A = 16'h00AE; B = 16'h0062; #100;
A = 16'h00AE; B = 16'h0063; #100;
A = 16'h00AE; B = 16'h0064; #100;
A = 16'h00AE; B = 16'h0065; #100;
A = 16'h00AE; B = 16'h0066; #100;
A = 16'h00AE; B = 16'h0067; #100;
A = 16'h00AE; B = 16'h0068; #100;
A = 16'h00AE; B = 16'h0069; #100;
A = 16'h00AE; B = 16'h006A; #100;
A = 16'h00AE; B = 16'h006B; #100;
A = 16'h00AE; B = 16'h006C; #100;
A = 16'h00AE; B = 16'h006D; #100;
A = 16'h00AE; B = 16'h006E; #100;
A = 16'h00AE; B = 16'h006F; #100;
A = 16'h00AE; B = 16'h0070; #100;
A = 16'h00AE; B = 16'h0071; #100;
A = 16'h00AE; B = 16'h0072; #100;
A = 16'h00AE; B = 16'h0073; #100;
A = 16'h00AE; B = 16'h0074; #100;
A = 16'h00AE; B = 16'h0075; #100;
A = 16'h00AE; B = 16'h0076; #100;
A = 16'h00AE; B = 16'h0077; #100;
A = 16'h00AE; B = 16'h0078; #100;
A = 16'h00AE; B = 16'h0079; #100;
A = 16'h00AE; B = 16'h007A; #100;
A = 16'h00AE; B = 16'h007B; #100;
A = 16'h00AE; B = 16'h007C; #100;
A = 16'h00AE; B = 16'h007D; #100;
A = 16'h00AE; B = 16'h007E; #100;
A = 16'h00AE; B = 16'h007F; #100;
A = 16'h00AE; B = 16'h0080; #100;
A = 16'h00AE; B = 16'h0081; #100;
A = 16'h00AE; B = 16'h0082; #100;
A = 16'h00AE; B = 16'h0083; #100;
A = 16'h00AE; B = 16'h0084; #100;
A = 16'h00AE; B = 16'h0085; #100;
A = 16'h00AE; B = 16'h0086; #100;
A = 16'h00AE; B = 16'h0087; #100;
A = 16'h00AE; B = 16'h0088; #100;
A = 16'h00AE; B = 16'h0089; #100;
A = 16'h00AE; B = 16'h008A; #100;
A = 16'h00AE; B = 16'h008B; #100;
A = 16'h00AE; B = 16'h008C; #100;
A = 16'h00AE; B = 16'h008D; #100;
A = 16'h00AE; B = 16'h008E; #100;
A = 16'h00AE; B = 16'h008F; #100;
A = 16'h00AE; B = 16'h0090; #100;
A = 16'h00AE; B = 16'h0091; #100;
A = 16'h00AE; B = 16'h0092; #100;
A = 16'h00AE; B = 16'h0093; #100;
A = 16'h00AE; B = 16'h0094; #100;
A = 16'h00AE; B = 16'h0095; #100;
A = 16'h00AE; B = 16'h0096; #100;
A = 16'h00AE; B = 16'h0097; #100;
A = 16'h00AE; B = 16'h0098; #100;
A = 16'h00AE; B = 16'h0099; #100;
A = 16'h00AE; B = 16'h009A; #100;
A = 16'h00AE; B = 16'h009B; #100;
A = 16'h00AE; B = 16'h009C; #100;
A = 16'h00AE; B = 16'h009D; #100;
A = 16'h00AE; B = 16'h009E; #100;
A = 16'h00AE; B = 16'h009F; #100;
A = 16'h00AE; B = 16'h00A0; #100;
A = 16'h00AE; B = 16'h00A1; #100;
A = 16'h00AE; B = 16'h00A2; #100;
A = 16'h00AE; B = 16'h00A3; #100;
A = 16'h00AE; B = 16'h00A4; #100;
A = 16'h00AE; B = 16'h00A5; #100;
A = 16'h00AE; B = 16'h00A6; #100;
A = 16'h00AE; B = 16'h00A7; #100;
A = 16'h00AE; B = 16'h00A8; #100;
A = 16'h00AE; B = 16'h00A9; #100;
A = 16'h00AE; B = 16'h00AA; #100;
A = 16'h00AE; B = 16'h00AB; #100;
A = 16'h00AE; B = 16'h00AC; #100;
A = 16'h00AE; B = 16'h00AD; #100;
A = 16'h00AE; B = 16'h00AE; #100;
A = 16'h00AE; B = 16'h00AF; #100;
A = 16'h00AE; B = 16'h00B0; #100;
A = 16'h00AE; B = 16'h00B1; #100;
A = 16'h00AE; B = 16'h00B2; #100;
A = 16'h00AE; B = 16'h00B3; #100;
A = 16'h00AE; B = 16'h00B4; #100;
A = 16'h00AE; B = 16'h00B5; #100;
A = 16'h00AE; B = 16'h00B6; #100;
A = 16'h00AE; B = 16'h00B7; #100;
A = 16'h00AE; B = 16'h00B8; #100;
A = 16'h00AE; B = 16'h00B9; #100;
A = 16'h00AE; B = 16'h00BA; #100;
A = 16'h00AE; B = 16'h00BB; #100;
A = 16'h00AE; B = 16'h00BC; #100;
A = 16'h00AE; B = 16'h00BD; #100;
A = 16'h00AE; B = 16'h00BE; #100;
A = 16'h00AE; B = 16'h00BF; #100;
A = 16'h00AE; B = 16'h00C0; #100;
A = 16'h00AE; B = 16'h00C1; #100;
A = 16'h00AE; B = 16'h00C2; #100;
A = 16'h00AE; B = 16'h00C3; #100;
A = 16'h00AE; B = 16'h00C4; #100;
A = 16'h00AE; B = 16'h00C5; #100;
A = 16'h00AE; B = 16'h00C6; #100;
A = 16'h00AE; B = 16'h00C7; #100;
A = 16'h00AE; B = 16'h00C8; #100;
A = 16'h00AE; B = 16'h00C9; #100;
A = 16'h00AE; B = 16'h00CA; #100;
A = 16'h00AE; B = 16'h00CB; #100;
A = 16'h00AE; B = 16'h00CC; #100;
A = 16'h00AE; B = 16'h00CD; #100;
A = 16'h00AE; B = 16'h00CE; #100;
A = 16'h00AE; B = 16'h00CF; #100;
A = 16'h00AE; B = 16'h00D0; #100;
A = 16'h00AE; B = 16'h00D1; #100;
A = 16'h00AE; B = 16'h00D2; #100;
A = 16'h00AE; B = 16'h00D3; #100;
A = 16'h00AE; B = 16'h00D4; #100;
A = 16'h00AE; B = 16'h00D5; #100;
A = 16'h00AE; B = 16'h00D6; #100;
A = 16'h00AE; B = 16'h00D7; #100;
A = 16'h00AE; B = 16'h00D8; #100;
A = 16'h00AE; B = 16'h00D9; #100;
A = 16'h00AE; B = 16'h00DA; #100;
A = 16'h00AE; B = 16'h00DB; #100;
A = 16'h00AE; B = 16'h00DC; #100;
A = 16'h00AE; B = 16'h00DD; #100;
A = 16'h00AE; B = 16'h00DE; #100;
A = 16'h00AE; B = 16'h00DF; #100;
A = 16'h00AE; B = 16'h00E0; #100;
A = 16'h00AE; B = 16'h00E1; #100;
A = 16'h00AE; B = 16'h00E2; #100;
A = 16'h00AE; B = 16'h00E3; #100;
A = 16'h00AE; B = 16'h00E4; #100;
A = 16'h00AE; B = 16'h00E5; #100;
A = 16'h00AE; B = 16'h00E6; #100;
A = 16'h00AE; B = 16'h00E7; #100;
A = 16'h00AE; B = 16'h00E8; #100;
A = 16'h00AE; B = 16'h00E9; #100;
A = 16'h00AE; B = 16'h00EA; #100;
A = 16'h00AE; B = 16'h00EB; #100;
A = 16'h00AE; B = 16'h00EC; #100;
A = 16'h00AE; B = 16'h00ED; #100;
A = 16'h00AE; B = 16'h00EE; #100;
A = 16'h00AE; B = 16'h00EF; #100;
A = 16'h00AE; B = 16'h00F0; #100;
A = 16'h00AE; B = 16'h00F1; #100;
A = 16'h00AE; B = 16'h00F2; #100;
A = 16'h00AE; B = 16'h00F3; #100;
A = 16'h00AE; B = 16'h00F4; #100;
A = 16'h00AE; B = 16'h00F5; #100;
A = 16'h00AE; B = 16'h00F6; #100;
A = 16'h00AE; B = 16'h00F7; #100;
A = 16'h00AE; B = 16'h00F8; #100;
A = 16'h00AE; B = 16'h00F9; #100;
A = 16'h00AE; B = 16'h00FA; #100;
A = 16'h00AE; B = 16'h00FB; #100;
A = 16'h00AE; B = 16'h00FC; #100;
A = 16'h00AE; B = 16'h00FD; #100;
A = 16'h00AE; B = 16'h00FE; #100;
A = 16'h00AE; B = 16'h00FF; #100;
A = 16'h00AF; B = 16'h000; #100;
A = 16'h00AF; B = 16'h001; #100;
A = 16'h00AF; B = 16'h002; #100;
A = 16'h00AF; B = 16'h003; #100;
A = 16'h00AF; B = 16'h004; #100;
A = 16'h00AF; B = 16'h005; #100;
A = 16'h00AF; B = 16'h006; #100;
A = 16'h00AF; B = 16'h007; #100;
A = 16'h00AF; B = 16'h008; #100;
A = 16'h00AF; B = 16'h009; #100;
A = 16'h00AF; B = 16'h00A; #100;
A = 16'h00AF; B = 16'h00B; #100;
A = 16'h00AF; B = 16'h00C; #100;
A = 16'h00AF; B = 16'h00D; #100;
A = 16'h00AF; B = 16'h00E; #100;
A = 16'h00AF; B = 16'h00F; #100;
A = 16'h00AF; B = 16'h0010; #100;
A = 16'h00AF; B = 16'h0011; #100;
A = 16'h00AF; B = 16'h0012; #100;
A = 16'h00AF; B = 16'h0013; #100;
A = 16'h00AF; B = 16'h0014; #100;
A = 16'h00AF; B = 16'h0015; #100;
A = 16'h00AF; B = 16'h0016; #100;
A = 16'h00AF; B = 16'h0017; #100;
A = 16'h00AF; B = 16'h0018; #100;
A = 16'h00AF; B = 16'h0019; #100;
A = 16'h00AF; B = 16'h001A; #100;
A = 16'h00AF; B = 16'h001B; #100;
A = 16'h00AF; B = 16'h001C; #100;
A = 16'h00AF; B = 16'h001D; #100;
A = 16'h00AF; B = 16'h001E; #100;
A = 16'h00AF; B = 16'h001F; #100;
A = 16'h00AF; B = 16'h0020; #100;
A = 16'h00AF; B = 16'h0021; #100;
A = 16'h00AF; B = 16'h0022; #100;
A = 16'h00AF; B = 16'h0023; #100;
A = 16'h00AF; B = 16'h0024; #100;
A = 16'h00AF; B = 16'h0025; #100;
A = 16'h00AF; B = 16'h0026; #100;
A = 16'h00AF; B = 16'h0027; #100;
A = 16'h00AF; B = 16'h0028; #100;
A = 16'h00AF; B = 16'h0029; #100;
A = 16'h00AF; B = 16'h002A; #100;
A = 16'h00AF; B = 16'h002B; #100;
A = 16'h00AF; B = 16'h002C; #100;
A = 16'h00AF; B = 16'h002D; #100;
A = 16'h00AF; B = 16'h002E; #100;
A = 16'h00AF; B = 16'h002F; #100;
A = 16'h00AF; B = 16'h0030; #100;
A = 16'h00AF; B = 16'h0031; #100;
A = 16'h00AF; B = 16'h0032; #100;
A = 16'h00AF; B = 16'h0033; #100;
A = 16'h00AF; B = 16'h0034; #100;
A = 16'h00AF; B = 16'h0035; #100;
A = 16'h00AF; B = 16'h0036; #100;
A = 16'h00AF; B = 16'h0037; #100;
A = 16'h00AF; B = 16'h0038; #100;
A = 16'h00AF; B = 16'h0039; #100;
A = 16'h00AF; B = 16'h003A; #100;
A = 16'h00AF; B = 16'h003B; #100;
A = 16'h00AF; B = 16'h003C; #100;
A = 16'h00AF; B = 16'h003D; #100;
A = 16'h00AF; B = 16'h003E; #100;
A = 16'h00AF; B = 16'h003F; #100;
A = 16'h00AF; B = 16'h0040; #100;
A = 16'h00AF; B = 16'h0041; #100;
A = 16'h00AF; B = 16'h0042; #100;
A = 16'h00AF; B = 16'h0043; #100;
A = 16'h00AF; B = 16'h0044; #100;
A = 16'h00AF; B = 16'h0045; #100;
A = 16'h00AF; B = 16'h0046; #100;
A = 16'h00AF; B = 16'h0047; #100;
A = 16'h00AF; B = 16'h0048; #100;
A = 16'h00AF; B = 16'h0049; #100;
A = 16'h00AF; B = 16'h004A; #100;
A = 16'h00AF; B = 16'h004B; #100;
A = 16'h00AF; B = 16'h004C; #100;
A = 16'h00AF; B = 16'h004D; #100;
A = 16'h00AF; B = 16'h004E; #100;
A = 16'h00AF; B = 16'h004F; #100;
A = 16'h00AF; B = 16'h0050; #100;
A = 16'h00AF; B = 16'h0051; #100;
A = 16'h00AF; B = 16'h0052; #100;
A = 16'h00AF; B = 16'h0053; #100;
A = 16'h00AF; B = 16'h0054; #100;
A = 16'h00AF; B = 16'h0055; #100;
A = 16'h00AF; B = 16'h0056; #100;
A = 16'h00AF; B = 16'h0057; #100;
A = 16'h00AF; B = 16'h0058; #100;
A = 16'h00AF; B = 16'h0059; #100;
A = 16'h00AF; B = 16'h005A; #100;
A = 16'h00AF; B = 16'h005B; #100;
A = 16'h00AF; B = 16'h005C; #100;
A = 16'h00AF; B = 16'h005D; #100;
A = 16'h00AF; B = 16'h005E; #100;
A = 16'h00AF; B = 16'h005F; #100;
A = 16'h00AF; B = 16'h0060; #100;
A = 16'h00AF; B = 16'h0061; #100;
A = 16'h00AF; B = 16'h0062; #100;
A = 16'h00AF; B = 16'h0063; #100;
A = 16'h00AF; B = 16'h0064; #100;
A = 16'h00AF; B = 16'h0065; #100;
A = 16'h00AF; B = 16'h0066; #100;
A = 16'h00AF; B = 16'h0067; #100;
A = 16'h00AF; B = 16'h0068; #100;
A = 16'h00AF; B = 16'h0069; #100;
A = 16'h00AF; B = 16'h006A; #100;
A = 16'h00AF; B = 16'h006B; #100;
A = 16'h00AF; B = 16'h006C; #100;
A = 16'h00AF; B = 16'h006D; #100;
A = 16'h00AF; B = 16'h006E; #100;
A = 16'h00AF; B = 16'h006F; #100;
A = 16'h00AF; B = 16'h0070; #100;
A = 16'h00AF; B = 16'h0071; #100;
A = 16'h00AF; B = 16'h0072; #100;
A = 16'h00AF; B = 16'h0073; #100;
A = 16'h00AF; B = 16'h0074; #100;
A = 16'h00AF; B = 16'h0075; #100;
A = 16'h00AF; B = 16'h0076; #100;
A = 16'h00AF; B = 16'h0077; #100;
A = 16'h00AF; B = 16'h0078; #100;
A = 16'h00AF; B = 16'h0079; #100;
A = 16'h00AF; B = 16'h007A; #100;
A = 16'h00AF; B = 16'h007B; #100;
A = 16'h00AF; B = 16'h007C; #100;
A = 16'h00AF; B = 16'h007D; #100;
A = 16'h00AF; B = 16'h007E; #100;
A = 16'h00AF; B = 16'h007F; #100;
A = 16'h00AF; B = 16'h0080; #100;
A = 16'h00AF; B = 16'h0081; #100;
A = 16'h00AF; B = 16'h0082; #100;
A = 16'h00AF; B = 16'h0083; #100;
A = 16'h00AF; B = 16'h0084; #100;
A = 16'h00AF; B = 16'h0085; #100;
A = 16'h00AF; B = 16'h0086; #100;
A = 16'h00AF; B = 16'h0087; #100;
A = 16'h00AF; B = 16'h0088; #100;
A = 16'h00AF; B = 16'h0089; #100;
A = 16'h00AF; B = 16'h008A; #100;
A = 16'h00AF; B = 16'h008B; #100;
A = 16'h00AF; B = 16'h008C; #100;
A = 16'h00AF; B = 16'h008D; #100;
A = 16'h00AF; B = 16'h008E; #100;
A = 16'h00AF; B = 16'h008F; #100;
A = 16'h00AF; B = 16'h0090; #100;
A = 16'h00AF; B = 16'h0091; #100;
A = 16'h00AF; B = 16'h0092; #100;
A = 16'h00AF; B = 16'h0093; #100;
A = 16'h00AF; B = 16'h0094; #100;
A = 16'h00AF; B = 16'h0095; #100;
A = 16'h00AF; B = 16'h0096; #100;
A = 16'h00AF; B = 16'h0097; #100;
A = 16'h00AF; B = 16'h0098; #100;
A = 16'h00AF; B = 16'h0099; #100;
A = 16'h00AF; B = 16'h009A; #100;
A = 16'h00AF; B = 16'h009B; #100;
A = 16'h00AF; B = 16'h009C; #100;
A = 16'h00AF; B = 16'h009D; #100;
A = 16'h00AF; B = 16'h009E; #100;
A = 16'h00AF; B = 16'h009F; #100;
A = 16'h00AF; B = 16'h00A0; #100;
A = 16'h00AF; B = 16'h00A1; #100;
A = 16'h00AF; B = 16'h00A2; #100;
A = 16'h00AF; B = 16'h00A3; #100;
A = 16'h00AF; B = 16'h00A4; #100;
A = 16'h00AF; B = 16'h00A5; #100;
A = 16'h00AF; B = 16'h00A6; #100;
A = 16'h00AF; B = 16'h00A7; #100;
A = 16'h00AF; B = 16'h00A8; #100;
A = 16'h00AF; B = 16'h00A9; #100;
A = 16'h00AF; B = 16'h00AA; #100;
A = 16'h00AF; B = 16'h00AB; #100;
A = 16'h00AF; B = 16'h00AC; #100;
A = 16'h00AF; B = 16'h00AD; #100;
A = 16'h00AF; B = 16'h00AE; #100;
A = 16'h00AF; B = 16'h00AF; #100;
A = 16'h00AF; B = 16'h00B0; #100;
A = 16'h00AF; B = 16'h00B1; #100;
A = 16'h00AF; B = 16'h00B2; #100;
A = 16'h00AF; B = 16'h00B3; #100;
A = 16'h00AF; B = 16'h00B4; #100;
A = 16'h00AF; B = 16'h00B5; #100;
A = 16'h00AF; B = 16'h00B6; #100;
A = 16'h00AF; B = 16'h00B7; #100;
A = 16'h00AF; B = 16'h00B8; #100;
A = 16'h00AF; B = 16'h00B9; #100;
A = 16'h00AF; B = 16'h00BA; #100;
A = 16'h00AF; B = 16'h00BB; #100;
A = 16'h00AF; B = 16'h00BC; #100;
A = 16'h00AF; B = 16'h00BD; #100;
A = 16'h00AF; B = 16'h00BE; #100;
A = 16'h00AF; B = 16'h00BF; #100;
A = 16'h00AF; B = 16'h00C0; #100;
A = 16'h00AF; B = 16'h00C1; #100;
A = 16'h00AF; B = 16'h00C2; #100;
A = 16'h00AF; B = 16'h00C3; #100;
A = 16'h00AF; B = 16'h00C4; #100;
A = 16'h00AF; B = 16'h00C5; #100;
A = 16'h00AF; B = 16'h00C6; #100;
A = 16'h00AF; B = 16'h00C7; #100;
A = 16'h00AF; B = 16'h00C8; #100;
A = 16'h00AF; B = 16'h00C9; #100;
A = 16'h00AF; B = 16'h00CA; #100;
A = 16'h00AF; B = 16'h00CB; #100;
A = 16'h00AF; B = 16'h00CC; #100;
A = 16'h00AF; B = 16'h00CD; #100;
A = 16'h00AF; B = 16'h00CE; #100;
A = 16'h00AF; B = 16'h00CF; #100;
A = 16'h00AF; B = 16'h00D0; #100;
A = 16'h00AF; B = 16'h00D1; #100;
A = 16'h00AF; B = 16'h00D2; #100;
A = 16'h00AF; B = 16'h00D3; #100;
A = 16'h00AF; B = 16'h00D4; #100;
A = 16'h00AF; B = 16'h00D5; #100;
A = 16'h00AF; B = 16'h00D6; #100;
A = 16'h00AF; B = 16'h00D7; #100;
A = 16'h00AF; B = 16'h00D8; #100;
A = 16'h00AF; B = 16'h00D9; #100;
A = 16'h00AF; B = 16'h00DA; #100;
A = 16'h00AF; B = 16'h00DB; #100;
A = 16'h00AF; B = 16'h00DC; #100;
A = 16'h00AF; B = 16'h00DD; #100;
A = 16'h00AF; B = 16'h00DE; #100;
A = 16'h00AF; B = 16'h00DF; #100;
A = 16'h00AF; B = 16'h00E0; #100;
A = 16'h00AF; B = 16'h00E1; #100;
A = 16'h00AF; B = 16'h00E2; #100;
A = 16'h00AF; B = 16'h00E3; #100;
A = 16'h00AF; B = 16'h00E4; #100;
A = 16'h00AF; B = 16'h00E5; #100;
A = 16'h00AF; B = 16'h00E6; #100;
A = 16'h00AF; B = 16'h00E7; #100;
A = 16'h00AF; B = 16'h00E8; #100;
A = 16'h00AF; B = 16'h00E9; #100;
A = 16'h00AF; B = 16'h00EA; #100;
A = 16'h00AF; B = 16'h00EB; #100;
A = 16'h00AF; B = 16'h00EC; #100;
A = 16'h00AF; B = 16'h00ED; #100;
A = 16'h00AF; B = 16'h00EE; #100;
A = 16'h00AF; B = 16'h00EF; #100;
A = 16'h00AF; B = 16'h00F0; #100;
A = 16'h00AF; B = 16'h00F1; #100;
A = 16'h00AF; B = 16'h00F2; #100;
A = 16'h00AF; B = 16'h00F3; #100;
A = 16'h00AF; B = 16'h00F4; #100;
A = 16'h00AF; B = 16'h00F5; #100;
A = 16'h00AF; B = 16'h00F6; #100;
A = 16'h00AF; B = 16'h00F7; #100;
A = 16'h00AF; B = 16'h00F8; #100;
A = 16'h00AF; B = 16'h00F9; #100;
A = 16'h00AF; B = 16'h00FA; #100;
A = 16'h00AF; B = 16'h00FB; #100;
A = 16'h00AF; B = 16'h00FC; #100;
A = 16'h00AF; B = 16'h00FD; #100;
A = 16'h00AF; B = 16'h00FE; #100;
A = 16'h00AF; B = 16'h00FF; #100;
A = 16'h00B0; B = 16'h000; #100;
A = 16'h00B0; B = 16'h001; #100;
A = 16'h00B0; B = 16'h002; #100;
A = 16'h00B0; B = 16'h003; #100;
A = 16'h00B0; B = 16'h004; #100;
A = 16'h00B0; B = 16'h005; #100;
A = 16'h00B0; B = 16'h006; #100;
A = 16'h00B0; B = 16'h007; #100;
A = 16'h00B0; B = 16'h008; #100;
A = 16'h00B0; B = 16'h009; #100;
A = 16'h00B0; B = 16'h00A; #100;
A = 16'h00B0; B = 16'h00B; #100;
A = 16'h00B0; B = 16'h00C; #100;
A = 16'h00B0; B = 16'h00D; #100;
A = 16'h00B0; B = 16'h00E; #100;
A = 16'h00B0; B = 16'h00F; #100;
A = 16'h00B0; B = 16'h0010; #100;
A = 16'h00B0; B = 16'h0011; #100;
A = 16'h00B0; B = 16'h0012; #100;
A = 16'h00B0; B = 16'h0013; #100;
A = 16'h00B0; B = 16'h0014; #100;
A = 16'h00B0; B = 16'h0015; #100;
A = 16'h00B0; B = 16'h0016; #100;
A = 16'h00B0; B = 16'h0017; #100;
A = 16'h00B0; B = 16'h0018; #100;
A = 16'h00B0; B = 16'h0019; #100;
A = 16'h00B0; B = 16'h001A; #100;
A = 16'h00B0; B = 16'h001B; #100;
A = 16'h00B0; B = 16'h001C; #100;
A = 16'h00B0; B = 16'h001D; #100;
A = 16'h00B0; B = 16'h001E; #100;
A = 16'h00B0; B = 16'h001F; #100;
A = 16'h00B0; B = 16'h0020; #100;
A = 16'h00B0; B = 16'h0021; #100;
A = 16'h00B0; B = 16'h0022; #100;
A = 16'h00B0; B = 16'h0023; #100;
A = 16'h00B0; B = 16'h0024; #100;
A = 16'h00B0; B = 16'h0025; #100;
A = 16'h00B0; B = 16'h0026; #100;
A = 16'h00B0; B = 16'h0027; #100;
A = 16'h00B0; B = 16'h0028; #100;
A = 16'h00B0; B = 16'h0029; #100;
A = 16'h00B0; B = 16'h002A; #100;
A = 16'h00B0; B = 16'h002B; #100;
A = 16'h00B0; B = 16'h002C; #100;
A = 16'h00B0; B = 16'h002D; #100;
A = 16'h00B0; B = 16'h002E; #100;
A = 16'h00B0; B = 16'h002F; #100;
A = 16'h00B0; B = 16'h0030; #100;
A = 16'h00B0; B = 16'h0031; #100;
A = 16'h00B0; B = 16'h0032; #100;
A = 16'h00B0; B = 16'h0033; #100;
A = 16'h00B0; B = 16'h0034; #100;
A = 16'h00B0; B = 16'h0035; #100;
A = 16'h00B0; B = 16'h0036; #100;
A = 16'h00B0; B = 16'h0037; #100;
A = 16'h00B0; B = 16'h0038; #100;
A = 16'h00B0; B = 16'h0039; #100;
A = 16'h00B0; B = 16'h003A; #100;
A = 16'h00B0; B = 16'h003B; #100;
A = 16'h00B0; B = 16'h003C; #100;
A = 16'h00B0; B = 16'h003D; #100;
A = 16'h00B0; B = 16'h003E; #100;
A = 16'h00B0; B = 16'h003F; #100;
A = 16'h00B0; B = 16'h0040; #100;
A = 16'h00B0; B = 16'h0041; #100;
A = 16'h00B0; B = 16'h0042; #100;
A = 16'h00B0; B = 16'h0043; #100;
A = 16'h00B0; B = 16'h0044; #100;
A = 16'h00B0; B = 16'h0045; #100;
A = 16'h00B0; B = 16'h0046; #100;
A = 16'h00B0; B = 16'h0047; #100;
A = 16'h00B0; B = 16'h0048; #100;
A = 16'h00B0; B = 16'h0049; #100;
A = 16'h00B0; B = 16'h004A; #100;
A = 16'h00B0; B = 16'h004B; #100;
A = 16'h00B0; B = 16'h004C; #100;
A = 16'h00B0; B = 16'h004D; #100;
A = 16'h00B0; B = 16'h004E; #100;
A = 16'h00B0; B = 16'h004F; #100;
A = 16'h00B0; B = 16'h0050; #100;
A = 16'h00B0; B = 16'h0051; #100;
A = 16'h00B0; B = 16'h0052; #100;
A = 16'h00B0; B = 16'h0053; #100;
A = 16'h00B0; B = 16'h0054; #100;
A = 16'h00B0; B = 16'h0055; #100;
A = 16'h00B0; B = 16'h0056; #100;
A = 16'h00B0; B = 16'h0057; #100;
A = 16'h00B0; B = 16'h0058; #100;
A = 16'h00B0; B = 16'h0059; #100;
A = 16'h00B0; B = 16'h005A; #100;
A = 16'h00B0; B = 16'h005B; #100;
A = 16'h00B0; B = 16'h005C; #100;
A = 16'h00B0; B = 16'h005D; #100;
A = 16'h00B0; B = 16'h005E; #100;
A = 16'h00B0; B = 16'h005F; #100;
A = 16'h00B0; B = 16'h0060; #100;
A = 16'h00B0; B = 16'h0061; #100;
A = 16'h00B0; B = 16'h0062; #100;
A = 16'h00B0; B = 16'h0063; #100;
A = 16'h00B0; B = 16'h0064; #100;
A = 16'h00B0; B = 16'h0065; #100;
A = 16'h00B0; B = 16'h0066; #100;
A = 16'h00B0; B = 16'h0067; #100;
A = 16'h00B0; B = 16'h0068; #100;
A = 16'h00B0; B = 16'h0069; #100;
A = 16'h00B0; B = 16'h006A; #100;
A = 16'h00B0; B = 16'h006B; #100;
A = 16'h00B0; B = 16'h006C; #100;
A = 16'h00B0; B = 16'h006D; #100;
A = 16'h00B0; B = 16'h006E; #100;
A = 16'h00B0; B = 16'h006F; #100;
A = 16'h00B0; B = 16'h0070; #100;
A = 16'h00B0; B = 16'h0071; #100;
A = 16'h00B0; B = 16'h0072; #100;
A = 16'h00B0; B = 16'h0073; #100;
A = 16'h00B0; B = 16'h0074; #100;
A = 16'h00B0; B = 16'h0075; #100;
A = 16'h00B0; B = 16'h0076; #100;
A = 16'h00B0; B = 16'h0077; #100;
A = 16'h00B0; B = 16'h0078; #100;
A = 16'h00B0; B = 16'h0079; #100;
A = 16'h00B0; B = 16'h007A; #100;
A = 16'h00B0; B = 16'h007B; #100;
A = 16'h00B0; B = 16'h007C; #100;
A = 16'h00B0; B = 16'h007D; #100;
A = 16'h00B0; B = 16'h007E; #100;
A = 16'h00B0; B = 16'h007F; #100;
A = 16'h00B0; B = 16'h0080; #100;
A = 16'h00B0; B = 16'h0081; #100;
A = 16'h00B0; B = 16'h0082; #100;
A = 16'h00B0; B = 16'h0083; #100;
A = 16'h00B0; B = 16'h0084; #100;
A = 16'h00B0; B = 16'h0085; #100;
A = 16'h00B0; B = 16'h0086; #100;
A = 16'h00B0; B = 16'h0087; #100;
A = 16'h00B0; B = 16'h0088; #100;
A = 16'h00B0; B = 16'h0089; #100;
A = 16'h00B0; B = 16'h008A; #100;
A = 16'h00B0; B = 16'h008B; #100;
A = 16'h00B0; B = 16'h008C; #100;
A = 16'h00B0; B = 16'h008D; #100;
A = 16'h00B0; B = 16'h008E; #100;
A = 16'h00B0; B = 16'h008F; #100;
A = 16'h00B0; B = 16'h0090; #100;
A = 16'h00B0; B = 16'h0091; #100;
A = 16'h00B0; B = 16'h0092; #100;
A = 16'h00B0; B = 16'h0093; #100;
A = 16'h00B0; B = 16'h0094; #100;
A = 16'h00B0; B = 16'h0095; #100;
A = 16'h00B0; B = 16'h0096; #100;
A = 16'h00B0; B = 16'h0097; #100;
A = 16'h00B0; B = 16'h0098; #100;
A = 16'h00B0; B = 16'h0099; #100;
A = 16'h00B0; B = 16'h009A; #100;
A = 16'h00B0; B = 16'h009B; #100;
A = 16'h00B0; B = 16'h009C; #100;
A = 16'h00B0; B = 16'h009D; #100;
A = 16'h00B0; B = 16'h009E; #100;
A = 16'h00B0; B = 16'h009F; #100;
A = 16'h00B0; B = 16'h00A0; #100;
A = 16'h00B0; B = 16'h00A1; #100;
A = 16'h00B0; B = 16'h00A2; #100;
A = 16'h00B0; B = 16'h00A3; #100;
A = 16'h00B0; B = 16'h00A4; #100;
A = 16'h00B0; B = 16'h00A5; #100;
A = 16'h00B0; B = 16'h00A6; #100;
A = 16'h00B0; B = 16'h00A7; #100;
A = 16'h00B0; B = 16'h00A8; #100;
A = 16'h00B0; B = 16'h00A9; #100;
A = 16'h00B0; B = 16'h00AA; #100;
A = 16'h00B0; B = 16'h00AB; #100;
A = 16'h00B0; B = 16'h00AC; #100;
A = 16'h00B0; B = 16'h00AD; #100;
A = 16'h00B0; B = 16'h00AE; #100;
A = 16'h00B0; B = 16'h00AF; #100;
A = 16'h00B0; B = 16'h00B0; #100;
A = 16'h00B0; B = 16'h00B1; #100;
A = 16'h00B0; B = 16'h00B2; #100;
A = 16'h00B0; B = 16'h00B3; #100;
A = 16'h00B0; B = 16'h00B4; #100;
A = 16'h00B0; B = 16'h00B5; #100;
A = 16'h00B0; B = 16'h00B6; #100;
A = 16'h00B0; B = 16'h00B7; #100;
A = 16'h00B0; B = 16'h00B8; #100;
A = 16'h00B0; B = 16'h00B9; #100;
A = 16'h00B0; B = 16'h00BA; #100;
A = 16'h00B0; B = 16'h00BB; #100;
A = 16'h00B0; B = 16'h00BC; #100;
A = 16'h00B0; B = 16'h00BD; #100;
A = 16'h00B0; B = 16'h00BE; #100;
A = 16'h00B0; B = 16'h00BF; #100;
A = 16'h00B0; B = 16'h00C0; #100;
A = 16'h00B0; B = 16'h00C1; #100;
A = 16'h00B0; B = 16'h00C2; #100;
A = 16'h00B0; B = 16'h00C3; #100;
A = 16'h00B0; B = 16'h00C4; #100;
A = 16'h00B0; B = 16'h00C5; #100;
A = 16'h00B0; B = 16'h00C6; #100;
A = 16'h00B0; B = 16'h00C7; #100;
A = 16'h00B0; B = 16'h00C8; #100;
A = 16'h00B0; B = 16'h00C9; #100;
A = 16'h00B0; B = 16'h00CA; #100;
A = 16'h00B0; B = 16'h00CB; #100;
A = 16'h00B0; B = 16'h00CC; #100;
A = 16'h00B0; B = 16'h00CD; #100;
A = 16'h00B0; B = 16'h00CE; #100;
A = 16'h00B0; B = 16'h00CF; #100;
A = 16'h00B0; B = 16'h00D0; #100;
A = 16'h00B0; B = 16'h00D1; #100;
A = 16'h00B0; B = 16'h00D2; #100;
A = 16'h00B0; B = 16'h00D3; #100;
A = 16'h00B0; B = 16'h00D4; #100;
A = 16'h00B0; B = 16'h00D5; #100;
A = 16'h00B0; B = 16'h00D6; #100;
A = 16'h00B0; B = 16'h00D7; #100;
A = 16'h00B0; B = 16'h00D8; #100;
A = 16'h00B0; B = 16'h00D9; #100;
A = 16'h00B0; B = 16'h00DA; #100;
A = 16'h00B0; B = 16'h00DB; #100;
A = 16'h00B0; B = 16'h00DC; #100;
A = 16'h00B0; B = 16'h00DD; #100;
A = 16'h00B0; B = 16'h00DE; #100;
A = 16'h00B0; B = 16'h00DF; #100;
A = 16'h00B0; B = 16'h00E0; #100;
A = 16'h00B0; B = 16'h00E1; #100;
A = 16'h00B0; B = 16'h00E2; #100;
A = 16'h00B0; B = 16'h00E3; #100;
A = 16'h00B0; B = 16'h00E4; #100;
A = 16'h00B0; B = 16'h00E5; #100;
A = 16'h00B0; B = 16'h00E6; #100;
A = 16'h00B0; B = 16'h00E7; #100;
A = 16'h00B0; B = 16'h00E8; #100;
A = 16'h00B0; B = 16'h00E9; #100;
A = 16'h00B0; B = 16'h00EA; #100;
A = 16'h00B0; B = 16'h00EB; #100;
A = 16'h00B0; B = 16'h00EC; #100;
A = 16'h00B0; B = 16'h00ED; #100;
A = 16'h00B0; B = 16'h00EE; #100;
A = 16'h00B0; B = 16'h00EF; #100;
A = 16'h00B0; B = 16'h00F0; #100;
A = 16'h00B0; B = 16'h00F1; #100;
A = 16'h00B0; B = 16'h00F2; #100;
A = 16'h00B0; B = 16'h00F3; #100;
A = 16'h00B0; B = 16'h00F4; #100;
A = 16'h00B0; B = 16'h00F5; #100;
A = 16'h00B0; B = 16'h00F6; #100;
A = 16'h00B0; B = 16'h00F7; #100;
A = 16'h00B0; B = 16'h00F8; #100;
A = 16'h00B0; B = 16'h00F9; #100;
A = 16'h00B0; B = 16'h00FA; #100;
A = 16'h00B0; B = 16'h00FB; #100;
A = 16'h00B0; B = 16'h00FC; #100;
A = 16'h00B0; B = 16'h00FD; #100;
A = 16'h00B0; B = 16'h00FE; #100;
A = 16'h00B0; B = 16'h00FF; #100;
A = 16'h00B1; B = 16'h000; #100;
A = 16'h00B1; B = 16'h001; #100;
A = 16'h00B1; B = 16'h002; #100;
A = 16'h00B1; B = 16'h003; #100;
A = 16'h00B1; B = 16'h004; #100;
A = 16'h00B1; B = 16'h005; #100;
A = 16'h00B1; B = 16'h006; #100;
A = 16'h00B1; B = 16'h007; #100;
A = 16'h00B1; B = 16'h008; #100;
A = 16'h00B1; B = 16'h009; #100;
A = 16'h00B1; B = 16'h00A; #100;
A = 16'h00B1; B = 16'h00B; #100;
A = 16'h00B1; B = 16'h00C; #100;
A = 16'h00B1; B = 16'h00D; #100;
A = 16'h00B1; B = 16'h00E; #100;
A = 16'h00B1; B = 16'h00F; #100;
A = 16'h00B1; B = 16'h0010; #100;
A = 16'h00B1; B = 16'h0011; #100;
A = 16'h00B1; B = 16'h0012; #100;
A = 16'h00B1; B = 16'h0013; #100;
A = 16'h00B1; B = 16'h0014; #100;
A = 16'h00B1; B = 16'h0015; #100;
A = 16'h00B1; B = 16'h0016; #100;
A = 16'h00B1; B = 16'h0017; #100;
A = 16'h00B1; B = 16'h0018; #100;
A = 16'h00B1; B = 16'h0019; #100;
A = 16'h00B1; B = 16'h001A; #100;
A = 16'h00B1; B = 16'h001B; #100;
A = 16'h00B1; B = 16'h001C; #100;
A = 16'h00B1; B = 16'h001D; #100;
A = 16'h00B1; B = 16'h001E; #100;
A = 16'h00B1; B = 16'h001F; #100;
A = 16'h00B1; B = 16'h0020; #100;
A = 16'h00B1; B = 16'h0021; #100;
A = 16'h00B1; B = 16'h0022; #100;
A = 16'h00B1; B = 16'h0023; #100;
A = 16'h00B1; B = 16'h0024; #100;
A = 16'h00B1; B = 16'h0025; #100;
A = 16'h00B1; B = 16'h0026; #100;
A = 16'h00B1; B = 16'h0027; #100;
A = 16'h00B1; B = 16'h0028; #100;
A = 16'h00B1; B = 16'h0029; #100;
A = 16'h00B1; B = 16'h002A; #100;
A = 16'h00B1; B = 16'h002B; #100;
A = 16'h00B1; B = 16'h002C; #100;
A = 16'h00B1; B = 16'h002D; #100;
A = 16'h00B1; B = 16'h002E; #100;
A = 16'h00B1; B = 16'h002F; #100;
A = 16'h00B1; B = 16'h0030; #100;
A = 16'h00B1; B = 16'h0031; #100;
A = 16'h00B1; B = 16'h0032; #100;
A = 16'h00B1; B = 16'h0033; #100;
A = 16'h00B1; B = 16'h0034; #100;
A = 16'h00B1; B = 16'h0035; #100;
A = 16'h00B1; B = 16'h0036; #100;
A = 16'h00B1; B = 16'h0037; #100;
A = 16'h00B1; B = 16'h0038; #100;
A = 16'h00B1; B = 16'h0039; #100;
A = 16'h00B1; B = 16'h003A; #100;
A = 16'h00B1; B = 16'h003B; #100;
A = 16'h00B1; B = 16'h003C; #100;
A = 16'h00B1; B = 16'h003D; #100;
A = 16'h00B1; B = 16'h003E; #100;
A = 16'h00B1; B = 16'h003F; #100;
A = 16'h00B1; B = 16'h0040; #100;
A = 16'h00B1; B = 16'h0041; #100;
A = 16'h00B1; B = 16'h0042; #100;
A = 16'h00B1; B = 16'h0043; #100;
A = 16'h00B1; B = 16'h0044; #100;
A = 16'h00B1; B = 16'h0045; #100;
A = 16'h00B1; B = 16'h0046; #100;
A = 16'h00B1; B = 16'h0047; #100;
A = 16'h00B1; B = 16'h0048; #100;
A = 16'h00B1; B = 16'h0049; #100;
A = 16'h00B1; B = 16'h004A; #100;
A = 16'h00B1; B = 16'h004B; #100;
A = 16'h00B1; B = 16'h004C; #100;
A = 16'h00B1; B = 16'h004D; #100;
A = 16'h00B1; B = 16'h004E; #100;
A = 16'h00B1; B = 16'h004F; #100;
A = 16'h00B1; B = 16'h0050; #100;
A = 16'h00B1; B = 16'h0051; #100;
A = 16'h00B1; B = 16'h0052; #100;
A = 16'h00B1; B = 16'h0053; #100;
A = 16'h00B1; B = 16'h0054; #100;
A = 16'h00B1; B = 16'h0055; #100;
A = 16'h00B1; B = 16'h0056; #100;
A = 16'h00B1; B = 16'h0057; #100;
A = 16'h00B1; B = 16'h0058; #100;
A = 16'h00B1; B = 16'h0059; #100;
A = 16'h00B1; B = 16'h005A; #100;
A = 16'h00B1; B = 16'h005B; #100;
A = 16'h00B1; B = 16'h005C; #100;
A = 16'h00B1; B = 16'h005D; #100;
A = 16'h00B1; B = 16'h005E; #100;
A = 16'h00B1; B = 16'h005F; #100;
A = 16'h00B1; B = 16'h0060; #100;
A = 16'h00B1; B = 16'h0061; #100;
A = 16'h00B1; B = 16'h0062; #100;
A = 16'h00B1; B = 16'h0063; #100;
A = 16'h00B1; B = 16'h0064; #100;
A = 16'h00B1; B = 16'h0065; #100;
A = 16'h00B1; B = 16'h0066; #100;
A = 16'h00B1; B = 16'h0067; #100;
A = 16'h00B1; B = 16'h0068; #100;
A = 16'h00B1; B = 16'h0069; #100;
A = 16'h00B1; B = 16'h006A; #100;
A = 16'h00B1; B = 16'h006B; #100;
A = 16'h00B1; B = 16'h006C; #100;
A = 16'h00B1; B = 16'h006D; #100;
A = 16'h00B1; B = 16'h006E; #100;
A = 16'h00B1; B = 16'h006F; #100;
A = 16'h00B1; B = 16'h0070; #100;
A = 16'h00B1; B = 16'h0071; #100;
A = 16'h00B1; B = 16'h0072; #100;
A = 16'h00B1; B = 16'h0073; #100;
A = 16'h00B1; B = 16'h0074; #100;
A = 16'h00B1; B = 16'h0075; #100;
A = 16'h00B1; B = 16'h0076; #100;
A = 16'h00B1; B = 16'h0077; #100;
A = 16'h00B1; B = 16'h0078; #100;
A = 16'h00B1; B = 16'h0079; #100;
A = 16'h00B1; B = 16'h007A; #100;
A = 16'h00B1; B = 16'h007B; #100;
A = 16'h00B1; B = 16'h007C; #100;
A = 16'h00B1; B = 16'h007D; #100;
A = 16'h00B1; B = 16'h007E; #100;
A = 16'h00B1; B = 16'h007F; #100;
A = 16'h00B1; B = 16'h0080; #100;
A = 16'h00B1; B = 16'h0081; #100;
A = 16'h00B1; B = 16'h0082; #100;
A = 16'h00B1; B = 16'h0083; #100;
A = 16'h00B1; B = 16'h0084; #100;
A = 16'h00B1; B = 16'h0085; #100;
A = 16'h00B1; B = 16'h0086; #100;
A = 16'h00B1; B = 16'h0087; #100;
A = 16'h00B1; B = 16'h0088; #100;
A = 16'h00B1; B = 16'h0089; #100;
A = 16'h00B1; B = 16'h008A; #100;
A = 16'h00B1; B = 16'h008B; #100;
A = 16'h00B1; B = 16'h008C; #100;
A = 16'h00B1; B = 16'h008D; #100;
A = 16'h00B1; B = 16'h008E; #100;
A = 16'h00B1; B = 16'h008F; #100;
A = 16'h00B1; B = 16'h0090; #100;
A = 16'h00B1; B = 16'h0091; #100;
A = 16'h00B1; B = 16'h0092; #100;
A = 16'h00B1; B = 16'h0093; #100;
A = 16'h00B1; B = 16'h0094; #100;
A = 16'h00B1; B = 16'h0095; #100;
A = 16'h00B1; B = 16'h0096; #100;
A = 16'h00B1; B = 16'h0097; #100;
A = 16'h00B1; B = 16'h0098; #100;
A = 16'h00B1; B = 16'h0099; #100;
A = 16'h00B1; B = 16'h009A; #100;
A = 16'h00B1; B = 16'h009B; #100;
A = 16'h00B1; B = 16'h009C; #100;
A = 16'h00B1; B = 16'h009D; #100;
A = 16'h00B1; B = 16'h009E; #100;
A = 16'h00B1; B = 16'h009F; #100;
A = 16'h00B1; B = 16'h00A0; #100;
A = 16'h00B1; B = 16'h00A1; #100;
A = 16'h00B1; B = 16'h00A2; #100;
A = 16'h00B1; B = 16'h00A3; #100;
A = 16'h00B1; B = 16'h00A4; #100;
A = 16'h00B1; B = 16'h00A5; #100;
A = 16'h00B1; B = 16'h00A6; #100;
A = 16'h00B1; B = 16'h00A7; #100;
A = 16'h00B1; B = 16'h00A8; #100;
A = 16'h00B1; B = 16'h00A9; #100;
A = 16'h00B1; B = 16'h00AA; #100;
A = 16'h00B1; B = 16'h00AB; #100;
A = 16'h00B1; B = 16'h00AC; #100;
A = 16'h00B1; B = 16'h00AD; #100;
A = 16'h00B1; B = 16'h00AE; #100;
A = 16'h00B1; B = 16'h00AF; #100;
A = 16'h00B1; B = 16'h00B0; #100;
A = 16'h00B1; B = 16'h00B1; #100;
A = 16'h00B1; B = 16'h00B2; #100;
A = 16'h00B1; B = 16'h00B3; #100;
A = 16'h00B1; B = 16'h00B4; #100;
A = 16'h00B1; B = 16'h00B5; #100;
A = 16'h00B1; B = 16'h00B6; #100;
A = 16'h00B1; B = 16'h00B7; #100;
A = 16'h00B1; B = 16'h00B8; #100;
A = 16'h00B1; B = 16'h00B9; #100;
A = 16'h00B1; B = 16'h00BA; #100;
A = 16'h00B1; B = 16'h00BB; #100;
A = 16'h00B1; B = 16'h00BC; #100;
A = 16'h00B1; B = 16'h00BD; #100;
A = 16'h00B1; B = 16'h00BE; #100;
A = 16'h00B1; B = 16'h00BF; #100;
A = 16'h00B1; B = 16'h00C0; #100;
A = 16'h00B1; B = 16'h00C1; #100;
A = 16'h00B1; B = 16'h00C2; #100;
A = 16'h00B1; B = 16'h00C3; #100;
A = 16'h00B1; B = 16'h00C4; #100;
A = 16'h00B1; B = 16'h00C5; #100;
A = 16'h00B1; B = 16'h00C6; #100;
A = 16'h00B1; B = 16'h00C7; #100;
A = 16'h00B1; B = 16'h00C8; #100;
A = 16'h00B1; B = 16'h00C9; #100;
A = 16'h00B1; B = 16'h00CA; #100;
A = 16'h00B1; B = 16'h00CB; #100;
A = 16'h00B1; B = 16'h00CC; #100;
A = 16'h00B1; B = 16'h00CD; #100;
A = 16'h00B1; B = 16'h00CE; #100;
A = 16'h00B1; B = 16'h00CF; #100;
A = 16'h00B1; B = 16'h00D0; #100;
A = 16'h00B1; B = 16'h00D1; #100;
A = 16'h00B1; B = 16'h00D2; #100;
A = 16'h00B1; B = 16'h00D3; #100;
A = 16'h00B1; B = 16'h00D4; #100;
A = 16'h00B1; B = 16'h00D5; #100;
A = 16'h00B1; B = 16'h00D6; #100;
A = 16'h00B1; B = 16'h00D7; #100;
A = 16'h00B1; B = 16'h00D8; #100;
A = 16'h00B1; B = 16'h00D9; #100;
A = 16'h00B1; B = 16'h00DA; #100;
A = 16'h00B1; B = 16'h00DB; #100;
A = 16'h00B1; B = 16'h00DC; #100;
A = 16'h00B1; B = 16'h00DD; #100;
A = 16'h00B1; B = 16'h00DE; #100;
A = 16'h00B1; B = 16'h00DF; #100;
A = 16'h00B1; B = 16'h00E0; #100;
A = 16'h00B1; B = 16'h00E1; #100;
A = 16'h00B1; B = 16'h00E2; #100;
A = 16'h00B1; B = 16'h00E3; #100;
A = 16'h00B1; B = 16'h00E4; #100;
A = 16'h00B1; B = 16'h00E5; #100;
A = 16'h00B1; B = 16'h00E6; #100;
A = 16'h00B1; B = 16'h00E7; #100;
A = 16'h00B1; B = 16'h00E8; #100;
A = 16'h00B1; B = 16'h00E9; #100;
A = 16'h00B1; B = 16'h00EA; #100;
A = 16'h00B1; B = 16'h00EB; #100;
A = 16'h00B1; B = 16'h00EC; #100;
A = 16'h00B1; B = 16'h00ED; #100;
A = 16'h00B1; B = 16'h00EE; #100;
A = 16'h00B1; B = 16'h00EF; #100;
A = 16'h00B1; B = 16'h00F0; #100;
A = 16'h00B1; B = 16'h00F1; #100;
A = 16'h00B1; B = 16'h00F2; #100;
A = 16'h00B1; B = 16'h00F3; #100;
A = 16'h00B1; B = 16'h00F4; #100;
A = 16'h00B1; B = 16'h00F5; #100;
A = 16'h00B1; B = 16'h00F6; #100;
A = 16'h00B1; B = 16'h00F7; #100;
A = 16'h00B1; B = 16'h00F8; #100;
A = 16'h00B1; B = 16'h00F9; #100;
A = 16'h00B1; B = 16'h00FA; #100;
A = 16'h00B1; B = 16'h00FB; #100;
A = 16'h00B1; B = 16'h00FC; #100;
A = 16'h00B1; B = 16'h00FD; #100;
A = 16'h00B1; B = 16'h00FE; #100;
A = 16'h00B1; B = 16'h00FF; #100;
A = 16'h00B2; B = 16'h000; #100;
A = 16'h00B2; B = 16'h001; #100;
A = 16'h00B2; B = 16'h002; #100;
A = 16'h00B2; B = 16'h003; #100;
A = 16'h00B2; B = 16'h004; #100;
A = 16'h00B2; B = 16'h005; #100;
A = 16'h00B2; B = 16'h006; #100;
A = 16'h00B2; B = 16'h007; #100;
A = 16'h00B2; B = 16'h008; #100;
A = 16'h00B2; B = 16'h009; #100;
A = 16'h00B2; B = 16'h00A; #100;
A = 16'h00B2; B = 16'h00B; #100;
A = 16'h00B2; B = 16'h00C; #100;
A = 16'h00B2; B = 16'h00D; #100;
A = 16'h00B2; B = 16'h00E; #100;
A = 16'h00B2; B = 16'h00F; #100;
A = 16'h00B2; B = 16'h0010; #100;
A = 16'h00B2; B = 16'h0011; #100;
A = 16'h00B2; B = 16'h0012; #100;
A = 16'h00B2; B = 16'h0013; #100;
A = 16'h00B2; B = 16'h0014; #100;
A = 16'h00B2; B = 16'h0015; #100;
A = 16'h00B2; B = 16'h0016; #100;
A = 16'h00B2; B = 16'h0017; #100;
A = 16'h00B2; B = 16'h0018; #100;
A = 16'h00B2; B = 16'h0019; #100;
A = 16'h00B2; B = 16'h001A; #100;
A = 16'h00B2; B = 16'h001B; #100;
A = 16'h00B2; B = 16'h001C; #100;
A = 16'h00B2; B = 16'h001D; #100;
A = 16'h00B2; B = 16'h001E; #100;
A = 16'h00B2; B = 16'h001F; #100;
A = 16'h00B2; B = 16'h0020; #100;
A = 16'h00B2; B = 16'h0021; #100;
A = 16'h00B2; B = 16'h0022; #100;
A = 16'h00B2; B = 16'h0023; #100;
A = 16'h00B2; B = 16'h0024; #100;
A = 16'h00B2; B = 16'h0025; #100;
A = 16'h00B2; B = 16'h0026; #100;
A = 16'h00B2; B = 16'h0027; #100;
A = 16'h00B2; B = 16'h0028; #100;
A = 16'h00B2; B = 16'h0029; #100;
A = 16'h00B2; B = 16'h002A; #100;
A = 16'h00B2; B = 16'h002B; #100;
A = 16'h00B2; B = 16'h002C; #100;
A = 16'h00B2; B = 16'h002D; #100;
A = 16'h00B2; B = 16'h002E; #100;
A = 16'h00B2; B = 16'h002F; #100;
A = 16'h00B2; B = 16'h0030; #100;
A = 16'h00B2; B = 16'h0031; #100;
A = 16'h00B2; B = 16'h0032; #100;
A = 16'h00B2; B = 16'h0033; #100;
A = 16'h00B2; B = 16'h0034; #100;
A = 16'h00B2; B = 16'h0035; #100;
A = 16'h00B2; B = 16'h0036; #100;
A = 16'h00B2; B = 16'h0037; #100;
A = 16'h00B2; B = 16'h0038; #100;
A = 16'h00B2; B = 16'h0039; #100;
A = 16'h00B2; B = 16'h003A; #100;
A = 16'h00B2; B = 16'h003B; #100;
A = 16'h00B2; B = 16'h003C; #100;
A = 16'h00B2; B = 16'h003D; #100;
A = 16'h00B2; B = 16'h003E; #100;
A = 16'h00B2; B = 16'h003F; #100;
A = 16'h00B2; B = 16'h0040; #100;
A = 16'h00B2; B = 16'h0041; #100;
A = 16'h00B2; B = 16'h0042; #100;
A = 16'h00B2; B = 16'h0043; #100;
A = 16'h00B2; B = 16'h0044; #100;
A = 16'h00B2; B = 16'h0045; #100;
A = 16'h00B2; B = 16'h0046; #100;
A = 16'h00B2; B = 16'h0047; #100;
A = 16'h00B2; B = 16'h0048; #100;
A = 16'h00B2; B = 16'h0049; #100;
A = 16'h00B2; B = 16'h004A; #100;
A = 16'h00B2; B = 16'h004B; #100;
A = 16'h00B2; B = 16'h004C; #100;
A = 16'h00B2; B = 16'h004D; #100;
A = 16'h00B2; B = 16'h004E; #100;
A = 16'h00B2; B = 16'h004F; #100;
A = 16'h00B2; B = 16'h0050; #100;
A = 16'h00B2; B = 16'h0051; #100;
A = 16'h00B2; B = 16'h0052; #100;
A = 16'h00B2; B = 16'h0053; #100;
A = 16'h00B2; B = 16'h0054; #100;
A = 16'h00B2; B = 16'h0055; #100;
A = 16'h00B2; B = 16'h0056; #100;
A = 16'h00B2; B = 16'h0057; #100;
A = 16'h00B2; B = 16'h0058; #100;
A = 16'h00B2; B = 16'h0059; #100;
A = 16'h00B2; B = 16'h005A; #100;
A = 16'h00B2; B = 16'h005B; #100;
A = 16'h00B2; B = 16'h005C; #100;
A = 16'h00B2; B = 16'h005D; #100;
A = 16'h00B2; B = 16'h005E; #100;
A = 16'h00B2; B = 16'h005F; #100;
A = 16'h00B2; B = 16'h0060; #100;
A = 16'h00B2; B = 16'h0061; #100;
A = 16'h00B2; B = 16'h0062; #100;
A = 16'h00B2; B = 16'h0063; #100;
A = 16'h00B2; B = 16'h0064; #100;
A = 16'h00B2; B = 16'h0065; #100;
A = 16'h00B2; B = 16'h0066; #100;
A = 16'h00B2; B = 16'h0067; #100;
A = 16'h00B2; B = 16'h0068; #100;
A = 16'h00B2; B = 16'h0069; #100;
A = 16'h00B2; B = 16'h006A; #100;
A = 16'h00B2; B = 16'h006B; #100;
A = 16'h00B2; B = 16'h006C; #100;
A = 16'h00B2; B = 16'h006D; #100;
A = 16'h00B2; B = 16'h006E; #100;
A = 16'h00B2; B = 16'h006F; #100;
A = 16'h00B2; B = 16'h0070; #100;
A = 16'h00B2; B = 16'h0071; #100;
A = 16'h00B2; B = 16'h0072; #100;
A = 16'h00B2; B = 16'h0073; #100;
A = 16'h00B2; B = 16'h0074; #100;
A = 16'h00B2; B = 16'h0075; #100;
A = 16'h00B2; B = 16'h0076; #100;
A = 16'h00B2; B = 16'h0077; #100;
A = 16'h00B2; B = 16'h0078; #100;
A = 16'h00B2; B = 16'h0079; #100;
A = 16'h00B2; B = 16'h007A; #100;
A = 16'h00B2; B = 16'h007B; #100;
A = 16'h00B2; B = 16'h007C; #100;
A = 16'h00B2; B = 16'h007D; #100;
A = 16'h00B2; B = 16'h007E; #100;
A = 16'h00B2; B = 16'h007F; #100;
A = 16'h00B2; B = 16'h0080; #100;
A = 16'h00B2; B = 16'h0081; #100;
A = 16'h00B2; B = 16'h0082; #100;
A = 16'h00B2; B = 16'h0083; #100;
A = 16'h00B2; B = 16'h0084; #100;
A = 16'h00B2; B = 16'h0085; #100;
A = 16'h00B2; B = 16'h0086; #100;
A = 16'h00B2; B = 16'h0087; #100;
A = 16'h00B2; B = 16'h0088; #100;
A = 16'h00B2; B = 16'h0089; #100;
A = 16'h00B2; B = 16'h008A; #100;
A = 16'h00B2; B = 16'h008B; #100;
A = 16'h00B2; B = 16'h008C; #100;
A = 16'h00B2; B = 16'h008D; #100;
A = 16'h00B2; B = 16'h008E; #100;
A = 16'h00B2; B = 16'h008F; #100;
A = 16'h00B2; B = 16'h0090; #100;
A = 16'h00B2; B = 16'h0091; #100;
A = 16'h00B2; B = 16'h0092; #100;
A = 16'h00B2; B = 16'h0093; #100;
A = 16'h00B2; B = 16'h0094; #100;
A = 16'h00B2; B = 16'h0095; #100;
A = 16'h00B2; B = 16'h0096; #100;
A = 16'h00B2; B = 16'h0097; #100;
A = 16'h00B2; B = 16'h0098; #100;
A = 16'h00B2; B = 16'h0099; #100;
A = 16'h00B2; B = 16'h009A; #100;
A = 16'h00B2; B = 16'h009B; #100;
A = 16'h00B2; B = 16'h009C; #100;
A = 16'h00B2; B = 16'h009D; #100;
A = 16'h00B2; B = 16'h009E; #100;
A = 16'h00B2; B = 16'h009F; #100;
A = 16'h00B2; B = 16'h00A0; #100;
A = 16'h00B2; B = 16'h00A1; #100;
A = 16'h00B2; B = 16'h00A2; #100;
A = 16'h00B2; B = 16'h00A3; #100;
A = 16'h00B2; B = 16'h00A4; #100;
A = 16'h00B2; B = 16'h00A5; #100;
A = 16'h00B2; B = 16'h00A6; #100;
A = 16'h00B2; B = 16'h00A7; #100;
A = 16'h00B2; B = 16'h00A8; #100;
A = 16'h00B2; B = 16'h00A9; #100;
A = 16'h00B2; B = 16'h00AA; #100;
A = 16'h00B2; B = 16'h00AB; #100;
A = 16'h00B2; B = 16'h00AC; #100;
A = 16'h00B2; B = 16'h00AD; #100;
A = 16'h00B2; B = 16'h00AE; #100;
A = 16'h00B2; B = 16'h00AF; #100;
A = 16'h00B2; B = 16'h00B0; #100;
A = 16'h00B2; B = 16'h00B1; #100;
A = 16'h00B2; B = 16'h00B2; #100;
A = 16'h00B2; B = 16'h00B3; #100;
A = 16'h00B2; B = 16'h00B4; #100;
A = 16'h00B2; B = 16'h00B5; #100;
A = 16'h00B2; B = 16'h00B6; #100;
A = 16'h00B2; B = 16'h00B7; #100;
A = 16'h00B2; B = 16'h00B8; #100;
A = 16'h00B2; B = 16'h00B9; #100;
A = 16'h00B2; B = 16'h00BA; #100;
A = 16'h00B2; B = 16'h00BB; #100;
A = 16'h00B2; B = 16'h00BC; #100;
A = 16'h00B2; B = 16'h00BD; #100;
A = 16'h00B2; B = 16'h00BE; #100;
A = 16'h00B2; B = 16'h00BF; #100;
A = 16'h00B2; B = 16'h00C0; #100;
A = 16'h00B2; B = 16'h00C1; #100;
A = 16'h00B2; B = 16'h00C2; #100;
A = 16'h00B2; B = 16'h00C3; #100;
A = 16'h00B2; B = 16'h00C4; #100;
A = 16'h00B2; B = 16'h00C5; #100;
A = 16'h00B2; B = 16'h00C6; #100;
A = 16'h00B2; B = 16'h00C7; #100;
A = 16'h00B2; B = 16'h00C8; #100;
A = 16'h00B2; B = 16'h00C9; #100;
A = 16'h00B2; B = 16'h00CA; #100;
A = 16'h00B2; B = 16'h00CB; #100;
A = 16'h00B2; B = 16'h00CC; #100;
A = 16'h00B2; B = 16'h00CD; #100;
A = 16'h00B2; B = 16'h00CE; #100;
A = 16'h00B2; B = 16'h00CF; #100;
A = 16'h00B2; B = 16'h00D0; #100;
A = 16'h00B2; B = 16'h00D1; #100;
A = 16'h00B2; B = 16'h00D2; #100;
A = 16'h00B2; B = 16'h00D3; #100;
A = 16'h00B2; B = 16'h00D4; #100;
A = 16'h00B2; B = 16'h00D5; #100;
A = 16'h00B2; B = 16'h00D6; #100;
A = 16'h00B2; B = 16'h00D7; #100;
A = 16'h00B2; B = 16'h00D8; #100;
A = 16'h00B2; B = 16'h00D9; #100;
A = 16'h00B2; B = 16'h00DA; #100;
A = 16'h00B2; B = 16'h00DB; #100;
A = 16'h00B2; B = 16'h00DC; #100;
A = 16'h00B2; B = 16'h00DD; #100;
A = 16'h00B2; B = 16'h00DE; #100;
A = 16'h00B2; B = 16'h00DF; #100;
A = 16'h00B2; B = 16'h00E0; #100;
A = 16'h00B2; B = 16'h00E1; #100;
A = 16'h00B2; B = 16'h00E2; #100;
A = 16'h00B2; B = 16'h00E3; #100;
A = 16'h00B2; B = 16'h00E4; #100;
A = 16'h00B2; B = 16'h00E5; #100;
A = 16'h00B2; B = 16'h00E6; #100;
A = 16'h00B2; B = 16'h00E7; #100;
A = 16'h00B2; B = 16'h00E8; #100;
A = 16'h00B2; B = 16'h00E9; #100;
A = 16'h00B2; B = 16'h00EA; #100;
A = 16'h00B2; B = 16'h00EB; #100;
A = 16'h00B2; B = 16'h00EC; #100;
A = 16'h00B2; B = 16'h00ED; #100;
A = 16'h00B2; B = 16'h00EE; #100;
A = 16'h00B2; B = 16'h00EF; #100;
A = 16'h00B2; B = 16'h00F0; #100;
A = 16'h00B2; B = 16'h00F1; #100;
A = 16'h00B2; B = 16'h00F2; #100;
A = 16'h00B2; B = 16'h00F3; #100;
A = 16'h00B2; B = 16'h00F4; #100;
A = 16'h00B2; B = 16'h00F5; #100;
A = 16'h00B2; B = 16'h00F6; #100;
A = 16'h00B2; B = 16'h00F7; #100;
A = 16'h00B2; B = 16'h00F8; #100;
A = 16'h00B2; B = 16'h00F9; #100;
A = 16'h00B2; B = 16'h00FA; #100;
A = 16'h00B2; B = 16'h00FB; #100;
A = 16'h00B2; B = 16'h00FC; #100;
A = 16'h00B2; B = 16'h00FD; #100;
A = 16'h00B2; B = 16'h00FE; #100;
A = 16'h00B2; B = 16'h00FF; #100;
A = 16'h00B3; B = 16'h000; #100;
A = 16'h00B3; B = 16'h001; #100;
A = 16'h00B3; B = 16'h002; #100;
A = 16'h00B3; B = 16'h003; #100;
A = 16'h00B3; B = 16'h004; #100;
A = 16'h00B3; B = 16'h005; #100;
A = 16'h00B3; B = 16'h006; #100;
A = 16'h00B3; B = 16'h007; #100;
A = 16'h00B3; B = 16'h008; #100;
A = 16'h00B3; B = 16'h009; #100;
A = 16'h00B3; B = 16'h00A; #100;
A = 16'h00B3; B = 16'h00B; #100;
A = 16'h00B3; B = 16'h00C; #100;
A = 16'h00B3; B = 16'h00D; #100;
A = 16'h00B3; B = 16'h00E; #100;
A = 16'h00B3; B = 16'h00F; #100;
A = 16'h00B3; B = 16'h0010; #100;
A = 16'h00B3; B = 16'h0011; #100;
A = 16'h00B3; B = 16'h0012; #100;
A = 16'h00B3; B = 16'h0013; #100;
A = 16'h00B3; B = 16'h0014; #100;
A = 16'h00B3; B = 16'h0015; #100;
A = 16'h00B3; B = 16'h0016; #100;
A = 16'h00B3; B = 16'h0017; #100;
A = 16'h00B3; B = 16'h0018; #100;
A = 16'h00B3; B = 16'h0019; #100;
A = 16'h00B3; B = 16'h001A; #100;
A = 16'h00B3; B = 16'h001B; #100;
A = 16'h00B3; B = 16'h001C; #100;
A = 16'h00B3; B = 16'h001D; #100;
A = 16'h00B3; B = 16'h001E; #100;
A = 16'h00B3; B = 16'h001F; #100;
A = 16'h00B3; B = 16'h0020; #100;
A = 16'h00B3; B = 16'h0021; #100;
A = 16'h00B3; B = 16'h0022; #100;
A = 16'h00B3; B = 16'h0023; #100;
A = 16'h00B3; B = 16'h0024; #100;
A = 16'h00B3; B = 16'h0025; #100;
A = 16'h00B3; B = 16'h0026; #100;
A = 16'h00B3; B = 16'h0027; #100;
A = 16'h00B3; B = 16'h0028; #100;
A = 16'h00B3; B = 16'h0029; #100;
A = 16'h00B3; B = 16'h002A; #100;
A = 16'h00B3; B = 16'h002B; #100;
A = 16'h00B3; B = 16'h002C; #100;
A = 16'h00B3; B = 16'h002D; #100;
A = 16'h00B3; B = 16'h002E; #100;
A = 16'h00B3; B = 16'h002F; #100;
A = 16'h00B3; B = 16'h0030; #100;
A = 16'h00B3; B = 16'h0031; #100;
A = 16'h00B3; B = 16'h0032; #100;
A = 16'h00B3; B = 16'h0033; #100;
A = 16'h00B3; B = 16'h0034; #100;
A = 16'h00B3; B = 16'h0035; #100;
A = 16'h00B3; B = 16'h0036; #100;
A = 16'h00B3; B = 16'h0037; #100;
A = 16'h00B3; B = 16'h0038; #100;
A = 16'h00B3; B = 16'h0039; #100;
A = 16'h00B3; B = 16'h003A; #100;
A = 16'h00B3; B = 16'h003B; #100;
A = 16'h00B3; B = 16'h003C; #100;
A = 16'h00B3; B = 16'h003D; #100;
A = 16'h00B3; B = 16'h003E; #100;
A = 16'h00B3; B = 16'h003F; #100;
A = 16'h00B3; B = 16'h0040; #100;
A = 16'h00B3; B = 16'h0041; #100;
A = 16'h00B3; B = 16'h0042; #100;
A = 16'h00B3; B = 16'h0043; #100;
A = 16'h00B3; B = 16'h0044; #100;
A = 16'h00B3; B = 16'h0045; #100;
A = 16'h00B3; B = 16'h0046; #100;
A = 16'h00B3; B = 16'h0047; #100;
A = 16'h00B3; B = 16'h0048; #100;
A = 16'h00B3; B = 16'h0049; #100;
A = 16'h00B3; B = 16'h004A; #100;
A = 16'h00B3; B = 16'h004B; #100;
A = 16'h00B3; B = 16'h004C; #100;
A = 16'h00B3; B = 16'h004D; #100;
A = 16'h00B3; B = 16'h004E; #100;
A = 16'h00B3; B = 16'h004F; #100;
A = 16'h00B3; B = 16'h0050; #100;
A = 16'h00B3; B = 16'h0051; #100;
A = 16'h00B3; B = 16'h0052; #100;
A = 16'h00B3; B = 16'h0053; #100;
A = 16'h00B3; B = 16'h0054; #100;
A = 16'h00B3; B = 16'h0055; #100;
A = 16'h00B3; B = 16'h0056; #100;
A = 16'h00B3; B = 16'h0057; #100;
A = 16'h00B3; B = 16'h0058; #100;
A = 16'h00B3; B = 16'h0059; #100;
A = 16'h00B3; B = 16'h005A; #100;
A = 16'h00B3; B = 16'h005B; #100;
A = 16'h00B3; B = 16'h005C; #100;
A = 16'h00B3; B = 16'h005D; #100;
A = 16'h00B3; B = 16'h005E; #100;
A = 16'h00B3; B = 16'h005F; #100;
A = 16'h00B3; B = 16'h0060; #100;
A = 16'h00B3; B = 16'h0061; #100;
A = 16'h00B3; B = 16'h0062; #100;
A = 16'h00B3; B = 16'h0063; #100;
A = 16'h00B3; B = 16'h0064; #100;
A = 16'h00B3; B = 16'h0065; #100;
A = 16'h00B3; B = 16'h0066; #100;
A = 16'h00B3; B = 16'h0067; #100;
A = 16'h00B3; B = 16'h0068; #100;
A = 16'h00B3; B = 16'h0069; #100;
A = 16'h00B3; B = 16'h006A; #100;
A = 16'h00B3; B = 16'h006B; #100;
A = 16'h00B3; B = 16'h006C; #100;
A = 16'h00B3; B = 16'h006D; #100;
A = 16'h00B3; B = 16'h006E; #100;
A = 16'h00B3; B = 16'h006F; #100;
A = 16'h00B3; B = 16'h0070; #100;
A = 16'h00B3; B = 16'h0071; #100;
A = 16'h00B3; B = 16'h0072; #100;
A = 16'h00B3; B = 16'h0073; #100;
A = 16'h00B3; B = 16'h0074; #100;
A = 16'h00B3; B = 16'h0075; #100;
A = 16'h00B3; B = 16'h0076; #100;
A = 16'h00B3; B = 16'h0077; #100;
A = 16'h00B3; B = 16'h0078; #100;
A = 16'h00B3; B = 16'h0079; #100;
A = 16'h00B3; B = 16'h007A; #100;
A = 16'h00B3; B = 16'h007B; #100;
A = 16'h00B3; B = 16'h007C; #100;
A = 16'h00B3; B = 16'h007D; #100;
A = 16'h00B3; B = 16'h007E; #100;
A = 16'h00B3; B = 16'h007F; #100;
A = 16'h00B3; B = 16'h0080; #100;
A = 16'h00B3; B = 16'h0081; #100;
A = 16'h00B3; B = 16'h0082; #100;
A = 16'h00B3; B = 16'h0083; #100;
A = 16'h00B3; B = 16'h0084; #100;
A = 16'h00B3; B = 16'h0085; #100;
A = 16'h00B3; B = 16'h0086; #100;
A = 16'h00B3; B = 16'h0087; #100;
A = 16'h00B3; B = 16'h0088; #100;
A = 16'h00B3; B = 16'h0089; #100;
A = 16'h00B3; B = 16'h008A; #100;
A = 16'h00B3; B = 16'h008B; #100;
A = 16'h00B3; B = 16'h008C; #100;
A = 16'h00B3; B = 16'h008D; #100;
A = 16'h00B3; B = 16'h008E; #100;
A = 16'h00B3; B = 16'h008F; #100;
A = 16'h00B3; B = 16'h0090; #100;
A = 16'h00B3; B = 16'h0091; #100;
A = 16'h00B3; B = 16'h0092; #100;
A = 16'h00B3; B = 16'h0093; #100;
A = 16'h00B3; B = 16'h0094; #100;
A = 16'h00B3; B = 16'h0095; #100;
A = 16'h00B3; B = 16'h0096; #100;
A = 16'h00B3; B = 16'h0097; #100;
A = 16'h00B3; B = 16'h0098; #100;
A = 16'h00B3; B = 16'h0099; #100;
A = 16'h00B3; B = 16'h009A; #100;
A = 16'h00B3; B = 16'h009B; #100;
A = 16'h00B3; B = 16'h009C; #100;
A = 16'h00B3; B = 16'h009D; #100;
A = 16'h00B3; B = 16'h009E; #100;
A = 16'h00B3; B = 16'h009F; #100;
A = 16'h00B3; B = 16'h00A0; #100;
A = 16'h00B3; B = 16'h00A1; #100;
A = 16'h00B3; B = 16'h00A2; #100;
A = 16'h00B3; B = 16'h00A3; #100;
A = 16'h00B3; B = 16'h00A4; #100;
A = 16'h00B3; B = 16'h00A5; #100;
A = 16'h00B3; B = 16'h00A6; #100;
A = 16'h00B3; B = 16'h00A7; #100;
A = 16'h00B3; B = 16'h00A8; #100;
A = 16'h00B3; B = 16'h00A9; #100;
A = 16'h00B3; B = 16'h00AA; #100;
A = 16'h00B3; B = 16'h00AB; #100;
A = 16'h00B3; B = 16'h00AC; #100;
A = 16'h00B3; B = 16'h00AD; #100;
A = 16'h00B3; B = 16'h00AE; #100;
A = 16'h00B3; B = 16'h00AF; #100;
A = 16'h00B3; B = 16'h00B0; #100;
A = 16'h00B3; B = 16'h00B1; #100;
A = 16'h00B3; B = 16'h00B2; #100;
A = 16'h00B3; B = 16'h00B3; #100;
A = 16'h00B3; B = 16'h00B4; #100;
A = 16'h00B3; B = 16'h00B5; #100;
A = 16'h00B3; B = 16'h00B6; #100;
A = 16'h00B3; B = 16'h00B7; #100;
A = 16'h00B3; B = 16'h00B8; #100;
A = 16'h00B3; B = 16'h00B9; #100;
A = 16'h00B3; B = 16'h00BA; #100;
A = 16'h00B3; B = 16'h00BB; #100;
A = 16'h00B3; B = 16'h00BC; #100;
A = 16'h00B3; B = 16'h00BD; #100;
A = 16'h00B3; B = 16'h00BE; #100;
A = 16'h00B3; B = 16'h00BF; #100;
A = 16'h00B3; B = 16'h00C0; #100;
A = 16'h00B3; B = 16'h00C1; #100;
A = 16'h00B3; B = 16'h00C2; #100;
A = 16'h00B3; B = 16'h00C3; #100;
A = 16'h00B3; B = 16'h00C4; #100;
A = 16'h00B3; B = 16'h00C5; #100;
A = 16'h00B3; B = 16'h00C6; #100;
A = 16'h00B3; B = 16'h00C7; #100;
A = 16'h00B3; B = 16'h00C8; #100;
A = 16'h00B3; B = 16'h00C9; #100;
A = 16'h00B3; B = 16'h00CA; #100;
A = 16'h00B3; B = 16'h00CB; #100;
A = 16'h00B3; B = 16'h00CC; #100;
A = 16'h00B3; B = 16'h00CD; #100;
A = 16'h00B3; B = 16'h00CE; #100;
A = 16'h00B3; B = 16'h00CF; #100;
A = 16'h00B3; B = 16'h00D0; #100;
A = 16'h00B3; B = 16'h00D1; #100;
A = 16'h00B3; B = 16'h00D2; #100;
A = 16'h00B3; B = 16'h00D3; #100;
A = 16'h00B3; B = 16'h00D4; #100;
A = 16'h00B3; B = 16'h00D5; #100;
A = 16'h00B3; B = 16'h00D6; #100;
A = 16'h00B3; B = 16'h00D7; #100;
A = 16'h00B3; B = 16'h00D8; #100;
A = 16'h00B3; B = 16'h00D9; #100;
A = 16'h00B3; B = 16'h00DA; #100;
A = 16'h00B3; B = 16'h00DB; #100;
A = 16'h00B3; B = 16'h00DC; #100;
A = 16'h00B3; B = 16'h00DD; #100;
A = 16'h00B3; B = 16'h00DE; #100;
A = 16'h00B3; B = 16'h00DF; #100;
A = 16'h00B3; B = 16'h00E0; #100;
A = 16'h00B3; B = 16'h00E1; #100;
A = 16'h00B3; B = 16'h00E2; #100;
A = 16'h00B3; B = 16'h00E3; #100;
A = 16'h00B3; B = 16'h00E4; #100;
A = 16'h00B3; B = 16'h00E5; #100;
A = 16'h00B3; B = 16'h00E6; #100;
A = 16'h00B3; B = 16'h00E7; #100;
A = 16'h00B3; B = 16'h00E8; #100;
A = 16'h00B3; B = 16'h00E9; #100;
A = 16'h00B3; B = 16'h00EA; #100;
A = 16'h00B3; B = 16'h00EB; #100;
A = 16'h00B3; B = 16'h00EC; #100;
A = 16'h00B3; B = 16'h00ED; #100;
A = 16'h00B3; B = 16'h00EE; #100;
A = 16'h00B3; B = 16'h00EF; #100;
A = 16'h00B3; B = 16'h00F0; #100;
A = 16'h00B3; B = 16'h00F1; #100;
A = 16'h00B3; B = 16'h00F2; #100;
A = 16'h00B3; B = 16'h00F3; #100;
A = 16'h00B3; B = 16'h00F4; #100;
A = 16'h00B3; B = 16'h00F5; #100;
A = 16'h00B3; B = 16'h00F6; #100;
A = 16'h00B3; B = 16'h00F7; #100;
A = 16'h00B3; B = 16'h00F8; #100;
A = 16'h00B3; B = 16'h00F9; #100;
A = 16'h00B3; B = 16'h00FA; #100;
A = 16'h00B3; B = 16'h00FB; #100;
A = 16'h00B3; B = 16'h00FC; #100;
A = 16'h00B3; B = 16'h00FD; #100;
A = 16'h00B3; B = 16'h00FE; #100;
A = 16'h00B3; B = 16'h00FF; #100;
A = 16'h00B4; B = 16'h000; #100;
A = 16'h00B4; B = 16'h001; #100;
A = 16'h00B4; B = 16'h002; #100;
A = 16'h00B4; B = 16'h003; #100;
A = 16'h00B4; B = 16'h004; #100;
A = 16'h00B4; B = 16'h005; #100;
A = 16'h00B4; B = 16'h006; #100;
A = 16'h00B4; B = 16'h007; #100;
A = 16'h00B4; B = 16'h008; #100;
A = 16'h00B4; B = 16'h009; #100;
A = 16'h00B4; B = 16'h00A; #100;
A = 16'h00B4; B = 16'h00B; #100;
A = 16'h00B4; B = 16'h00C; #100;
A = 16'h00B4; B = 16'h00D; #100;
A = 16'h00B4; B = 16'h00E; #100;
A = 16'h00B4; B = 16'h00F; #100;
A = 16'h00B4; B = 16'h0010; #100;
A = 16'h00B4; B = 16'h0011; #100;
A = 16'h00B4; B = 16'h0012; #100;
A = 16'h00B4; B = 16'h0013; #100;
A = 16'h00B4; B = 16'h0014; #100;
A = 16'h00B4; B = 16'h0015; #100;
A = 16'h00B4; B = 16'h0016; #100;
A = 16'h00B4; B = 16'h0017; #100;
A = 16'h00B4; B = 16'h0018; #100;
A = 16'h00B4; B = 16'h0019; #100;
A = 16'h00B4; B = 16'h001A; #100;
A = 16'h00B4; B = 16'h001B; #100;
A = 16'h00B4; B = 16'h001C; #100;
A = 16'h00B4; B = 16'h001D; #100;
A = 16'h00B4; B = 16'h001E; #100;
A = 16'h00B4; B = 16'h001F; #100;
A = 16'h00B4; B = 16'h0020; #100;
A = 16'h00B4; B = 16'h0021; #100;
A = 16'h00B4; B = 16'h0022; #100;
A = 16'h00B4; B = 16'h0023; #100;
A = 16'h00B4; B = 16'h0024; #100;
A = 16'h00B4; B = 16'h0025; #100;
A = 16'h00B4; B = 16'h0026; #100;
A = 16'h00B4; B = 16'h0027; #100;
A = 16'h00B4; B = 16'h0028; #100;
A = 16'h00B4; B = 16'h0029; #100;
A = 16'h00B4; B = 16'h002A; #100;
A = 16'h00B4; B = 16'h002B; #100;
A = 16'h00B4; B = 16'h002C; #100;
A = 16'h00B4; B = 16'h002D; #100;
A = 16'h00B4; B = 16'h002E; #100;
A = 16'h00B4; B = 16'h002F; #100;
A = 16'h00B4; B = 16'h0030; #100;
A = 16'h00B4; B = 16'h0031; #100;
A = 16'h00B4; B = 16'h0032; #100;
A = 16'h00B4; B = 16'h0033; #100;
A = 16'h00B4; B = 16'h0034; #100;
A = 16'h00B4; B = 16'h0035; #100;
A = 16'h00B4; B = 16'h0036; #100;
A = 16'h00B4; B = 16'h0037; #100;
A = 16'h00B4; B = 16'h0038; #100;
A = 16'h00B4; B = 16'h0039; #100;
A = 16'h00B4; B = 16'h003A; #100;
A = 16'h00B4; B = 16'h003B; #100;
A = 16'h00B4; B = 16'h003C; #100;
A = 16'h00B4; B = 16'h003D; #100;
A = 16'h00B4; B = 16'h003E; #100;
A = 16'h00B4; B = 16'h003F; #100;
A = 16'h00B4; B = 16'h0040; #100;
A = 16'h00B4; B = 16'h0041; #100;
A = 16'h00B4; B = 16'h0042; #100;
A = 16'h00B4; B = 16'h0043; #100;
A = 16'h00B4; B = 16'h0044; #100;
A = 16'h00B4; B = 16'h0045; #100;
A = 16'h00B4; B = 16'h0046; #100;
A = 16'h00B4; B = 16'h0047; #100;
A = 16'h00B4; B = 16'h0048; #100;
A = 16'h00B4; B = 16'h0049; #100;
A = 16'h00B4; B = 16'h004A; #100;
A = 16'h00B4; B = 16'h004B; #100;
A = 16'h00B4; B = 16'h004C; #100;
A = 16'h00B4; B = 16'h004D; #100;
A = 16'h00B4; B = 16'h004E; #100;
A = 16'h00B4; B = 16'h004F; #100;
A = 16'h00B4; B = 16'h0050; #100;
A = 16'h00B4; B = 16'h0051; #100;
A = 16'h00B4; B = 16'h0052; #100;
A = 16'h00B4; B = 16'h0053; #100;
A = 16'h00B4; B = 16'h0054; #100;
A = 16'h00B4; B = 16'h0055; #100;
A = 16'h00B4; B = 16'h0056; #100;
A = 16'h00B4; B = 16'h0057; #100;
A = 16'h00B4; B = 16'h0058; #100;
A = 16'h00B4; B = 16'h0059; #100;
A = 16'h00B4; B = 16'h005A; #100;
A = 16'h00B4; B = 16'h005B; #100;
A = 16'h00B4; B = 16'h005C; #100;
A = 16'h00B4; B = 16'h005D; #100;
A = 16'h00B4; B = 16'h005E; #100;
A = 16'h00B4; B = 16'h005F; #100;
A = 16'h00B4; B = 16'h0060; #100;
A = 16'h00B4; B = 16'h0061; #100;
A = 16'h00B4; B = 16'h0062; #100;
A = 16'h00B4; B = 16'h0063; #100;
A = 16'h00B4; B = 16'h0064; #100;
A = 16'h00B4; B = 16'h0065; #100;
A = 16'h00B4; B = 16'h0066; #100;
A = 16'h00B4; B = 16'h0067; #100;
A = 16'h00B4; B = 16'h0068; #100;
A = 16'h00B4; B = 16'h0069; #100;
A = 16'h00B4; B = 16'h006A; #100;
A = 16'h00B4; B = 16'h006B; #100;
A = 16'h00B4; B = 16'h006C; #100;
A = 16'h00B4; B = 16'h006D; #100;
A = 16'h00B4; B = 16'h006E; #100;
A = 16'h00B4; B = 16'h006F; #100;
A = 16'h00B4; B = 16'h0070; #100;
A = 16'h00B4; B = 16'h0071; #100;
A = 16'h00B4; B = 16'h0072; #100;
A = 16'h00B4; B = 16'h0073; #100;
A = 16'h00B4; B = 16'h0074; #100;
A = 16'h00B4; B = 16'h0075; #100;
A = 16'h00B4; B = 16'h0076; #100;
A = 16'h00B4; B = 16'h0077; #100;
A = 16'h00B4; B = 16'h0078; #100;
A = 16'h00B4; B = 16'h0079; #100;
A = 16'h00B4; B = 16'h007A; #100;
A = 16'h00B4; B = 16'h007B; #100;
A = 16'h00B4; B = 16'h007C; #100;
A = 16'h00B4; B = 16'h007D; #100;
A = 16'h00B4; B = 16'h007E; #100;
A = 16'h00B4; B = 16'h007F; #100;
A = 16'h00B4; B = 16'h0080; #100;
A = 16'h00B4; B = 16'h0081; #100;
A = 16'h00B4; B = 16'h0082; #100;
A = 16'h00B4; B = 16'h0083; #100;
A = 16'h00B4; B = 16'h0084; #100;
A = 16'h00B4; B = 16'h0085; #100;
A = 16'h00B4; B = 16'h0086; #100;
A = 16'h00B4; B = 16'h0087; #100;
A = 16'h00B4; B = 16'h0088; #100;
A = 16'h00B4; B = 16'h0089; #100;
A = 16'h00B4; B = 16'h008A; #100;
A = 16'h00B4; B = 16'h008B; #100;
A = 16'h00B4; B = 16'h008C; #100;
A = 16'h00B4; B = 16'h008D; #100;
A = 16'h00B4; B = 16'h008E; #100;
A = 16'h00B4; B = 16'h008F; #100;
A = 16'h00B4; B = 16'h0090; #100;
A = 16'h00B4; B = 16'h0091; #100;
A = 16'h00B4; B = 16'h0092; #100;
A = 16'h00B4; B = 16'h0093; #100;
A = 16'h00B4; B = 16'h0094; #100;
A = 16'h00B4; B = 16'h0095; #100;
A = 16'h00B4; B = 16'h0096; #100;
A = 16'h00B4; B = 16'h0097; #100;
A = 16'h00B4; B = 16'h0098; #100;
A = 16'h00B4; B = 16'h0099; #100;
A = 16'h00B4; B = 16'h009A; #100;
A = 16'h00B4; B = 16'h009B; #100;
A = 16'h00B4; B = 16'h009C; #100;
A = 16'h00B4; B = 16'h009D; #100;
A = 16'h00B4; B = 16'h009E; #100;
A = 16'h00B4; B = 16'h009F; #100;
A = 16'h00B4; B = 16'h00A0; #100;
A = 16'h00B4; B = 16'h00A1; #100;
A = 16'h00B4; B = 16'h00A2; #100;
A = 16'h00B4; B = 16'h00A3; #100;
A = 16'h00B4; B = 16'h00A4; #100;
A = 16'h00B4; B = 16'h00A5; #100;
A = 16'h00B4; B = 16'h00A6; #100;
A = 16'h00B4; B = 16'h00A7; #100;
A = 16'h00B4; B = 16'h00A8; #100;
A = 16'h00B4; B = 16'h00A9; #100;
A = 16'h00B4; B = 16'h00AA; #100;
A = 16'h00B4; B = 16'h00AB; #100;
A = 16'h00B4; B = 16'h00AC; #100;
A = 16'h00B4; B = 16'h00AD; #100;
A = 16'h00B4; B = 16'h00AE; #100;
A = 16'h00B4; B = 16'h00AF; #100;
A = 16'h00B4; B = 16'h00B0; #100;
A = 16'h00B4; B = 16'h00B1; #100;
A = 16'h00B4; B = 16'h00B2; #100;
A = 16'h00B4; B = 16'h00B3; #100;
A = 16'h00B4; B = 16'h00B4; #100;
A = 16'h00B4; B = 16'h00B5; #100;
A = 16'h00B4; B = 16'h00B6; #100;
A = 16'h00B4; B = 16'h00B7; #100;
A = 16'h00B4; B = 16'h00B8; #100;
A = 16'h00B4; B = 16'h00B9; #100;
A = 16'h00B4; B = 16'h00BA; #100;
A = 16'h00B4; B = 16'h00BB; #100;
A = 16'h00B4; B = 16'h00BC; #100;
A = 16'h00B4; B = 16'h00BD; #100;
A = 16'h00B4; B = 16'h00BE; #100;
A = 16'h00B4; B = 16'h00BF; #100;
A = 16'h00B4; B = 16'h00C0; #100;
A = 16'h00B4; B = 16'h00C1; #100;
A = 16'h00B4; B = 16'h00C2; #100;
A = 16'h00B4; B = 16'h00C3; #100;
A = 16'h00B4; B = 16'h00C4; #100;
A = 16'h00B4; B = 16'h00C5; #100;
A = 16'h00B4; B = 16'h00C6; #100;
A = 16'h00B4; B = 16'h00C7; #100;
A = 16'h00B4; B = 16'h00C8; #100;
A = 16'h00B4; B = 16'h00C9; #100;
A = 16'h00B4; B = 16'h00CA; #100;
A = 16'h00B4; B = 16'h00CB; #100;
A = 16'h00B4; B = 16'h00CC; #100;
A = 16'h00B4; B = 16'h00CD; #100;
A = 16'h00B4; B = 16'h00CE; #100;
A = 16'h00B4; B = 16'h00CF; #100;
A = 16'h00B4; B = 16'h00D0; #100;
A = 16'h00B4; B = 16'h00D1; #100;
A = 16'h00B4; B = 16'h00D2; #100;
A = 16'h00B4; B = 16'h00D3; #100;
A = 16'h00B4; B = 16'h00D4; #100;
A = 16'h00B4; B = 16'h00D5; #100;
A = 16'h00B4; B = 16'h00D6; #100;
A = 16'h00B4; B = 16'h00D7; #100;
A = 16'h00B4; B = 16'h00D8; #100;
A = 16'h00B4; B = 16'h00D9; #100;
A = 16'h00B4; B = 16'h00DA; #100;
A = 16'h00B4; B = 16'h00DB; #100;
A = 16'h00B4; B = 16'h00DC; #100;
A = 16'h00B4; B = 16'h00DD; #100;
A = 16'h00B4; B = 16'h00DE; #100;
A = 16'h00B4; B = 16'h00DF; #100;
A = 16'h00B4; B = 16'h00E0; #100;
A = 16'h00B4; B = 16'h00E1; #100;
A = 16'h00B4; B = 16'h00E2; #100;
A = 16'h00B4; B = 16'h00E3; #100;
A = 16'h00B4; B = 16'h00E4; #100;
A = 16'h00B4; B = 16'h00E5; #100;
A = 16'h00B4; B = 16'h00E6; #100;
A = 16'h00B4; B = 16'h00E7; #100;
A = 16'h00B4; B = 16'h00E8; #100;
A = 16'h00B4; B = 16'h00E9; #100;
A = 16'h00B4; B = 16'h00EA; #100;
A = 16'h00B4; B = 16'h00EB; #100;
A = 16'h00B4; B = 16'h00EC; #100;
A = 16'h00B4; B = 16'h00ED; #100;
A = 16'h00B4; B = 16'h00EE; #100;
A = 16'h00B4; B = 16'h00EF; #100;
A = 16'h00B4; B = 16'h00F0; #100;
A = 16'h00B4; B = 16'h00F1; #100;
A = 16'h00B4; B = 16'h00F2; #100;
A = 16'h00B4; B = 16'h00F3; #100;
A = 16'h00B4; B = 16'h00F4; #100;
A = 16'h00B4; B = 16'h00F5; #100;
A = 16'h00B4; B = 16'h00F6; #100;
A = 16'h00B4; B = 16'h00F7; #100;
A = 16'h00B4; B = 16'h00F8; #100;
A = 16'h00B4; B = 16'h00F9; #100;
A = 16'h00B4; B = 16'h00FA; #100;
A = 16'h00B4; B = 16'h00FB; #100;
A = 16'h00B4; B = 16'h00FC; #100;
A = 16'h00B4; B = 16'h00FD; #100;
A = 16'h00B4; B = 16'h00FE; #100;
A = 16'h00B4; B = 16'h00FF; #100;
A = 16'h00B5; B = 16'h000; #100;
A = 16'h00B5; B = 16'h001; #100;
A = 16'h00B5; B = 16'h002; #100;
A = 16'h00B5; B = 16'h003; #100;
A = 16'h00B5; B = 16'h004; #100;
A = 16'h00B5; B = 16'h005; #100;
A = 16'h00B5; B = 16'h006; #100;
A = 16'h00B5; B = 16'h007; #100;
A = 16'h00B5; B = 16'h008; #100;
A = 16'h00B5; B = 16'h009; #100;
A = 16'h00B5; B = 16'h00A; #100;
A = 16'h00B5; B = 16'h00B; #100;
A = 16'h00B5; B = 16'h00C; #100;
A = 16'h00B5; B = 16'h00D; #100;
A = 16'h00B5; B = 16'h00E; #100;
A = 16'h00B5; B = 16'h00F; #100;
A = 16'h00B5; B = 16'h0010; #100;
A = 16'h00B5; B = 16'h0011; #100;
A = 16'h00B5; B = 16'h0012; #100;
A = 16'h00B5; B = 16'h0013; #100;
A = 16'h00B5; B = 16'h0014; #100;
A = 16'h00B5; B = 16'h0015; #100;
A = 16'h00B5; B = 16'h0016; #100;
A = 16'h00B5; B = 16'h0017; #100;
A = 16'h00B5; B = 16'h0018; #100;
A = 16'h00B5; B = 16'h0019; #100;
A = 16'h00B5; B = 16'h001A; #100;
A = 16'h00B5; B = 16'h001B; #100;
A = 16'h00B5; B = 16'h001C; #100;
A = 16'h00B5; B = 16'h001D; #100;
A = 16'h00B5; B = 16'h001E; #100;
A = 16'h00B5; B = 16'h001F; #100;
A = 16'h00B5; B = 16'h0020; #100;
A = 16'h00B5; B = 16'h0021; #100;
A = 16'h00B5; B = 16'h0022; #100;
A = 16'h00B5; B = 16'h0023; #100;
A = 16'h00B5; B = 16'h0024; #100;
A = 16'h00B5; B = 16'h0025; #100;
A = 16'h00B5; B = 16'h0026; #100;
A = 16'h00B5; B = 16'h0027; #100;
A = 16'h00B5; B = 16'h0028; #100;
A = 16'h00B5; B = 16'h0029; #100;
A = 16'h00B5; B = 16'h002A; #100;
A = 16'h00B5; B = 16'h002B; #100;
A = 16'h00B5; B = 16'h002C; #100;
A = 16'h00B5; B = 16'h002D; #100;
A = 16'h00B5; B = 16'h002E; #100;
A = 16'h00B5; B = 16'h002F; #100;
A = 16'h00B5; B = 16'h0030; #100;
A = 16'h00B5; B = 16'h0031; #100;
A = 16'h00B5; B = 16'h0032; #100;
A = 16'h00B5; B = 16'h0033; #100;
A = 16'h00B5; B = 16'h0034; #100;
A = 16'h00B5; B = 16'h0035; #100;
A = 16'h00B5; B = 16'h0036; #100;
A = 16'h00B5; B = 16'h0037; #100;
A = 16'h00B5; B = 16'h0038; #100;
A = 16'h00B5; B = 16'h0039; #100;
A = 16'h00B5; B = 16'h003A; #100;
A = 16'h00B5; B = 16'h003B; #100;
A = 16'h00B5; B = 16'h003C; #100;
A = 16'h00B5; B = 16'h003D; #100;
A = 16'h00B5; B = 16'h003E; #100;
A = 16'h00B5; B = 16'h003F; #100;
A = 16'h00B5; B = 16'h0040; #100;
A = 16'h00B5; B = 16'h0041; #100;
A = 16'h00B5; B = 16'h0042; #100;
A = 16'h00B5; B = 16'h0043; #100;
A = 16'h00B5; B = 16'h0044; #100;
A = 16'h00B5; B = 16'h0045; #100;
A = 16'h00B5; B = 16'h0046; #100;
A = 16'h00B5; B = 16'h0047; #100;
A = 16'h00B5; B = 16'h0048; #100;
A = 16'h00B5; B = 16'h0049; #100;
A = 16'h00B5; B = 16'h004A; #100;
A = 16'h00B5; B = 16'h004B; #100;
A = 16'h00B5; B = 16'h004C; #100;
A = 16'h00B5; B = 16'h004D; #100;
A = 16'h00B5; B = 16'h004E; #100;
A = 16'h00B5; B = 16'h004F; #100;
A = 16'h00B5; B = 16'h0050; #100;
A = 16'h00B5; B = 16'h0051; #100;
A = 16'h00B5; B = 16'h0052; #100;
A = 16'h00B5; B = 16'h0053; #100;
A = 16'h00B5; B = 16'h0054; #100;
A = 16'h00B5; B = 16'h0055; #100;
A = 16'h00B5; B = 16'h0056; #100;
A = 16'h00B5; B = 16'h0057; #100;
A = 16'h00B5; B = 16'h0058; #100;
A = 16'h00B5; B = 16'h0059; #100;
A = 16'h00B5; B = 16'h005A; #100;
A = 16'h00B5; B = 16'h005B; #100;
A = 16'h00B5; B = 16'h005C; #100;
A = 16'h00B5; B = 16'h005D; #100;
A = 16'h00B5; B = 16'h005E; #100;
A = 16'h00B5; B = 16'h005F; #100;
A = 16'h00B5; B = 16'h0060; #100;
A = 16'h00B5; B = 16'h0061; #100;
A = 16'h00B5; B = 16'h0062; #100;
A = 16'h00B5; B = 16'h0063; #100;
A = 16'h00B5; B = 16'h0064; #100;
A = 16'h00B5; B = 16'h0065; #100;
A = 16'h00B5; B = 16'h0066; #100;
A = 16'h00B5; B = 16'h0067; #100;
A = 16'h00B5; B = 16'h0068; #100;
A = 16'h00B5; B = 16'h0069; #100;
A = 16'h00B5; B = 16'h006A; #100;
A = 16'h00B5; B = 16'h006B; #100;
A = 16'h00B5; B = 16'h006C; #100;
A = 16'h00B5; B = 16'h006D; #100;
A = 16'h00B5; B = 16'h006E; #100;
A = 16'h00B5; B = 16'h006F; #100;
A = 16'h00B5; B = 16'h0070; #100;
A = 16'h00B5; B = 16'h0071; #100;
A = 16'h00B5; B = 16'h0072; #100;
A = 16'h00B5; B = 16'h0073; #100;
A = 16'h00B5; B = 16'h0074; #100;
A = 16'h00B5; B = 16'h0075; #100;
A = 16'h00B5; B = 16'h0076; #100;
A = 16'h00B5; B = 16'h0077; #100;
A = 16'h00B5; B = 16'h0078; #100;
A = 16'h00B5; B = 16'h0079; #100;
A = 16'h00B5; B = 16'h007A; #100;
A = 16'h00B5; B = 16'h007B; #100;
A = 16'h00B5; B = 16'h007C; #100;
A = 16'h00B5; B = 16'h007D; #100;
A = 16'h00B5; B = 16'h007E; #100;
A = 16'h00B5; B = 16'h007F; #100;
A = 16'h00B5; B = 16'h0080; #100;
A = 16'h00B5; B = 16'h0081; #100;
A = 16'h00B5; B = 16'h0082; #100;
A = 16'h00B5; B = 16'h0083; #100;
A = 16'h00B5; B = 16'h0084; #100;
A = 16'h00B5; B = 16'h0085; #100;
A = 16'h00B5; B = 16'h0086; #100;
A = 16'h00B5; B = 16'h0087; #100;
A = 16'h00B5; B = 16'h0088; #100;
A = 16'h00B5; B = 16'h0089; #100;
A = 16'h00B5; B = 16'h008A; #100;
A = 16'h00B5; B = 16'h008B; #100;
A = 16'h00B5; B = 16'h008C; #100;
A = 16'h00B5; B = 16'h008D; #100;
A = 16'h00B5; B = 16'h008E; #100;
A = 16'h00B5; B = 16'h008F; #100;
A = 16'h00B5; B = 16'h0090; #100;
A = 16'h00B5; B = 16'h0091; #100;
A = 16'h00B5; B = 16'h0092; #100;
A = 16'h00B5; B = 16'h0093; #100;
A = 16'h00B5; B = 16'h0094; #100;
A = 16'h00B5; B = 16'h0095; #100;
A = 16'h00B5; B = 16'h0096; #100;
A = 16'h00B5; B = 16'h0097; #100;
A = 16'h00B5; B = 16'h0098; #100;
A = 16'h00B5; B = 16'h0099; #100;
A = 16'h00B5; B = 16'h009A; #100;
A = 16'h00B5; B = 16'h009B; #100;
A = 16'h00B5; B = 16'h009C; #100;
A = 16'h00B5; B = 16'h009D; #100;
A = 16'h00B5; B = 16'h009E; #100;
A = 16'h00B5; B = 16'h009F; #100;
A = 16'h00B5; B = 16'h00A0; #100;
A = 16'h00B5; B = 16'h00A1; #100;
A = 16'h00B5; B = 16'h00A2; #100;
A = 16'h00B5; B = 16'h00A3; #100;
A = 16'h00B5; B = 16'h00A4; #100;
A = 16'h00B5; B = 16'h00A5; #100;
A = 16'h00B5; B = 16'h00A6; #100;
A = 16'h00B5; B = 16'h00A7; #100;
A = 16'h00B5; B = 16'h00A8; #100;
A = 16'h00B5; B = 16'h00A9; #100;
A = 16'h00B5; B = 16'h00AA; #100;
A = 16'h00B5; B = 16'h00AB; #100;
A = 16'h00B5; B = 16'h00AC; #100;
A = 16'h00B5; B = 16'h00AD; #100;
A = 16'h00B5; B = 16'h00AE; #100;
A = 16'h00B5; B = 16'h00AF; #100;
A = 16'h00B5; B = 16'h00B0; #100;
A = 16'h00B5; B = 16'h00B1; #100;
A = 16'h00B5; B = 16'h00B2; #100;
A = 16'h00B5; B = 16'h00B3; #100;
A = 16'h00B5; B = 16'h00B4; #100;
A = 16'h00B5; B = 16'h00B5; #100;
A = 16'h00B5; B = 16'h00B6; #100;
A = 16'h00B5; B = 16'h00B7; #100;
A = 16'h00B5; B = 16'h00B8; #100;
A = 16'h00B5; B = 16'h00B9; #100;
A = 16'h00B5; B = 16'h00BA; #100;
A = 16'h00B5; B = 16'h00BB; #100;
A = 16'h00B5; B = 16'h00BC; #100;
A = 16'h00B5; B = 16'h00BD; #100;
A = 16'h00B5; B = 16'h00BE; #100;
A = 16'h00B5; B = 16'h00BF; #100;
A = 16'h00B5; B = 16'h00C0; #100;
A = 16'h00B5; B = 16'h00C1; #100;
A = 16'h00B5; B = 16'h00C2; #100;
A = 16'h00B5; B = 16'h00C3; #100;
A = 16'h00B5; B = 16'h00C4; #100;
A = 16'h00B5; B = 16'h00C5; #100;
A = 16'h00B5; B = 16'h00C6; #100;
A = 16'h00B5; B = 16'h00C7; #100;
A = 16'h00B5; B = 16'h00C8; #100;
A = 16'h00B5; B = 16'h00C9; #100;
A = 16'h00B5; B = 16'h00CA; #100;
A = 16'h00B5; B = 16'h00CB; #100;
A = 16'h00B5; B = 16'h00CC; #100;
A = 16'h00B5; B = 16'h00CD; #100;
A = 16'h00B5; B = 16'h00CE; #100;
A = 16'h00B5; B = 16'h00CF; #100;
A = 16'h00B5; B = 16'h00D0; #100;
A = 16'h00B5; B = 16'h00D1; #100;
A = 16'h00B5; B = 16'h00D2; #100;
A = 16'h00B5; B = 16'h00D3; #100;
A = 16'h00B5; B = 16'h00D4; #100;
A = 16'h00B5; B = 16'h00D5; #100;
A = 16'h00B5; B = 16'h00D6; #100;
A = 16'h00B5; B = 16'h00D7; #100;
A = 16'h00B5; B = 16'h00D8; #100;
A = 16'h00B5; B = 16'h00D9; #100;
A = 16'h00B5; B = 16'h00DA; #100;
A = 16'h00B5; B = 16'h00DB; #100;
A = 16'h00B5; B = 16'h00DC; #100;
A = 16'h00B5; B = 16'h00DD; #100;
A = 16'h00B5; B = 16'h00DE; #100;
A = 16'h00B5; B = 16'h00DF; #100;
A = 16'h00B5; B = 16'h00E0; #100;
A = 16'h00B5; B = 16'h00E1; #100;
A = 16'h00B5; B = 16'h00E2; #100;
A = 16'h00B5; B = 16'h00E3; #100;
A = 16'h00B5; B = 16'h00E4; #100;
A = 16'h00B5; B = 16'h00E5; #100;
A = 16'h00B5; B = 16'h00E6; #100;
A = 16'h00B5; B = 16'h00E7; #100;
A = 16'h00B5; B = 16'h00E8; #100;
A = 16'h00B5; B = 16'h00E9; #100;
A = 16'h00B5; B = 16'h00EA; #100;
A = 16'h00B5; B = 16'h00EB; #100;
A = 16'h00B5; B = 16'h00EC; #100;
A = 16'h00B5; B = 16'h00ED; #100;
A = 16'h00B5; B = 16'h00EE; #100;
A = 16'h00B5; B = 16'h00EF; #100;
A = 16'h00B5; B = 16'h00F0; #100;
A = 16'h00B5; B = 16'h00F1; #100;
A = 16'h00B5; B = 16'h00F2; #100;
A = 16'h00B5; B = 16'h00F3; #100;
A = 16'h00B5; B = 16'h00F4; #100;
A = 16'h00B5; B = 16'h00F5; #100;
A = 16'h00B5; B = 16'h00F6; #100;
A = 16'h00B5; B = 16'h00F7; #100;
A = 16'h00B5; B = 16'h00F8; #100;
A = 16'h00B5; B = 16'h00F9; #100;
A = 16'h00B5; B = 16'h00FA; #100;
A = 16'h00B5; B = 16'h00FB; #100;
A = 16'h00B5; B = 16'h00FC; #100;
A = 16'h00B5; B = 16'h00FD; #100;
A = 16'h00B5; B = 16'h00FE; #100;
A = 16'h00B5; B = 16'h00FF; #100;
A = 16'h00B6; B = 16'h000; #100;
A = 16'h00B6; B = 16'h001; #100;
A = 16'h00B6; B = 16'h002; #100;
A = 16'h00B6; B = 16'h003; #100;
A = 16'h00B6; B = 16'h004; #100;
A = 16'h00B6; B = 16'h005; #100;
A = 16'h00B6; B = 16'h006; #100;
A = 16'h00B6; B = 16'h007; #100;
A = 16'h00B6; B = 16'h008; #100;
A = 16'h00B6; B = 16'h009; #100;
A = 16'h00B6; B = 16'h00A; #100;
A = 16'h00B6; B = 16'h00B; #100;
A = 16'h00B6; B = 16'h00C; #100;
A = 16'h00B6; B = 16'h00D; #100;
A = 16'h00B6; B = 16'h00E; #100;
A = 16'h00B6; B = 16'h00F; #100;
A = 16'h00B6; B = 16'h0010; #100;
A = 16'h00B6; B = 16'h0011; #100;
A = 16'h00B6; B = 16'h0012; #100;
A = 16'h00B6; B = 16'h0013; #100;
A = 16'h00B6; B = 16'h0014; #100;
A = 16'h00B6; B = 16'h0015; #100;
A = 16'h00B6; B = 16'h0016; #100;
A = 16'h00B6; B = 16'h0017; #100;
A = 16'h00B6; B = 16'h0018; #100;
A = 16'h00B6; B = 16'h0019; #100;
A = 16'h00B6; B = 16'h001A; #100;
A = 16'h00B6; B = 16'h001B; #100;
A = 16'h00B6; B = 16'h001C; #100;
A = 16'h00B6; B = 16'h001D; #100;
A = 16'h00B6; B = 16'h001E; #100;
A = 16'h00B6; B = 16'h001F; #100;
A = 16'h00B6; B = 16'h0020; #100;
A = 16'h00B6; B = 16'h0021; #100;
A = 16'h00B6; B = 16'h0022; #100;
A = 16'h00B6; B = 16'h0023; #100;
A = 16'h00B6; B = 16'h0024; #100;
A = 16'h00B6; B = 16'h0025; #100;
A = 16'h00B6; B = 16'h0026; #100;
A = 16'h00B6; B = 16'h0027; #100;
A = 16'h00B6; B = 16'h0028; #100;
A = 16'h00B6; B = 16'h0029; #100;
A = 16'h00B6; B = 16'h002A; #100;
A = 16'h00B6; B = 16'h002B; #100;
A = 16'h00B6; B = 16'h002C; #100;
A = 16'h00B6; B = 16'h002D; #100;
A = 16'h00B6; B = 16'h002E; #100;
A = 16'h00B6; B = 16'h002F; #100;
A = 16'h00B6; B = 16'h0030; #100;
A = 16'h00B6; B = 16'h0031; #100;
A = 16'h00B6; B = 16'h0032; #100;
A = 16'h00B6; B = 16'h0033; #100;
A = 16'h00B6; B = 16'h0034; #100;
A = 16'h00B6; B = 16'h0035; #100;
A = 16'h00B6; B = 16'h0036; #100;
A = 16'h00B6; B = 16'h0037; #100;
A = 16'h00B6; B = 16'h0038; #100;
A = 16'h00B6; B = 16'h0039; #100;
A = 16'h00B6; B = 16'h003A; #100;
A = 16'h00B6; B = 16'h003B; #100;
A = 16'h00B6; B = 16'h003C; #100;
A = 16'h00B6; B = 16'h003D; #100;
A = 16'h00B6; B = 16'h003E; #100;
A = 16'h00B6; B = 16'h003F; #100;
A = 16'h00B6; B = 16'h0040; #100;
A = 16'h00B6; B = 16'h0041; #100;
A = 16'h00B6; B = 16'h0042; #100;
A = 16'h00B6; B = 16'h0043; #100;
A = 16'h00B6; B = 16'h0044; #100;
A = 16'h00B6; B = 16'h0045; #100;
A = 16'h00B6; B = 16'h0046; #100;
A = 16'h00B6; B = 16'h0047; #100;
A = 16'h00B6; B = 16'h0048; #100;
A = 16'h00B6; B = 16'h0049; #100;
A = 16'h00B6; B = 16'h004A; #100;
A = 16'h00B6; B = 16'h004B; #100;
A = 16'h00B6; B = 16'h004C; #100;
A = 16'h00B6; B = 16'h004D; #100;
A = 16'h00B6; B = 16'h004E; #100;
A = 16'h00B6; B = 16'h004F; #100;
A = 16'h00B6; B = 16'h0050; #100;
A = 16'h00B6; B = 16'h0051; #100;
A = 16'h00B6; B = 16'h0052; #100;
A = 16'h00B6; B = 16'h0053; #100;
A = 16'h00B6; B = 16'h0054; #100;
A = 16'h00B6; B = 16'h0055; #100;
A = 16'h00B6; B = 16'h0056; #100;
A = 16'h00B6; B = 16'h0057; #100;
A = 16'h00B6; B = 16'h0058; #100;
A = 16'h00B6; B = 16'h0059; #100;
A = 16'h00B6; B = 16'h005A; #100;
A = 16'h00B6; B = 16'h005B; #100;
A = 16'h00B6; B = 16'h005C; #100;
A = 16'h00B6; B = 16'h005D; #100;
A = 16'h00B6; B = 16'h005E; #100;
A = 16'h00B6; B = 16'h005F; #100;
A = 16'h00B6; B = 16'h0060; #100;
A = 16'h00B6; B = 16'h0061; #100;
A = 16'h00B6; B = 16'h0062; #100;
A = 16'h00B6; B = 16'h0063; #100;
A = 16'h00B6; B = 16'h0064; #100;
A = 16'h00B6; B = 16'h0065; #100;
A = 16'h00B6; B = 16'h0066; #100;
A = 16'h00B6; B = 16'h0067; #100;
A = 16'h00B6; B = 16'h0068; #100;
A = 16'h00B6; B = 16'h0069; #100;
A = 16'h00B6; B = 16'h006A; #100;
A = 16'h00B6; B = 16'h006B; #100;
A = 16'h00B6; B = 16'h006C; #100;
A = 16'h00B6; B = 16'h006D; #100;
A = 16'h00B6; B = 16'h006E; #100;
A = 16'h00B6; B = 16'h006F; #100;
A = 16'h00B6; B = 16'h0070; #100;
A = 16'h00B6; B = 16'h0071; #100;
A = 16'h00B6; B = 16'h0072; #100;
A = 16'h00B6; B = 16'h0073; #100;
A = 16'h00B6; B = 16'h0074; #100;
A = 16'h00B6; B = 16'h0075; #100;
A = 16'h00B6; B = 16'h0076; #100;
A = 16'h00B6; B = 16'h0077; #100;
A = 16'h00B6; B = 16'h0078; #100;
A = 16'h00B6; B = 16'h0079; #100;
A = 16'h00B6; B = 16'h007A; #100;
A = 16'h00B6; B = 16'h007B; #100;
A = 16'h00B6; B = 16'h007C; #100;
A = 16'h00B6; B = 16'h007D; #100;
A = 16'h00B6; B = 16'h007E; #100;
A = 16'h00B6; B = 16'h007F; #100;
A = 16'h00B6; B = 16'h0080; #100;
A = 16'h00B6; B = 16'h0081; #100;
A = 16'h00B6; B = 16'h0082; #100;
A = 16'h00B6; B = 16'h0083; #100;
A = 16'h00B6; B = 16'h0084; #100;
A = 16'h00B6; B = 16'h0085; #100;
A = 16'h00B6; B = 16'h0086; #100;
A = 16'h00B6; B = 16'h0087; #100;
A = 16'h00B6; B = 16'h0088; #100;
A = 16'h00B6; B = 16'h0089; #100;
A = 16'h00B6; B = 16'h008A; #100;
A = 16'h00B6; B = 16'h008B; #100;
A = 16'h00B6; B = 16'h008C; #100;
A = 16'h00B6; B = 16'h008D; #100;
A = 16'h00B6; B = 16'h008E; #100;
A = 16'h00B6; B = 16'h008F; #100;
A = 16'h00B6; B = 16'h0090; #100;
A = 16'h00B6; B = 16'h0091; #100;
A = 16'h00B6; B = 16'h0092; #100;
A = 16'h00B6; B = 16'h0093; #100;
A = 16'h00B6; B = 16'h0094; #100;
A = 16'h00B6; B = 16'h0095; #100;
A = 16'h00B6; B = 16'h0096; #100;
A = 16'h00B6; B = 16'h0097; #100;
A = 16'h00B6; B = 16'h0098; #100;
A = 16'h00B6; B = 16'h0099; #100;
A = 16'h00B6; B = 16'h009A; #100;
A = 16'h00B6; B = 16'h009B; #100;
A = 16'h00B6; B = 16'h009C; #100;
A = 16'h00B6; B = 16'h009D; #100;
A = 16'h00B6; B = 16'h009E; #100;
A = 16'h00B6; B = 16'h009F; #100;
A = 16'h00B6; B = 16'h00A0; #100;
A = 16'h00B6; B = 16'h00A1; #100;
A = 16'h00B6; B = 16'h00A2; #100;
A = 16'h00B6; B = 16'h00A3; #100;
A = 16'h00B6; B = 16'h00A4; #100;
A = 16'h00B6; B = 16'h00A5; #100;
A = 16'h00B6; B = 16'h00A6; #100;
A = 16'h00B6; B = 16'h00A7; #100;
A = 16'h00B6; B = 16'h00A8; #100;
A = 16'h00B6; B = 16'h00A9; #100;
A = 16'h00B6; B = 16'h00AA; #100;
A = 16'h00B6; B = 16'h00AB; #100;
A = 16'h00B6; B = 16'h00AC; #100;
A = 16'h00B6; B = 16'h00AD; #100;
A = 16'h00B6; B = 16'h00AE; #100;
A = 16'h00B6; B = 16'h00AF; #100;
A = 16'h00B6; B = 16'h00B0; #100;
A = 16'h00B6; B = 16'h00B1; #100;
A = 16'h00B6; B = 16'h00B2; #100;
A = 16'h00B6; B = 16'h00B3; #100;
A = 16'h00B6; B = 16'h00B4; #100;
A = 16'h00B6; B = 16'h00B5; #100;
A = 16'h00B6; B = 16'h00B6; #100;
A = 16'h00B6; B = 16'h00B7; #100;
A = 16'h00B6; B = 16'h00B8; #100;
A = 16'h00B6; B = 16'h00B9; #100;
A = 16'h00B6; B = 16'h00BA; #100;
A = 16'h00B6; B = 16'h00BB; #100;
A = 16'h00B6; B = 16'h00BC; #100;
A = 16'h00B6; B = 16'h00BD; #100;
A = 16'h00B6; B = 16'h00BE; #100;
A = 16'h00B6; B = 16'h00BF; #100;
A = 16'h00B6; B = 16'h00C0; #100;
A = 16'h00B6; B = 16'h00C1; #100;
A = 16'h00B6; B = 16'h00C2; #100;
A = 16'h00B6; B = 16'h00C3; #100;
A = 16'h00B6; B = 16'h00C4; #100;
A = 16'h00B6; B = 16'h00C5; #100;
A = 16'h00B6; B = 16'h00C6; #100;
A = 16'h00B6; B = 16'h00C7; #100;
A = 16'h00B6; B = 16'h00C8; #100;
A = 16'h00B6; B = 16'h00C9; #100;
A = 16'h00B6; B = 16'h00CA; #100;
A = 16'h00B6; B = 16'h00CB; #100;
A = 16'h00B6; B = 16'h00CC; #100;
A = 16'h00B6; B = 16'h00CD; #100;
A = 16'h00B6; B = 16'h00CE; #100;
A = 16'h00B6; B = 16'h00CF; #100;
A = 16'h00B6; B = 16'h00D0; #100;
A = 16'h00B6; B = 16'h00D1; #100;
A = 16'h00B6; B = 16'h00D2; #100;
A = 16'h00B6; B = 16'h00D3; #100;
A = 16'h00B6; B = 16'h00D4; #100;
A = 16'h00B6; B = 16'h00D5; #100;
A = 16'h00B6; B = 16'h00D6; #100;
A = 16'h00B6; B = 16'h00D7; #100;
A = 16'h00B6; B = 16'h00D8; #100;
A = 16'h00B6; B = 16'h00D9; #100;
A = 16'h00B6; B = 16'h00DA; #100;
A = 16'h00B6; B = 16'h00DB; #100;
A = 16'h00B6; B = 16'h00DC; #100;
A = 16'h00B6; B = 16'h00DD; #100;
A = 16'h00B6; B = 16'h00DE; #100;
A = 16'h00B6; B = 16'h00DF; #100;
A = 16'h00B6; B = 16'h00E0; #100;
A = 16'h00B6; B = 16'h00E1; #100;
A = 16'h00B6; B = 16'h00E2; #100;
A = 16'h00B6; B = 16'h00E3; #100;
A = 16'h00B6; B = 16'h00E4; #100;
A = 16'h00B6; B = 16'h00E5; #100;
A = 16'h00B6; B = 16'h00E6; #100;
A = 16'h00B6; B = 16'h00E7; #100;
A = 16'h00B6; B = 16'h00E8; #100;
A = 16'h00B6; B = 16'h00E9; #100;
A = 16'h00B6; B = 16'h00EA; #100;
A = 16'h00B6; B = 16'h00EB; #100;
A = 16'h00B6; B = 16'h00EC; #100;
A = 16'h00B6; B = 16'h00ED; #100;
A = 16'h00B6; B = 16'h00EE; #100;
A = 16'h00B6; B = 16'h00EF; #100;
A = 16'h00B6; B = 16'h00F0; #100;
A = 16'h00B6; B = 16'h00F1; #100;
A = 16'h00B6; B = 16'h00F2; #100;
A = 16'h00B6; B = 16'h00F3; #100;
A = 16'h00B6; B = 16'h00F4; #100;
A = 16'h00B6; B = 16'h00F5; #100;
A = 16'h00B6; B = 16'h00F6; #100;
A = 16'h00B6; B = 16'h00F7; #100;
A = 16'h00B6; B = 16'h00F8; #100;
A = 16'h00B6; B = 16'h00F9; #100;
A = 16'h00B6; B = 16'h00FA; #100;
A = 16'h00B6; B = 16'h00FB; #100;
A = 16'h00B6; B = 16'h00FC; #100;
A = 16'h00B6; B = 16'h00FD; #100;
A = 16'h00B6; B = 16'h00FE; #100;
A = 16'h00B6; B = 16'h00FF; #100;
A = 16'h00B7; B = 16'h000; #100;
A = 16'h00B7; B = 16'h001; #100;
A = 16'h00B7; B = 16'h002; #100;
A = 16'h00B7; B = 16'h003; #100;
A = 16'h00B7; B = 16'h004; #100;
A = 16'h00B7; B = 16'h005; #100;
A = 16'h00B7; B = 16'h006; #100;
A = 16'h00B7; B = 16'h007; #100;
A = 16'h00B7; B = 16'h008; #100;
A = 16'h00B7; B = 16'h009; #100;
A = 16'h00B7; B = 16'h00A; #100;
A = 16'h00B7; B = 16'h00B; #100;
A = 16'h00B7; B = 16'h00C; #100;
A = 16'h00B7; B = 16'h00D; #100;
A = 16'h00B7; B = 16'h00E; #100;
A = 16'h00B7; B = 16'h00F; #100;
A = 16'h00B7; B = 16'h0010; #100;
A = 16'h00B7; B = 16'h0011; #100;
A = 16'h00B7; B = 16'h0012; #100;
A = 16'h00B7; B = 16'h0013; #100;
A = 16'h00B7; B = 16'h0014; #100;
A = 16'h00B7; B = 16'h0015; #100;
A = 16'h00B7; B = 16'h0016; #100;
A = 16'h00B7; B = 16'h0017; #100;
A = 16'h00B7; B = 16'h0018; #100;
A = 16'h00B7; B = 16'h0019; #100;
A = 16'h00B7; B = 16'h001A; #100;
A = 16'h00B7; B = 16'h001B; #100;
A = 16'h00B7; B = 16'h001C; #100;
A = 16'h00B7; B = 16'h001D; #100;
A = 16'h00B7; B = 16'h001E; #100;
A = 16'h00B7; B = 16'h001F; #100;
A = 16'h00B7; B = 16'h0020; #100;
A = 16'h00B7; B = 16'h0021; #100;
A = 16'h00B7; B = 16'h0022; #100;
A = 16'h00B7; B = 16'h0023; #100;
A = 16'h00B7; B = 16'h0024; #100;
A = 16'h00B7; B = 16'h0025; #100;
A = 16'h00B7; B = 16'h0026; #100;
A = 16'h00B7; B = 16'h0027; #100;
A = 16'h00B7; B = 16'h0028; #100;
A = 16'h00B7; B = 16'h0029; #100;
A = 16'h00B7; B = 16'h002A; #100;
A = 16'h00B7; B = 16'h002B; #100;
A = 16'h00B7; B = 16'h002C; #100;
A = 16'h00B7; B = 16'h002D; #100;
A = 16'h00B7; B = 16'h002E; #100;
A = 16'h00B7; B = 16'h002F; #100;
A = 16'h00B7; B = 16'h0030; #100;
A = 16'h00B7; B = 16'h0031; #100;
A = 16'h00B7; B = 16'h0032; #100;
A = 16'h00B7; B = 16'h0033; #100;
A = 16'h00B7; B = 16'h0034; #100;
A = 16'h00B7; B = 16'h0035; #100;
A = 16'h00B7; B = 16'h0036; #100;
A = 16'h00B7; B = 16'h0037; #100;
A = 16'h00B7; B = 16'h0038; #100;
A = 16'h00B7; B = 16'h0039; #100;
A = 16'h00B7; B = 16'h003A; #100;
A = 16'h00B7; B = 16'h003B; #100;
A = 16'h00B7; B = 16'h003C; #100;
A = 16'h00B7; B = 16'h003D; #100;
A = 16'h00B7; B = 16'h003E; #100;
A = 16'h00B7; B = 16'h003F; #100;
A = 16'h00B7; B = 16'h0040; #100;
A = 16'h00B7; B = 16'h0041; #100;
A = 16'h00B7; B = 16'h0042; #100;
A = 16'h00B7; B = 16'h0043; #100;
A = 16'h00B7; B = 16'h0044; #100;
A = 16'h00B7; B = 16'h0045; #100;
A = 16'h00B7; B = 16'h0046; #100;
A = 16'h00B7; B = 16'h0047; #100;
A = 16'h00B7; B = 16'h0048; #100;
A = 16'h00B7; B = 16'h0049; #100;
A = 16'h00B7; B = 16'h004A; #100;
A = 16'h00B7; B = 16'h004B; #100;
A = 16'h00B7; B = 16'h004C; #100;
A = 16'h00B7; B = 16'h004D; #100;
A = 16'h00B7; B = 16'h004E; #100;
A = 16'h00B7; B = 16'h004F; #100;
A = 16'h00B7; B = 16'h0050; #100;
A = 16'h00B7; B = 16'h0051; #100;
A = 16'h00B7; B = 16'h0052; #100;
A = 16'h00B7; B = 16'h0053; #100;
A = 16'h00B7; B = 16'h0054; #100;
A = 16'h00B7; B = 16'h0055; #100;
A = 16'h00B7; B = 16'h0056; #100;
A = 16'h00B7; B = 16'h0057; #100;
A = 16'h00B7; B = 16'h0058; #100;
A = 16'h00B7; B = 16'h0059; #100;
A = 16'h00B7; B = 16'h005A; #100;
A = 16'h00B7; B = 16'h005B; #100;
A = 16'h00B7; B = 16'h005C; #100;
A = 16'h00B7; B = 16'h005D; #100;
A = 16'h00B7; B = 16'h005E; #100;
A = 16'h00B7; B = 16'h005F; #100;
A = 16'h00B7; B = 16'h0060; #100;
A = 16'h00B7; B = 16'h0061; #100;
A = 16'h00B7; B = 16'h0062; #100;
A = 16'h00B7; B = 16'h0063; #100;
A = 16'h00B7; B = 16'h0064; #100;
A = 16'h00B7; B = 16'h0065; #100;
A = 16'h00B7; B = 16'h0066; #100;
A = 16'h00B7; B = 16'h0067; #100;
A = 16'h00B7; B = 16'h0068; #100;
A = 16'h00B7; B = 16'h0069; #100;
A = 16'h00B7; B = 16'h006A; #100;
A = 16'h00B7; B = 16'h006B; #100;
A = 16'h00B7; B = 16'h006C; #100;
A = 16'h00B7; B = 16'h006D; #100;
A = 16'h00B7; B = 16'h006E; #100;
A = 16'h00B7; B = 16'h006F; #100;
A = 16'h00B7; B = 16'h0070; #100;
A = 16'h00B7; B = 16'h0071; #100;
A = 16'h00B7; B = 16'h0072; #100;
A = 16'h00B7; B = 16'h0073; #100;
A = 16'h00B7; B = 16'h0074; #100;
A = 16'h00B7; B = 16'h0075; #100;
A = 16'h00B7; B = 16'h0076; #100;
A = 16'h00B7; B = 16'h0077; #100;
A = 16'h00B7; B = 16'h0078; #100;
A = 16'h00B7; B = 16'h0079; #100;
A = 16'h00B7; B = 16'h007A; #100;
A = 16'h00B7; B = 16'h007B; #100;
A = 16'h00B7; B = 16'h007C; #100;
A = 16'h00B7; B = 16'h007D; #100;
A = 16'h00B7; B = 16'h007E; #100;
A = 16'h00B7; B = 16'h007F; #100;
A = 16'h00B7; B = 16'h0080; #100;
A = 16'h00B7; B = 16'h0081; #100;
A = 16'h00B7; B = 16'h0082; #100;
A = 16'h00B7; B = 16'h0083; #100;
A = 16'h00B7; B = 16'h0084; #100;
A = 16'h00B7; B = 16'h0085; #100;
A = 16'h00B7; B = 16'h0086; #100;
A = 16'h00B7; B = 16'h0087; #100;
A = 16'h00B7; B = 16'h0088; #100;
A = 16'h00B7; B = 16'h0089; #100;
A = 16'h00B7; B = 16'h008A; #100;
A = 16'h00B7; B = 16'h008B; #100;
A = 16'h00B7; B = 16'h008C; #100;
A = 16'h00B7; B = 16'h008D; #100;
A = 16'h00B7; B = 16'h008E; #100;
A = 16'h00B7; B = 16'h008F; #100;
A = 16'h00B7; B = 16'h0090; #100;
A = 16'h00B7; B = 16'h0091; #100;
A = 16'h00B7; B = 16'h0092; #100;
A = 16'h00B7; B = 16'h0093; #100;
A = 16'h00B7; B = 16'h0094; #100;
A = 16'h00B7; B = 16'h0095; #100;
A = 16'h00B7; B = 16'h0096; #100;
A = 16'h00B7; B = 16'h0097; #100;
A = 16'h00B7; B = 16'h0098; #100;
A = 16'h00B7; B = 16'h0099; #100;
A = 16'h00B7; B = 16'h009A; #100;
A = 16'h00B7; B = 16'h009B; #100;
A = 16'h00B7; B = 16'h009C; #100;
A = 16'h00B7; B = 16'h009D; #100;
A = 16'h00B7; B = 16'h009E; #100;
A = 16'h00B7; B = 16'h009F; #100;
A = 16'h00B7; B = 16'h00A0; #100;
A = 16'h00B7; B = 16'h00A1; #100;
A = 16'h00B7; B = 16'h00A2; #100;
A = 16'h00B7; B = 16'h00A3; #100;
A = 16'h00B7; B = 16'h00A4; #100;
A = 16'h00B7; B = 16'h00A5; #100;
A = 16'h00B7; B = 16'h00A6; #100;
A = 16'h00B7; B = 16'h00A7; #100;
A = 16'h00B7; B = 16'h00A8; #100;
A = 16'h00B7; B = 16'h00A9; #100;
A = 16'h00B7; B = 16'h00AA; #100;
A = 16'h00B7; B = 16'h00AB; #100;
A = 16'h00B7; B = 16'h00AC; #100;
A = 16'h00B7; B = 16'h00AD; #100;
A = 16'h00B7; B = 16'h00AE; #100;
A = 16'h00B7; B = 16'h00AF; #100;
A = 16'h00B7; B = 16'h00B0; #100;
A = 16'h00B7; B = 16'h00B1; #100;
A = 16'h00B7; B = 16'h00B2; #100;
A = 16'h00B7; B = 16'h00B3; #100;
A = 16'h00B7; B = 16'h00B4; #100;
A = 16'h00B7; B = 16'h00B5; #100;
A = 16'h00B7; B = 16'h00B6; #100;
A = 16'h00B7; B = 16'h00B7; #100;
A = 16'h00B7; B = 16'h00B8; #100;
A = 16'h00B7; B = 16'h00B9; #100;
A = 16'h00B7; B = 16'h00BA; #100;
A = 16'h00B7; B = 16'h00BB; #100;
A = 16'h00B7; B = 16'h00BC; #100;
A = 16'h00B7; B = 16'h00BD; #100;
A = 16'h00B7; B = 16'h00BE; #100;
A = 16'h00B7; B = 16'h00BF; #100;
A = 16'h00B7; B = 16'h00C0; #100;
A = 16'h00B7; B = 16'h00C1; #100;
A = 16'h00B7; B = 16'h00C2; #100;
A = 16'h00B7; B = 16'h00C3; #100;
A = 16'h00B7; B = 16'h00C4; #100;
A = 16'h00B7; B = 16'h00C5; #100;
A = 16'h00B7; B = 16'h00C6; #100;
A = 16'h00B7; B = 16'h00C7; #100;
A = 16'h00B7; B = 16'h00C8; #100;
A = 16'h00B7; B = 16'h00C9; #100;
A = 16'h00B7; B = 16'h00CA; #100;
A = 16'h00B7; B = 16'h00CB; #100;
A = 16'h00B7; B = 16'h00CC; #100;
A = 16'h00B7; B = 16'h00CD; #100;
A = 16'h00B7; B = 16'h00CE; #100;
A = 16'h00B7; B = 16'h00CF; #100;
A = 16'h00B7; B = 16'h00D0; #100;
A = 16'h00B7; B = 16'h00D1; #100;
A = 16'h00B7; B = 16'h00D2; #100;
A = 16'h00B7; B = 16'h00D3; #100;
A = 16'h00B7; B = 16'h00D4; #100;
A = 16'h00B7; B = 16'h00D5; #100;
A = 16'h00B7; B = 16'h00D6; #100;
A = 16'h00B7; B = 16'h00D7; #100;
A = 16'h00B7; B = 16'h00D8; #100;
A = 16'h00B7; B = 16'h00D9; #100;
A = 16'h00B7; B = 16'h00DA; #100;
A = 16'h00B7; B = 16'h00DB; #100;
A = 16'h00B7; B = 16'h00DC; #100;
A = 16'h00B7; B = 16'h00DD; #100;
A = 16'h00B7; B = 16'h00DE; #100;
A = 16'h00B7; B = 16'h00DF; #100;
A = 16'h00B7; B = 16'h00E0; #100;
A = 16'h00B7; B = 16'h00E1; #100;
A = 16'h00B7; B = 16'h00E2; #100;
A = 16'h00B7; B = 16'h00E3; #100;
A = 16'h00B7; B = 16'h00E4; #100;
A = 16'h00B7; B = 16'h00E5; #100;
A = 16'h00B7; B = 16'h00E6; #100;
A = 16'h00B7; B = 16'h00E7; #100;
A = 16'h00B7; B = 16'h00E8; #100;
A = 16'h00B7; B = 16'h00E9; #100;
A = 16'h00B7; B = 16'h00EA; #100;
A = 16'h00B7; B = 16'h00EB; #100;
A = 16'h00B7; B = 16'h00EC; #100;
A = 16'h00B7; B = 16'h00ED; #100;
A = 16'h00B7; B = 16'h00EE; #100;
A = 16'h00B7; B = 16'h00EF; #100;
A = 16'h00B7; B = 16'h00F0; #100;
A = 16'h00B7; B = 16'h00F1; #100;
A = 16'h00B7; B = 16'h00F2; #100;
A = 16'h00B7; B = 16'h00F3; #100;
A = 16'h00B7; B = 16'h00F4; #100;
A = 16'h00B7; B = 16'h00F5; #100;
A = 16'h00B7; B = 16'h00F6; #100;
A = 16'h00B7; B = 16'h00F7; #100;
A = 16'h00B7; B = 16'h00F8; #100;
A = 16'h00B7; B = 16'h00F9; #100;
A = 16'h00B7; B = 16'h00FA; #100;
A = 16'h00B7; B = 16'h00FB; #100;
A = 16'h00B7; B = 16'h00FC; #100;
A = 16'h00B7; B = 16'h00FD; #100;
A = 16'h00B7; B = 16'h00FE; #100;
A = 16'h00B7; B = 16'h00FF; #100;
A = 16'h00B8; B = 16'h000; #100;
A = 16'h00B8; B = 16'h001; #100;
A = 16'h00B8; B = 16'h002; #100;
A = 16'h00B8; B = 16'h003; #100;
A = 16'h00B8; B = 16'h004; #100;
A = 16'h00B8; B = 16'h005; #100;
A = 16'h00B8; B = 16'h006; #100;
A = 16'h00B8; B = 16'h007; #100;
A = 16'h00B8; B = 16'h008; #100;
A = 16'h00B8; B = 16'h009; #100;
A = 16'h00B8; B = 16'h00A; #100;
A = 16'h00B8; B = 16'h00B; #100;
A = 16'h00B8; B = 16'h00C; #100;
A = 16'h00B8; B = 16'h00D; #100;
A = 16'h00B8; B = 16'h00E; #100;
A = 16'h00B8; B = 16'h00F; #100;
A = 16'h00B8; B = 16'h0010; #100;
A = 16'h00B8; B = 16'h0011; #100;
A = 16'h00B8; B = 16'h0012; #100;
A = 16'h00B8; B = 16'h0013; #100;
A = 16'h00B8; B = 16'h0014; #100;
A = 16'h00B8; B = 16'h0015; #100;
A = 16'h00B8; B = 16'h0016; #100;
A = 16'h00B8; B = 16'h0017; #100;
A = 16'h00B8; B = 16'h0018; #100;
A = 16'h00B8; B = 16'h0019; #100;
A = 16'h00B8; B = 16'h001A; #100;
A = 16'h00B8; B = 16'h001B; #100;
A = 16'h00B8; B = 16'h001C; #100;
A = 16'h00B8; B = 16'h001D; #100;
A = 16'h00B8; B = 16'h001E; #100;
A = 16'h00B8; B = 16'h001F; #100;
A = 16'h00B8; B = 16'h0020; #100;
A = 16'h00B8; B = 16'h0021; #100;
A = 16'h00B8; B = 16'h0022; #100;
A = 16'h00B8; B = 16'h0023; #100;
A = 16'h00B8; B = 16'h0024; #100;
A = 16'h00B8; B = 16'h0025; #100;
A = 16'h00B8; B = 16'h0026; #100;
A = 16'h00B8; B = 16'h0027; #100;
A = 16'h00B8; B = 16'h0028; #100;
A = 16'h00B8; B = 16'h0029; #100;
A = 16'h00B8; B = 16'h002A; #100;
A = 16'h00B8; B = 16'h002B; #100;
A = 16'h00B8; B = 16'h002C; #100;
A = 16'h00B8; B = 16'h002D; #100;
A = 16'h00B8; B = 16'h002E; #100;
A = 16'h00B8; B = 16'h002F; #100;
A = 16'h00B8; B = 16'h0030; #100;
A = 16'h00B8; B = 16'h0031; #100;
A = 16'h00B8; B = 16'h0032; #100;
A = 16'h00B8; B = 16'h0033; #100;
A = 16'h00B8; B = 16'h0034; #100;
A = 16'h00B8; B = 16'h0035; #100;
A = 16'h00B8; B = 16'h0036; #100;
A = 16'h00B8; B = 16'h0037; #100;
A = 16'h00B8; B = 16'h0038; #100;
A = 16'h00B8; B = 16'h0039; #100;
A = 16'h00B8; B = 16'h003A; #100;
A = 16'h00B8; B = 16'h003B; #100;
A = 16'h00B8; B = 16'h003C; #100;
A = 16'h00B8; B = 16'h003D; #100;
A = 16'h00B8; B = 16'h003E; #100;
A = 16'h00B8; B = 16'h003F; #100;
A = 16'h00B8; B = 16'h0040; #100;
A = 16'h00B8; B = 16'h0041; #100;
A = 16'h00B8; B = 16'h0042; #100;
A = 16'h00B8; B = 16'h0043; #100;
A = 16'h00B8; B = 16'h0044; #100;
A = 16'h00B8; B = 16'h0045; #100;
A = 16'h00B8; B = 16'h0046; #100;
A = 16'h00B8; B = 16'h0047; #100;
A = 16'h00B8; B = 16'h0048; #100;
A = 16'h00B8; B = 16'h0049; #100;
A = 16'h00B8; B = 16'h004A; #100;
A = 16'h00B8; B = 16'h004B; #100;
A = 16'h00B8; B = 16'h004C; #100;
A = 16'h00B8; B = 16'h004D; #100;
A = 16'h00B8; B = 16'h004E; #100;
A = 16'h00B8; B = 16'h004F; #100;
A = 16'h00B8; B = 16'h0050; #100;
A = 16'h00B8; B = 16'h0051; #100;
A = 16'h00B8; B = 16'h0052; #100;
A = 16'h00B8; B = 16'h0053; #100;
A = 16'h00B8; B = 16'h0054; #100;
A = 16'h00B8; B = 16'h0055; #100;
A = 16'h00B8; B = 16'h0056; #100;
A = 16'h00B8; B = 16'h0057; #100;
A = 16'h00B8; B = 16'h0058; #100;
A = 16'h00B8; B = 16'h0059; #100;
A = 16'h00B8; B = 16'h005A; #100;
A = 16'h00B8; B = 16'h005B; #100;
A = 16'h00B8; B = 16'h005C; #100;
A = 16'h00B8; B = 16'h005D; #100;
A = 16'h00B8; B = 16'h005E; #100;
A = 16'h00B8; B = 16'h005F; #100;
A = 16'h00B8; B = 16'h0060; #100;
A = 16'h00B8; B = 16'h0061; #100;
A = 16'h00B8; B = 16'h0062; #100;
A = 16'h00B8; B = 16'h0063; #100;
A = 16'h00B8; B = 16'h0064; #100;
A = 16'h00B8; B = 16'h0065; #100;
A = 16'h00B8; B = 16'h0066; #100;
A = 16'h00B8; B = 16'h0067; #100;
A = 16'h00B8; B = 16'h0068; #100;
A = 16'h00B8; B = 16'h0069; #100;
A = 16'h00B8; B = 16'h006A; #100;
A = 16'h00B8; B = 16'h006B; #100;
A = 16'h00B8; B = 16'h006C; #100;
A = 16'h00B8; B = 16'h006D; #100;
A = 16'h00B8; B = 16'h006E; #100;
A = 16'h00B8; B = 16'h006F; #100;
A = 16'h00B8; B = 16'h0070; #100;
A = 16'h00B8; B = 16'h0071; #100;
A = 16'h00B8; B = 16'h0072; #100;
A = 16'h00B8; B = 16'h0073; #100;
A = 16'h00B8; B = 16'h0074; #100;
A = 16'h00B8; B = 16'h0075; #100;
A = 16'h00B8; B = 16'h0076; #100;
A = 16'h00B8; B = 16'h0077; #100;
A = 16'h00B8; B = 16'h0078; #100;
A = 16'h00B8; B = 16'h0079; #100;
A = 16'h00B8; B = 16'h007A; #100;
A = 16'h00B8; B = 16'h007B; #100;
A = 16'h00B8; B = 16'h007C; #100;
A = 16'h00B8; B = 16'h007D; #100;
A = 16'h00B8; B = 16'h007E; #100;
A = 16'h00B8; B = 16'h007F; #100;
A = 16'h00B8; B = 16'h0080; #100;
A = 16'h00B8; B = 16'h0081; #100;
A = 16'h00B8; B = 16'h0082; #100;
A = 16'h00B8; B = 16'h0083; #100;
A = 16'h00B8; B = 16'h0084; #100;
A = 16'h00B8; B = 16'h0085; #100;
A = 16'h00B8; B = 16'h0086; #100;
A = 16'h00B8; B = 16'h0087; #100;
A = 16'h00B8; B = 16'h0088; #100;
A = 16'h00B8; B = 16'h0089; #100;
A = 16'h00B8; B = 16'h008A; #100;
A = 16'h00B8; B = 16'h008B; #100;
A = 16'h00B8; B = 16'h008C; #100;
A = 16'h00B8; B = 16'h008D; #100;
A = 16'h00B8; B = 16'h008E; #100;
A = 16'h00B8; B = 16'h008F; #100;
A = 16'h00B8; B = 16'h0090; #100;
A = 16'h00B8; B = 16'h0091; #100;
A = 16'h00B8; B = 16'h0092; #100;
A = 16'h00B8; B = 16'h0093; #100;
A = 16'h00B8; B = 16'h0094; #100;
A = 16'h00B8; B = 16'h0095; #100;
A = 16'h00B8; B = 16'h0096; #100;
A = 16'h00B8; B = 16'h0097; #100;
A = 16'h00B8; B = 16'h0098; #100;
A = 16'h00B8; B = 16'h0099; #100;
A = 16'h00B8; B = 16'h009A; #100;
A = 16'h00B8; B = 16'h009B; #100;
A = 16'h00B8; B = 16'h009C; #100;
A = 16'h00B8; B = 16'h009D; #100;
A = 16'h00B8; B = 16'h009E; #100;
A = 16'h00B8; B = 16'h009F; #100;
A = 16'h00B8; B = 16'h00A0; #100;
A = 16'h00B8; B = 16'h00A1; #100;
A = 16'h00B8; B = 16'h00A2; #100;
A = 16'h00B8; B = 16'h00A3; #100;
A = 16'h00B8; B = 16'h00A4; #100;
A = 16'h00B8; B = 16'h00A5; #100;
A = 16'h00B8; B = 16'h00A6; #100;
A = 16'h00B8; B = 16'h00A7; #100;
A = 16'h00B8; B = 16'h00A8; #100;
A = 16'h00B8; B = 16'h00A9; #100;
A = 16'h00B8; B = 16'h00AA; #100;
A = 16'h00B8; B = 16'h00AB; #100;
A = 16'h00B8; B = 16'h00AC; #100;
A = 16'h00B8; B = 16'h00AD; #100;
A = 16'h00B8; B = 16'h00AE; #100;
A = 16'h00B8; B = 16'h00AF; #100;
A = 16'h00B8; B = 16'h00B0; #100;
A = 16'h00B8; B = 16'h00B1; #100;
A = 16'h00B8; B = 16'h00B2; #100;
A = 16'h00B8; B = 16'h00B3; #100;
A = 16'h00B8; B = 16'h00B4; #100;
A = 16'h00B8; B = 16'h00B5; #100;
A = 16'h00B8; B = 16'h00B6; #100;
A = 16'h00B8; B = 16'h00B7; #100;
A = 16'h00B8; B = 16'h00B8; #100;
A = 16'h00B8; B = 16'h00B9; #100;
A = 16'h00B8; B = 16'h00BA; #100;
A = 16'h00B8; B = 16'h00BB; #100;
A = 16'h00B8; B = 16'h00BC; #100;
A = 16'h00B8; B = 16'h00BD; #100;
A = 16'h00B8; B = 16'h00BE; #100;
A = 16'h00B8; B = 16'h00BF; #100;
A = 16'h00B8; B = 16'h00C0; #100;
A = 16'h00B8; B = 16'h00C1; #100;
A = 16'h00B8; B = 16'h00C2; #100;
A = 16'h00B8; B = 16'h00C3; #100;
A = 16'h00B8; B = 16'h00C4; #100;
A = 16'h00B8; B = 16'h00C5; #100;
A = 16'h00B8; B = 16'h00C6; #100;
A = 16'h00B8; B = 16'h00C7; #100;
A = 16'h00B8; B = 16'h00C8; #100;
A = 16'h00B8; B = 16'h00C9; #100;
A = 16'h00B8; B = 16'h00CA; #100;
A = 16'h00B8; B = 16'h00CB; #100;
A = 16'h00B8; B = 16'h00CC; #100;
A = 16'h00B8; B = 16'h00CD; #100;
A = 16'h00B8; B = 16'h00CE; #100;
A = 16'h00B8; B = 16'h00CF; #100;
A = 16'h00B8; B = 16'h00D0; #100;
A = 16'h00B8; B = 16'h00D1; #100;
A = 16'h00B8; B = 16'h00D2; #100;
A = 16'h00B8; B = 16'h00D3; #100;
A = 16'h00B8; B = 16'h00D4; #100;
A = 16'h00B8; B = 16'h00D5; #100;
A = 16'h00B8; B = 16'h00D6; #100;
A = 16'h00B8; B = 16'h00D7; #100;
A = 16'h00B8; B = 16'h00D8; #100;
A = 16'h00B8; B = 16'h00D9; #100;
A = 16'h00B8; B = 16'h00DA; #100;
A = 16'h00B8; B = 16'h00DB; #100;
A = 16'h00B8; B = 16'h00DC; #100;
A = 16'h00B8; B = 16'h00DD; #100;
A = 16'h00B8; B = 16'h00DE; #100;
A = 16'h00B8; B = 16'h00DF; #100;
A = 16'h00B8; B = 16'h00E0; #100;
A = 16'h00B8; B = 16'h00E1; #100;
A = 16'h00B8; B = 16'h00E2; #100;
A = 16'h00B8; B = 16'h00E3; #100;
A = 16'h00B8; B = 16'h00E4; #100;
A = 16'h00B8; B = 16'h00E5; #100;
A = 16'h00B8; B = 16'h00E6; #100;
A = 16'h00B8; B = 16'h00E7; #100;
A = 16'h00B8; B = 16'h00E8; #100;
A = 16'h00B8; B = 16'h00E9; #100;
A = 16'h00B8; B = 16'h00EA; #100;
A = 16'h00B8; B = 16'h00EB; #100;
A = 16'h00B8; B = 16'h00EC; #100;
A = 16'h00B8; B = 16'h00ED; #100;
A = 16'h00B8; B = 16'h00EE; #100;
A = 16'h00B8; B = 16'h00EF; #100;
A = 16'h00B8; B = 16'h00F0; #100;
A = 16'h00B8; B = 16'h00F1; #100;
A = 16'h00B8; B = 16'h00F2; #100;
A = 16'h00B8; B = 16'h00F3; #100;
A = 16'h00B8; B = 16'h00F4; #100;
A = 16'h00B8; B = 16'h00F5; #100;
A = 16'h00B8; B = 16'h00F6; #100;
A = 16'h00B8; B = 16'h00F7; #100;
A = 16'h00B8; B = 16'h00F8; #100;
A = 16'h00B8; B = 16'h00F9; #100;
A = 16'h00B8; B = 16'h00FA; #100;
A = 16'h00B8; B = 16'h00FB; #100;
A = 16'h00B8; B = 16'h00FC; #100;
A = 16'h00B8; B = 16'h00FD; #100;
A = 16'h00B8; B = 16'h00FE; #100;
A = 16'h00B8; B = 16'h00FF; #100;
A = 16'h00B9; B = 16'h000; #100;
A = 16'h00B9; B = 16'h001; #100;
A = 16'h00B9; B = 16'h002; #100;
A = 16'h00B9; B = 16'h003; #100;
A = 16'h00B9; B = 16'h004; #100;
A = 16'h00B9; B = 16'h005; #100;
A = 16'h00B9; B = 16'h006; #100;
A = 16'h00B9; B = 16'h007; #100;
A = 16'h00B9; B = 16'h008; #100;
A = 16'h00B9; B = 16'h009; #100;
A = 16'h00B9; B = 16'h00A; #100;
A = 16'h00B9; B = 16'h00B; #100;
A = 16'h00B9; B = 16'h00C; #100;
A = 16'h00B9; B = 16'h00D; #100;
A = 16'h00B9; B = 16'h00E; #100;
A = 16'h00B9; B = 16'h00F; #100;
A = 16'h00B9; B = 16'h0010; #100;
A = 16'h00B9; B = 16'h0011; #100;
A = 16'h00B9; B = 16'h0012; #100;
A = 16'h00B9; B = 16'h0013; #100;
A = 16'h00B9; B = 16'h0014; #100;
A = 16'h00B9; B = 16'h0015; #100;
A = 16'h00B9; B = 16'h0016; #100;
A = 16'h00B9; B = 16'h0017; #100;
A = 16'h00B9; B = 16'h0018; #100;
A = 16'h00B9; B = 16'h0019; #100;
A = 16'h00B9; B = 16'h001A; #100;
A = 16'h00B9; B = 16'h001B; #100;
A = 16'h00B9; B = 16'h001C; #100;
A = 16'h00B9; B = 16'h001D; #100;
A = 16'h00B9; B = 16'h001E; #100;
A = 16'h00B9; B = 16'h001F; #100;
A = 16'h00B9; B = 16'h0020; #100;
A = 16'h00B9; B = 16'h0021; #100;
A = 16'h00B9; B = 16'h0022; #100;
A = 16'h00B9; B = 16'h0023; #100;
A = 16'h00B9; B = 16'h0024; #100;
A = 16'h00B9; B = 16'h0025; #100;
A = 16'h00B9; B = 16'h0026; #100;
A = 16'h00B9; B = 16'h0027; #100;
A = 16'h00B9; B = 16'h0028; #100;
A = 16'h00B9; B = 16'h0029; #100;
A = 16'h00B9; B = 16'h002A; #100;
A = 16'h00B9; B = 16'h002B; #100;
A = 16'h00B9; B = 16'h002C; #100;
A = 16'h00B9; B = 16'h002D; #100;
A = 16'h00B9; B = 16'h002E; #100;
A = 16'h00B9; B = 16'h002F; #100;
A = 16'h00B9; B = 16'h0030; #100;
A = 16'h00B9; B = 16'h0031; #100;
A = 16'h00B9; B = 16'h0032; #100;
A = 16'h00B9; B = 16'h0033; #100;
A = 16'h00B9; B = 16'h0034; #100;
A = 16'h00B9; B = 16'h0035; #100;
A = 16'h00B9; B = 16'h0036; #100;
A = 16'h00B9; B = 16'h0037; #100;
A = 16'h00B9; B = 16'h0038; #100;
A = 16'h00B9; B = 16'h0039; #100;
A = 16'h00B9; B = 16'h003A; #100;
A = 16'h00B9; B = 16'h003B; #100;
A = 16'h00B9; B = 16'h003C; #100;
A = 16'h00B9; B = 16'h003D; #100;
A = 16'h00B9; B = 16'h003E; #100;
A = 16'h00B9; B = 16'h003F; #100;
A = 16'h00B9; B = 16'h0040; #100;
A = 16'h00B9; B = 16'h0041; #100;
A = 16'h00B9; B = 16'h0042; #100;
A = 16'h00B9; B = 16'h0043; #100;
A = 16'h00B9; B = 16'h0044; #100;
A = 16'h00B9; B = 16'h0045; #100;
A = 16'h00B9; B = 16'h0046; #100;
A = 16'h00B9; B = 16'h0047; #100;
A = 16'h00B9; B = 16'h0048; #100;
A = 16'h00B9; B = 16'h0049; #100;
A = 16'h00B9; B = 16'h004A; #100;
A = 16'h00B9; B = 16'h004B; #100;
A = 16'h00B9; B = 16'h004C; #100;
A = 16'h00B9; B = 16'h004D; #100;
A = 16'h00B9; B = 16'h004E; #100;
A = 16'h00B9; B = 16'h004F; #100;
A = 16'h00B9; B = 16'h0050; #100;
A = 16'h00B9; B = 16'h0051; #100;
A = 16'h00B9; B = 16'h0052; #100;
A = 16'h00B9; B = 16'h0053; #100;
A = 16'h00B9; B = 16'h0054; #100;
A = 16'h00B9; B = 16'h0055; #100;
A = 16'h00B9; B = 16'h0056; #100;
A = 16'h00B9; B = 16'h0057; #100;
A = 16'h00B9; B = 16'h0058; #100;
A = 16'h00B9; B = 16'h0059; #100;
A = 16'h00B9; B = 16'h005A; #100;
A = 16'h00B9; B = 16'h005B; #100;
A = 16'h00B9; B = 16'h005C; #100;
A = 16'h00B9; B = 16'h005D; #100;
A = 16'h00B9; B = 16'h005E; #100;
A = 16'h00B9; B = 16'h005F; #100;
A = 16'h00B9; B = 16'h0060; #100;
A = 16'h00B9; B = 16'h0061; #100;
A = 16'h00B9; B = 16'h0062; #100;
A = 16'h00B9; B = 16'h0063; #100;
A = 16'h00B9; B = 16'h0064; #100;
A = 16'h00B9; B = 16'h0065; #100;
A = 16'h00B9; B = 16'h0066; #100;
A = 16'h00B9; B = 16'h0067; #100;
A = 16'h00B9; B = 16'h0068; #100;
A = 16'h00B9; B = 16'h0069; #100;
A = 16'h00B9; B = 16'h006A; #100;
A = 16'h00B9; B = 16'h006B; #100;
A = 16'h00B9; B = 16'h006C; #100;
A = 16'h00B9; B = 16'h006D; #100;
A = 16'h00B9; B = 16'h006E; #100;
A = 16'h00B9; B = 16'h006F; #100;
A = 16'h00B9; B = 16'h0070; #100;
A = 16'h00B9; B = 16'h0071; #100;
A = 16'h00B9; B = 16'h0072; #100;
A = 16'h00B9; B = 16'h0073; #100;
A = 16'h00B9; B = 16'h0074; #100;
A = 16'h00B9; B = 16'h0075; #100;
A = 16'h00B9; B = 16'h0076; #100;
A = 16'h00B9; B = 16'h0077; #100;
A = 16'h00B9; B = 16'h0078; #100;
A = 16'h00B9; B = 16'h0079; #100;
A = 16'h00B9; B = 16'h007A; #100;
A = 16'h00B9; B = 16'h007B; #100;
A = 16'h00B9; B = 16'h007C; #100;
A = 16'h00B9; B = 16'h007D; #100;
A = 16'h00B9; B = 16'h007E; #100;
A = 16'h00B9; B = 16'h007F; #100;
A = 16'h00B9; B = 16'h0080; #100;
A = 16'h00B9; B = 16'h0081; #100;
A = 16'h00B9; B = 16'h0082; #100;
A = 16'h00B9; B = 16'h0083; #100;
A = 16'h00B9; B = 16'h0084; #100;
A = 16'h00B9; B = 16'h0085; #100;
A = 16'h00B9; B = 16'h0086; #100;
A = 16'h00B9; B = 16'h0087; #100;
A = 16'h00B9; B = 16'h0088; #100;
A = 16'h00B9; B = 16'h0089; #100;
A = 16'h00B9; B = 16'h008A; #100;
A = 16'h00B9; B = 16'h008B; #100;
A = 16'h00B9; B = 16'h008C; #100;
A = 16'h00B9; B = 16'h008D; #100;
A = 16'h00B9; B = 16'h008E; #100;
A = 16'h00B9; B = 16'h008F; #100;
A = 16'h00B9; B = 16'h0090; #100;
A = 16'h00B9; B = 16'h0091; #100;
A = 16'h00B9; B = 16'h0092; #100;
A = 16'h00B9; B = 16'h0093; #100;
A = 16'h00B9; B = 16'h0094; #100;
A = 16'h00B9; B = 16'h0095; #100;
A = 16'h00B9; B = 16'h0096; #100;
A = 16'h00B9; B = 16'h0097; #100;
A = 16'h00B9; B = 16'h0098; #100;
A = 16'h00B9; B = 16'h0099; #100;
A = 16'h00B9; B = 16'h009A; #100;
A = 16'h00B9; B = 16'h009B; #100;
A = 16'h00B9; B = 16'h009C; #100;
A = 16'h00B9; B = 16'h009D; #100;
A = 16'h00B9; B = 16'h009E; #100;
A = 16'h00B9; B = 16'h009F; #100;
A = 16'h00B9; B = 16'h00A0; #100;
A = 16'h00B9; B = 16'h00A1; #100;
A = 16'h00B9; B = 16'h00A2; #100;
A = 16'h00B9; B = 16'h00A3; #100;
A = 16'h00B9; B = 16'h00A4; #100;
A = 16'h00B9; B = 16'h00A5; #100;
A = 16'h00B9; B = 16'h00A6; #100;
A = 16'h00B9; B = 16'h00A7; #100;
A = 16'h00B9; B = 16'h00A8; #100;
A = 16'h00B9; B = 16'h00A9; #100;
A = 16'h00B9; B = 16'h00AA; #100;
A = 16'h00B9; B = 16'h00AB; #100;
A = 16'h00B9; B = 16'h00AC; #100;
A = 16'h00B9; B = 16'h00AD; #100;
A = 16'h00B9; B = 16'h00AE; #100;
A = 16'h00B9; B = 16'h00AF; #100;
A = 16'h00B9; B = 16'h00B0; #100;
A = 16'h00B9; B = 16'h00B1; #100;
A = 16'h00B9; B = 16'h00B2; #100;
A = 16'h00B9; B = 16'h00B3; #100;
A = 16'h00B9; B = 16'h00B4; #100;
A = 16'h00B9; B = 16'h00B5; #100;
A = 16'h00B9; B = 16'h00B6; #100;
A = 16'h00B9; B = 16'h00B7; #100;
A = 16'h00B9; B = 16'h00B8; #100;
A = 16'h00B9; B = 16'h00B9; #100;
A = 16'h00B9; B = 16'h00BA; #100;
A = 16'h00B9; B = 16'h00BB; #100;
A = 16'h00B9; B = 16'h00BC; #100;
A = 16'h00B9; B = 16'h00BD; #100;
A = 16'h00B9; B = 16'h00BE; #100;
A = 16'h00B9; B = 16'h00BF; #100;
A = 16'h00B9; B = 16'h00C0; #100;
A = 16'h00B9; B = 16'h00C1; #100;
A = 16'h00B9; B = 16'h00C2; #100;
A = 16'h00B9; B = 16'h00C3; #100;
A = 16'h00B9; B = 16'h00C4; #100;
A = 16'h00B9; B = 16'h00C5; #100;
A = 16'h00B9; B = 16'h00C6; #100;
A = 16'h00B9; B = 16'h00C7; #100;
A = 16'h00B9; B = 16'h00C8; #100;
A = 16'h00B9; B = 16'h00C9; #100;
A = 16'h00B9; B = 16'h00CA; #100;
A = 16'h00B9; B = 16'h00CB; #100;
A = 16'h00B9; B = 16'h00CC; #100;
A = 16'h00B9; B = 16'h00CD; #100;
A = 16'h00B9; B = 16'h00CE; #100;
A = 16'h00B9; B = 16'h00CF; #100;
A = 16'h00B9; B = 16'h00D0; #100;
A = 16'h00B9; B = 16'h00D1; #100;
A = 16'h00B9; B = 16'h00D2; #100;
A = 16'h00B9; B = 16'h00D3; #100;
A = 16'h00B9; B = 16'h00D4; #100;
A = 16'h00B9; B = 16'h00D5; #100;
A = 16'h00B9; B = 16'h00D6; #100;
A = 16'h00B9; B = 16'h00D7; #100;
A = 16'h00B9; B = 16'h00D8; #100;
A = 16'h00B9; B = 16'h00D9; #100;
A = 16'h00B9; B = 16'h00DA; #100;
A = 16'h00B9; B = 16'h00DB; #100;
A = 16'h00B9; B = 16'h00DC; #100;
A = 16'h00B9; B = 16'h00DD; #100;
A = 16'h00B9; B = 16'h00DE; #100;
A = 16'h00B9; B = 16'h00DF; #100;
A = 16'h00B9; B = 16'h00E0; #100;
A = 16'h00B9; B = 16'h00E1; #100;
A = 16'h00B9; B = 16'h00E2; #100;
A = 16'h00B9; B = 16'h00E3; #100;
A = 16'h00B9; B = 16'h00E4; #100;
A = 16'h00B9; B = 16'h00E5; #100;
A = 16'h00B9; B = 16'h00E6; #100;
A = 16'h00B9; B = 16'h00E7; #100;
A = 16'h00B9; B = 16'h00E8; #100;
A = 16'h00B9; B = 16'h00E9; #100;
A = 16'h00B9; B = 16'h00EA; #100;
A = 16'h00B9; B = 16'h00EB; #100;
A = 16'h00B9; B = 16'h00EC; #100;
A = 16'h00B9; B = 16'h00ED; #100;
A = 16'h00B9; B = 16'h00EE; #100;
A = 16'h00B9; B = 16'h00EF; #100;
A = 16'h00B9; B = 16'h00F0; #100;
A = 16'h00B9; B = 16'h00F1; #100;
A = 16'h00B9; B = 16'h00F2; #100;
A = 16'h00B9; B = 16'h00F3; #100;
A = 16'h00B9; B = 16'h00F4; #100;
A = 16'h00B9; B = 16'h00F5; #100;
A = 16'h00B9; B = 16'h00F6; #100;
A = 16'h00B9; B = 16'h00F7; #100;
A = 16'h00B9; B = 16'h00F8; #100;
A = 16'h00B9; B = 16'h00F9; #100;
A = 16'h00B9; B = 16'h00FA; #100;
A = 16'h00B9; B = 16'h00FB; #100;
A = 16'h00B9; B = 16'h00FC; #100;
A = 16'h00B9; B = 16'h00FD; #100;
A = 16'h00B9; B = 16'h00FE; #100;
A = 16'h00B9; B = 16'h00FF; #100;
A = 16'h00BA; B = 16'h000; #100;
A = 16'h00BA; B = 16'h001; #100;
A = 16'h00BA; B = 16'h002; #100;
A = 16'h00BA; B = 16'h003; #100;
A = 16'h00BA; B = 16'h004; #100;
A = 16'h00BA; B = 16'h005; #100;
A = 16'h00BA; B = 16'h006; #100;
A = 16'h00BA; B = 16'h007; #100;
A = 16'h00BA; B = 16'h008; #100;
A = 16'h00BA; B = 16'h009; #100;
A = 16'h00BA; B = 16'h00A; #100;
A = 16'h00BA; B = 16'h00B; #100;
A = 16'h00BA; B = 16'h00C; #100;
A = 16'h00BA; B = 16'h00D; #100;
A = 16'h00BA; B = 16'h00E; #100;
A = 16'h00BA; B = 16'h00F; #100;
A = 16'h00BA; B = 16'h0010; #100;
A = 16'h00BA; B = 16'h0011; #100;
A = 16'h00BA; B = 16'h0012; #100;
A = 16'h00BA; B = 16'h0013; #100;
A = 16'h00BA; B = 16'h0014; #100;
A = 16'h00BA; B = 16'h0015; #100;
A = 16'h00BA; B = 16'h0016; #100;
A = 16'h00BA; B = 16'h0017; #100;
A = 16'h00BA; B = 16'h0018; #100;
A = 16'h00BA; B = 16'h0019; #100;
A = 16'h00BA; B = 16'h001A; #100;
A = 16'h00BA; B = 16'h001B; #100;
A = 16'h00BA; B = 16'h001C; #100;
A = 16'h00BA; B = 16'h001D; #100;
A = 16'h00BA; B = 16'h001E; #100;
A = 16'h00BA; B = 16'h001F; #100;
A = 16'h00BA; B = 16'h0020; #100;
A = 16'h00BA; B = 16'h0021; #100;
A = 16'h00BA; B = 16'h0022; #100;
A = 16'h00BA; B = 16'h0023; #100;
A = 16'h00BA; B = 16'h0024; #100;
A = 16'h00BA; B = 16'h0025; #100;
A = 16'h00BA; B = 16'h0026; #100;
A = 16'h00BA; B = 16'h0027; #100;
A = 16'h00BA; B = 16'h0028; #100;
A = 16'h00BA; B = 16'h0029; #100;
A = 16'h00BA; B = 16'h002A; #100;
A = 16'h00BA; B = 16'h002B; #100;
A = 16'h00BA; B = 16'h002C; #100;
A = 16'h00BA; B = 16'h002D; #100;
A = 16'h00BA; B = 16'h002E; #100;
A = 16'h00BA; B = 16'h002F; #100;
A = 16'h00BA; B = 16'h0030; #100;
A = 16'h00BA; B = 16'h0031; #100;
A = 16'h00BA; B = 16'h0032; #100;
A = 16'h00BA; B = 16'h0033; #100;
A = 16'h00BA; B = 16'h0034; #100;
A = 16'h00BA; B = 16'h0035; #100;
A = 16'h00BA; B = 16'h0036; #100;
A = 16'h00BA; B = 16'h0037; #100;
A = 16'h00BA; B = 16'h0038; #100;
A = 16'h00BA; B = 16'h0039; #100;
A = 16'h00BA; B = 16'h003A; #100;
A = 16'h00BA; B = 16'h003B; #100;
A = 16'h00BA; B = 16'h003C; #100;
A = 16'h00BA; B = 16'h003D; #100;
A = 16'h00BA; B = 16'h003E; #100;
A = 16'h00BA; B = 16'h003F; #100;
A = 16'h00BA; B = 16'h0040; #100;
A = 16'h00BA; B = 16'h0041; #100;
A = 16'h00BA; B = 16'h0042; #100;
A = 16'h00BA; B = 16'h0043; #100;
A = 16'h00BA; B = 16'h0044; #100;
A = 16'h00BA; B = 16'h0045; #100;
A = 16'h00BA; B = 16'h0046; #100;
A = 16'h00BA; B = 16'h0047; #100;
A = 16'h00BA; B = 16'h0048; #100;
A = 16'h00BA; B = 16'h0049; #100;
A = 16'h00BA; B = 16'h004A; #100;
A = 16'h00BA; B = 16'h004B; #100;
A = 16'h00BA; B = 16'h004C; #100;
A = 16'h00BA; B = 16'h004D; #100;
A = 16'h00BA; B = 16'h004E; #100;
A = 16'h00BA; B = 16'h004F; #100;
A = 16'h00BA; B = 16'h0050; #100;
A = 16'h00BA; B = 16'h0051; #100;
A = 16'h00BA; B = 16'h0052; #100;
A = 16'h00BA; B = 16'h0053; #100;
A = 16'h00BA; B = 16'h0054; #100;
A = 16'h00BA; B = 16'h0055; #100;
A = 16'h00BA; B = 16'h0056; #100;
A = 16'h00BA; B = 16'h0057; #100;
A = 16'h00BA; B = 16'h0058; #100;
A = 16'h00BA; B = 16'h0059; #100;
A = 16'h00BA; B = 16'h005A; #100;
A = 16'h00BA; B = 16'h005B; #100;
A = 16'h00BA; B = 16'h005C; #100;
A = 16'h00BA; B = 16'h005D; #100;
A = 16'h00BA; B = 16'h005E; #100;
A = 16'h00BA; B = 16'h005F; #100;
A = 16'h00BA; B = 16'h0060; #100;
A = 16'h00BA; B = 16'h0061; #100;
A = 16'h00BA; B = 16'h0062; #100;
A = 16'h00BA; B = 16'h0063; #100;
A = 16'h00BA; B = 16'h0064; #100;
A = 16'h00BA; B = 16'h0065; #100;
A = 16'h00BA; B = 16'h0066; #100;
A = 16'h00BA; B = 16'h0067; #100;
A = 16'h00BA; B = 16'h0068; #100;
A = 16'h00BA; B = 16'h0069; #100;
A = 16'h00BA; B = 16'h006A; #100;
A = 16'h00BA; B = 16'h006B; #100;
A = 16'h00BA; B = 16'h006C; #100;
A = 16'h00BA; B = 16'h006D; #100;
A = 16'h00BA; B = 16'h006E; #100;
A = 16'h00BA; B = 16'h006F; #100;
A = 16'h00BA; B = 16'h0070; #100;
A = 16'h00BA; B = 16'h0071; #100;
A = 16'h00BA; B = 16'h0072; #100;
A = 16'h00BA; B = 16'h0073; #100;
A = 16'h00BA; B = 16'h0074; #100;
A = 16'h00BA; B = 16'h0075; #100;
A = 16'h00BA; B = 16'h0076; #100;
A = 16'h00BA; B = 16'h0077; #100;
A = 16'h00BA; B = 16'h0078; #100;
A = 16'h00BA; B = 16'h0079; #100;
A = 16'h00BA; B = 16'h007A; #100;
A = 16'h00BA; B = 16'h007B; #100;
A = 16'h00BA; B = 16'h007C; #100;
A = 16'h00BA; B = 16'h007D; #100;
A = 16'h00BA; B = 16'h007E; #100;
A = 16'h00BA; B = 16'h007F; #100;
A = 16'h00BA; B = 16'h0080; #100;
A = 16'h00BA; B = 16'h0081; #100;
A = 16'h00BA; B = 16'h0082; #100;
A = 16'h00BA; B = 16'h0083; #100;
A = 16'h00BA; B = 16'h0084; #100;
A = 16'h00BA; B = 16'h0085; #100;
A = 16'h00BA; B = 16'h0086; #100;
A = 16'h00BA; B = 16'h0087; #100;
A = 16'h00BA; B = 16'h0088; #100;
A = 16'h00BA; B = 16'h0089; #100;
A = 16'h00BA; B = 16'h008A; #100;
A = 16'h00BA; B = 16'h008B; #100;
A = 16'h00BA; B = 16'h008C; #100;
A = 16'h00BA; B = 16'h008D; #100;
A = 16'h00BA; B = 16'h008E; #100;
A = 16'h00BA; B = 16'h008F; #100;
A = 16'h00BA; B = 16'h0090; #100;
A = 16'h00BA; B = 16'h0091; #100;
A = 16'h00BA; B = 16'h0092; #100;
A = 16'h00BA; B = 16'h0093; #100;
A = 16'h00BA; B = 16'h0094; #100;
A = 16'h00BA; B = 16'h0095; #100;
A = 16'h00BA; B = 16'h0096; #100;
A = 16'h00BA; B = 16'h0097; #100;
A = 16'h00BA; B = 16'h0098; #100;
A = 16'h00BA; B = 16'h0099; #100;
A = 16'h00BA; B = 16'h009A; #100;
A = 16'h00BA; B = 16'h009B; #100;
A = 16'h00BA; B = 16'h009C; #100;
A = 16'h00BA; B = 16'h009D; #100;
A = 16'h00BA; B = 16'h009E; #100;
A = 16'h00BA; B = 16'h009F; #100;
A = 16'h00BA; B = 16'h00A0; #100;
A = 16'h00BA; B = 16'h00A1; #100;
A = 16'h00BA; B = 16'h00A2; #100;
A = 16'h00BA; B = 16'h00A3; #100;
A = 16'h00BA; B = 16'h00A4; #100;
A = 16'h00BA; B = 16'h00A5; #100;
A = 16'h00BA; B = 16'h00A6; #100;
A = 16'h00BA; B = 16'h00A7; #100;
A = 16'h00BA; B = 16'h00A8; #100;
A = 16'h00BA; B = 16'h00A9; #100;
A = 16'h00BA; B = 16'h00AA; #100;
A = 16'h00BA; B = 16'h00AB; #100;
A = 16'h00BA; B = 16'h00AC; #100;
A = 16'h00BA; B = 16'h00AD; #100;
A = 16'h00BA; B = 16'h00AE; #100;
A = 16'h00BA; B = 16'h00AF; #100;
A = 16'h00BA; B = 16'h00B0; #100;
A = 16'h00BA; B = 16'h00B1; #100;
A = 16'h00BA; B = 16'h00B2; #100;
A = 16'h00BA; B = 16'h00B3; #100;
A = 16'h00BA; B = 16'h00B4; #100;
A = 16'h00BA; B = 16'h00B5; #100;
A = 16'h00BA; B = 16'h00B6; #100;
A = 16'h00BA; B = 16'h00B7; #100;
A = 16'h00BA; B = 16'h00B8; #100;
A = 16'h00BA; B = 16'h00B9; #100;
A = 16'h00BA; B = 16'h00BA; #100;
A = 16'h00BA; B = 16'h00BB; #100;
A = 16'h00BA; B = 16'h00BC; #100;
A = 16'h00BA; B = 16'h00BD; #100;
A = 16'h00BA; B = 16'h00BE; #100;
A = 16'h00BA; B = 16'h00BF; #100;
A = 16'h00BA; B = 16'h00C0; #100;
A = 16'h00BA; B = 16'h00C1; #100;
A = 16'h00BA; B = 16'h00C2; #100;
A = 16'h00BA; B = 16'h00C3; #100;
A = 16'h00BA; B = 16'h00C4; #100;
A = 16'h00BA; B = 16'h00C5; #100;
A = 16'h00BA; B = 16'h00C6; #100;
A = 16'h00BA; B = 16'h00C7; #100;
A = 16'h00BA; B = 16'h00C8; #100;
A = 16'h00BA; B = 16'h00C9; #100;
A = 16'h00BA; B = 16'h00CA; #100;
A = 16'h00BA; B = 16'h00CB; #100;
A = 16'h00BA; B = 16'h00CC; #100;
A = 16'h00BA; B = 16'h00CD; #100;
A = 16'h00BA; B = 16'h00CE; #100;
A = 16'h00BA; B = 16'h00CF; #100;
A = 16'h00BA; B = 16'h00D0; #100;
A = 16'h00BA; B = 16'h00D1; #100;
A = 16'h00BA; B = 16'h00D2; #100;
A = 16'h00BA; B = 16'h00D3; #100;
A = 16'h00BA; B = 16'h00D4; #100;
A = 16'h00BA; B = 16'h00D5; #100;
A = 16'h00BA; B = 16'h00D6; #100;
A = 16'h00BA; B = 16'h00D7; #100;
A = 16'h00BA; B = 16'h00D8; #100;
A = 16'h00BA; B = 16'h00D9; #100;
A = 16'h00BA; B = 16'h00DA; #100;
A = 16'h00BA; B = 16'h00DB; #100;
A = 16'h00BA; B = 16'h00DC; #100;
A = 16'h00BA; B = 16'h00DD; #100;
A = 16'h00BA; B = 16'h00DE; #100;
A = 16'h00BA; B = 16'h00DF; #100;
A = 16'h00BA; B = 16'h00E0; #100;
A = 16'h00BA; B = 16'h00E1; #100;
A = 16'h00BA; B = 16'h00E2; #100;
A = 16'h00BA; B = 16'h00E3; #100;
A = 16'h00BA; B = 16'h00E4; #100;
A = 16'h00BA; B = 16'h00E5; #100;
A = 16'h00BA; B = 16'h00E6; #100;
A = 16'h00BA; B = 16'h00E7; #100;
A = 16'h00BA; B = 16'h00E8; #100;
A = 16'h00BA; B = 16'h00E9; #100;
A = 16'h00BA; B = 16'h00EA; #100;
A = 16'h00BA; B = 16'h00EB; #100;
A = 16'h00BA; B = 16'h00EC; #100;
A = 16'h00BA; B = 16'h00ED; #100;
A = 16'h00BA; B = 16'h00EE; #100;
A = 16'h00BA; B = 16'h00EF; #100;
A = 16'h00BA; B = 16'h00F0; #100;
A = 16'h00BA; B = 16'h00F1; #100;
A = 16'h00BA; B = 16'h00F2; #100;
A = 16'h00BA; B = 16'h00F3; #100;
A = 16'h00BA; B = 16'h00F4; #100;
A = 16'h00BA; B = 16'h00F5; #100;
A = 16'h00BA; B = 16'h00F6; #100;
A = 16'h00BA; B = 16'h00F7; #100;
A = 16'h00BA; B = 16'h00F8; #100;
A = 16'h00BA; B = 16'h00F9; #100;
A = 16'h00BA; B = 16'h00FA; #100;
A = 16'h00BA; B = 16'h00FB; #100;
A = 16'h00BA; B = 16'h00FC; #100;
A = 16'h00BA; B = 16'h00FD; #100;
A = 16'h00BA; B = 16'h00FE; #100;
A = 16'h00BA; B = 16'h00FF; #100;
A = 16'h00BB; B = 16'h000; #100;
A = 16'h00BB; B = 16'h001; #100;
A = 16'h00BB; B = 16'h002; #100;
A = 16'h00BB; B = 16'h003; #100;
A = 16'h00BB; B = 16'h004; #100;
A = 16'h00BB; B = 16'h005; #100;
A = 16'h00BB; B = 16'h006; #100;
A = 16'h00BB; B = 16'h007; #100;
A = 16'h00BB; B = 16'h008; #100;
A = 16'h00BB; B = 16'h009; #100;
A = 16'h00BB; B = 16'h00A; #100;
A = 16'h00BB; B = 16'h00B; #100;
A = 16'h00BB; B = 16'h00C; #100;
A = 16'h00BB; B = 16'h00D; #100;
A = 16'h00BB; B = 16'h00E; #100;
A = 16'h00BB; B = 16'h00F; #100;
A = 16'h00BB; B = 16'h0010; #100;
A = 16'h00BB; B = 16'h0011; #100;
A = 16'h00BB; B = 16'h0012; #100;
A = 16'h00BB; B = 16'h0013; #100;
A = 16'h00BB; B = 16'h0014; #100;
A = 16'h00BB; B = 16'h0015; #100;
A = 16'h00BB; B = 16'h0016; #100;
A = 16'h00BB; B = 16'h0017; #100;
A = 16'h00BB; B = 16'h0018; #100;
A = 16'h00BB; B = 16'h0019; #100;
A = 16'h00BB; B = 16'h001A; #100;
A = 16'h00BB; B = 16'h001B; #100;
A = 16'h00BB; B = 16'h001C; #100;
A = 16'h00BB; B = 16'h001D; #100;
A = 16'h00BB; B = 16'h001E; #100;
A = 16'h00BB; B = 16'h001F; #100;
A = 16'h00BB; B = 16'h0020; #100;
A = 16'h00BB; B = 16'h0021; #100;
A = 16'h00BB; B = 16'h0022; #100;
A = 16'h00BB; B = 16'h0023; #100;
A = 16'h00BB; B = 16'h0024; #100;
A = 16'h00BB; B = 16'h0025; #100;
A = 16'h00BB; B = 16'h0026; #100;
A = 16'h00BB; B = 16'h0027; #100;
A = 16'h00BB; B = 16'h0028; #100;
A = 16'h00BB; B = 16'h0029; #100;
A = 16'h00BB; B = 16'h002A; #100;
A = 16'h00BB; B = 16'h002B; #100;
A = 16'h00BB; B = 16'h002C; #100;
A = 16'h00BB; B = 16'h002D; #100;
A = 16'h00BB; B = 16'h002E; #100;
A = 16'h00BB; B = 16'h002F; #100;
A = 16'h00BB; B = 16'h0030; #100;
A = 16'h00BB; B = 16'h0031; #100;
A = 16'h00BB; B = 16'h0032; #100;
A = 16'h00BB; B = 16'h0033; #100;
A = 16'h00BB; B = 16'h0034; #100;
A = 16'h00BB; B = 16'h0035; #100;
A = 16'h00BB; B = 16'h0036; #100;
A = 16'h00BB; B = 16'h0037; #100;
A = 16'h00BB; B = 16'h0038; #100;
A = 16'h00BB; B = 16'h0039; #100;
A = 16'h00BB; B = 16'h003A; #100;
A = 16'h00BB; B = 16'h003B; #100;
A = 16'h00BB; B = 16'h003C; #100;
A = 16'h00BB; B = 16'h003D; #100;
A = 16'h00BB; B = 16'h003E; #100;
A = 16'h00BB; B = 16'h003F; #100;
A = 16'h00BB; B = 16'h0040; #100;
A = 16'h00BB; B = 16'h0041; #100;
A = 16'h00BB; B = 16'h0042; #100;
A = 16'h00BB; B = 16'h0043; #100;
A = 16'h00BB; B = 16'h0044; #100;
A = 16'h00BB; B = 16'h0045; #100;
A = 16'h00BB; B = 16'h0046; #100;
A = 16'h00BB; B = 16'h0047; #100;
A = 16'h00BB; B = 16'h0048; #100;
A = 16'h00BB; B = 16'h0049; #100;
A = 16'h00BB; B = 16'h004A; #100;
A = 16'h00BB; B = 16'h004B; #100;
A = 16'h00BB; B = 16'h004C; #100;
A = 16'h00BB; B = 16'h004D; #100;
A = 16'h00BB; B = 16'h004E; #100;
A = 16'h00BB; B = 16'h004F; #100;
A = 16'h00BB; B = 16'h0050; #100;
A = 16'h00BB; B = 16'h0051; #100;
A = 16'h00BB; B = 16'h0052; #100;
A = 16'h00BB; B = 16'h0053; #100;
A = 16'h00BB; B = 16'h0054; #100;
A = 16'h00BB; B = 16'h0055; #100;
A = 16'h00BB; B = 16'h0056; #100;
A = 16'h00BB; B = 16'h0057; #100;
A = 16'h00BB; B = 16'h0058; #100;
A = 16'h00BB; B = 16'h0059; #100;
A = 16'h00BB; B = 16'h005A; #100;
A = 16'h00BB; B = 16'h005B; #100;
A = 16'h00BB; B = 16'h005C; #100;
A = 16'h00BB; B = 16'h005D; #100;
A = 16'h00BB; B = 16'h005E; #100;
A = 16'h00BB; B = 16'h005F; #100;
A = 16'h00BB; B = 16'h0060; #100;
A = 16'h00BB; B = 16'h0061; #100;
A = 16'h00BB; B = 16'h0062; #100;
A = 16'h00BB; B = 16'h0063; #100;
A = 16'h00BB; B = 16'h0064; #100;
A = 16'h00BB; B = 16'h0065; #100;
A = 16'h00BB; B = 16'h0066; #100;
A = 16'h00BB; B = 16'h0067; #100;
A = 16'h00BB; B = 16'h0068; #100;
A = 16'h00BB; B = 16'h0069; #100;
A = 16'h00BB; B = 16'h006A; #100;
A = 16'h00BB; B = 16'h006B; #100;
A = 16'h00BB; B = 16'h006C; #100;
A = 16'h00BB; B = 16'h006D; #100;
A = 16'h00BB; B = 16'h006E; #100;
A = 16'h00BB; B = 16'h006F; #100;
A = 16'h00BB; B = 16'h0070; #100;
A = 16'h00BB; B = 16'h0071; #100;
A = 16'h00BB; B = 16'h0072; #100;
A = 16'h00BB; B = 16'h0073; #100;
A = 16'h00BB; B = 16'h0074; #100;
A = 16'h00BB; B = 16'h0075; #100;
A = 16'h00BB; B = 16'h0076; #100;
A = 16'h00BB; B = 16'h0077; #100;
A = 16'h00BB; B = 16'h0078; #100;
A = 16'h00BB; B = 16'h0079; #100;
A = 16'h00BB; B = 16'h007A; #100;
A = 16'h00BB; B = 16'h007B; #100;
A = 16'h00BB; B = 16'h007C; #100;
A = 16'h00BB; B = 16'h007D; #100;
A = 16'h00BB; B = 16'h007E; #100;
A = 16'h00BB; B = 16'h007F; #100;
A = 16'h00BB; B = 16'h0080; #100;
A = 16'h00BB; B = 16'h0081; #100;
A = 16'h00BB; B = 16'h0082; #100;
A = 16'h00BB; B = 16'h0083; #100;
A = 16'h00BB; B = 16'h0084; #100;
A = 16'h00BB; B = 16'h0085; #100;
A = 16'h00BB; B = 16'h0086; #100;
A = 16'h00BB; B = 16'h0087; #100;
A = 16'h00BB; B = 16'h0088; #100;
A = 16'h00BB; B = 16'h0089; #100;
A = 16'h00BB; B = 16'h008A; #100;
A = 16'h00BB; B = 16'h008B; #100;
A = 16'h00BB; B = 16'h008C; #100;
A = 16'h00BB; B = 16'h008D; #100;
A = 16'h00BB; B = 16'h008E; #100;
A = 16'h00BB; B = 16'h008F; #100;
A = 16'h00BB; B = 16'h0090; #100;
A = 16'h00BB; B = 16'h0091; #100;
A = 16'h00BB; B = 16'h0092; #100;
A = 16'h00BB; B = 16'h0093; #100;
A = 16'h00BB; B = 16'h0094; #100;
A = 16'h00BB; B = 16'h0095; #100;
A = 16'h00BB; B = 16'h0096; #100;
A = 16'h00BB; B = 16'h0097; #100;
A = 16'h00BB; B = 16'h0098; #100;
A = 16'h00BB; B = 16'h0099; #100;
A = 16'h00BB; B = 16'h009A; #100;
A = 16'h00BB; B = 16'h009B; #100;
A = 16'h00BB; B = 16'h009C; #100;
A = 16'h00BB; B = 16'h009D; #100;
A = 16'h00BB; B = 16'h009E; #100;
A = 16'h00BB; B = 16'h009F; #100;
A = 16'h00BB; B = 16'h00A0; #100;
A = 16'h00BB; B = 16'h00A1; #100;
A = 16'h00BB; B = 16'h00A2; #100;
A = 16'h00BB; B = 16'h00A3; #100;
A = 16'h00BB; B = 16'h00A4; #100;
A = 16'h00BB; B = 16'h00A5; #100;
A = 16'h00BB; B = 16'h00A6; #100;
A = 16'h00BB; B = 16'h00A7; #100;
A = 16'h00BB; B = 16'h00A8; #100;
A = 16'h00BB; B = 16'h00A9; #100;
A = 16'h00BB; B = 16'h00AA; #100;
A = 16'h00BB; B = 16'h00AB; #100;
A = 16'h00BB; B = 16'h00AC; #100;
A = 16'h00BB; B = 16'h00AD; #100;
A = 16'h00BB; B = 16'h00AE; #100;
A = 16'h00BB; B = 16'h00AF; #100;
A = 16'h00BB; B = 16'h00B0; #100;
A = 16'h00BB; B = 16'h00B1; #100;
A = 16'h00BB; B = 16'h00B2; #100;
A = 16'h00BB; B = 16'h00B3; #100;
A = 16'h00BB; B = 16'h00B4; #100;
A = 16'h00BB; B = 16'h00B5; #100;
A = 16'h00BB; B = 16'h00B6; #100;
A = 16'h00BB; B = 16'h00B7; #100;
A = 16'h00BB; B = 16'h00B8; #100;
A = 16'h00BB; B = 16'h00B9; #100;
A = 16'h00BB; B = 16'h00BA; #100;
A = 16'h00BB; B = 16'h00BB; #100;
A = 16'h00BB; B = 16'h00BC; #100;
A = 16'h00BB; B = 16'h00BD; #100;
A = 16'h00BB; B = 16'h00BE; #100;
A = 16'h00BB; B = 16'h00BF; #100;
A = 16'h00BB; B = 16'h00C0; #100;
A = 16'h00BB; B = 16'h00C1; #100;
A = 16'h00BB; B = 16'h00C2; #100;
A = 16'h00BB; B = 16'h00C3; #100;
A = 16'h00BB; B = 16'h00C4; #100;
A = 16'h00BB; B = 16'h00C5; #100;
A = 16'h00BB; B = 16'h00C6; #100;
A = 16'h00BB; B = 16'h00C7; #100;
A = 16'h00BB; B = 16'h00C8; #100;
A = 16'h00BB; B = 16'h00C9; #100;
A = 16'h00BB; B = 16'h00CA; #100;
A = 16'h00BB; B = 16'h00CB; #100;
A = 16'h00BB; B = 16'h00CC; #100;
A = 16'h00BB; B = 16'h00CD; #100;
A = 16'h00BB; B = 16'h00CE; #100;
A = 16'h00BB; B = 16'h00CF; #100;
A = 16'h00BB; B = 16'h00D0; #100;
A = 16'h00BB; B = 16'h00D1; #100;
A = 16'h00BB; B = 16'h00D2; #100;
A = 16'h00BB; B = 16'h00D3; #100;
A = 16'h00BB; B = 16'h00D4; #100;
A = 16'h00BB; B = 16'h00D5; #100;
A = 16'h00BB; B = 16'h00D6; #100;
A = 16'h00BB; B = 16'h00D7; #100;
A = 16'h00BB; B = 16'h00D8; #100;
A = 16'h00BB; B = 16'h00D9; #100;
A = 16'h00BB; B = 16'h00DA; #100;
A = 16'h00BB; B = 16'h00DB; #100;
A = 16'h00BB; B = 16'h00DC; #100;
A = 16'h00BB; B = 16'h00DD; #100;
A = 16'h00BB; B = 16'h00DE; #100;
A = 16'h00BB; B = 16'h00DF; #100;
A = 16'h00BB; B = 16'h00E0; #100;
A = 16'h00BB; B = 16'h00E1; #100;
A = 16'h00BB; B = 16'h00E2; #100;
A = 16'h00BB; B = 16'h00E3; #100;
A = 16'h00BB; B = 16'h00E4; #100;
A = 16'h00BB; B = 16'h00E5; #100;
A = 16'h00BB; B = 16'h00E6; #100;
A = 16'h00BB; B = 16'h00E7; #100;
A = 16'h00BB; B = 16'h00E8; #100;
A = 16'h00BB; B = 16'h00E9; #100;
A = 16'h00BB; B = 16'h00EA; #100;
A = 16'h00BB; B = 16'h00EB; #100;
A = 16'h00BB; B = 16'h00EC; #100;
A = 16'h00BB; B = 16'h00ED; #100;
A = 16'h00BB; B = 16'h00EE; #100;
A = 16'h00BB; B = 16'h00EF; #100;
A = 16'h00BB; B = 16'h00F0; #100;
A = 16'h00BB; B = 16'h00F1; #100;
A = 16'h00BB; B = 16'h00F2; #100;
A = 16'h00BB; B = 16'h00F3; #100;
A = 16'h00BB; B = 16'h00F4; #100;
A = 16'h00BB; B = 16'h00F5; #100;
A = 16'h00BB; B = 16'h00F6; #100;
A = 16'h00BB; B = 16'h00F7; #100;
A = 16'h00BB; B = 16'h00F8; #100;
A = 16'h00BB; B = 16'h00F9; #100;
A = 16'h00BB; B = 16'h00FA; #100;
A = 16'h00BB; B = 16'h00FB; #100;
A = 16'h00BB; B = 16'h00FC; #100;
A = 16'h00BB; B = 16'h00FD; #100;
A = 16'h00BB; B = 16'h00FE; #100;
A = 16'h00BB; B = 16'h00FF; #100;
A = 16'h00BC; B = 16'h000; #100;
A = 16'h00BC; B = 16'h001; #100;
A = 16'h00BC; B = 16'h002; #100;
A = 16'h00BC; B = 16'h003; #100;
A = 16'h00BC; B = 16'h004; #100;
A = 16'h00BC; B = 16'h005; #100;
A = 16'h00BC; B = 16'h006; #100;
A = 16'h00BC; B = 16'h007; #100;
A = 16'h00BC; B = 16'h008; #100;
A = 16'h00BC; B = 16'h009; #100;
A = 16'h00BC; B = 16'h00A; #100;
A = 16'h00BC; B = 16'h00B; #100;
A = 16'h00BC; B = 16'h00C; #100;
A = 16'h00BC; B = 16'h00D; #100;
A = 16'h00BC; B = 16'h00E; #100;
A = 16'h00BC; B = 16'h00F; #100;
A = 16'h00BC; B = 16'h0010; #100;
A = 16'h00BC; B = 16'h0011; #100;
A = 16'h00BC; B = 16'h0012; #100;
A = 16'h00BC; B = 16'h0013; #100;
A = 16'h00BC; B = 16'h0014; #100;
A = 16'h00BC; B = 16'h0015; #100;
A = 16'h00BC; B = 16'h0016; #100;
A = 16'h00BC; B = 16'h0017; #100;
A = 16'h00BC; B = 16'h0018; #100;
A = 16'h00BC; B = 16'h0019; #100;
A = 16'h00BC; B = 16'h001A; #100;
A = 16'h00BC; B = 16'h001B; #100;
A = 16'h00BC; B = 16'h001C; #100;
A = 16'h00BC; B = 16'h001D; #100;
A = 16'h00BC; B = 16'h001E; #100;
A = 16'h00BC; B = 16'h001F; #100;
A = 16'h00BC; B = 16'h0020; #100;
A = 16'h00BC; B = 16'h0021; #100;
A = 16'h00BC; B = 16'h0022; #100;
A = 16'h00BC; B = 16'h0023; #100;
A = 16'h00BC; B = 16'h0024; #100;
A = 16'h00BC; B = 16'h0025; #100;
A = 16'h00BC; B = 16'h0026; #100;
A = 16'h00BC; B = 16'h0027; #100;
A = 16'h00BC; B = 16'h0028; #100;
A = 16'h00BC; B = 16'h0029; #100;
A = 16'h00BC; B = 16'h002A; #100;
A = 16'h00BC; B = 16'h002B; #100;
A = 16'h00BC; B = 16'h002C; #100;
A = 16'h00BC; B = 16'h002D; #100;
A = 16'h00BC; B = 16'h002E; #100;
A = 16'h00BC; B = 16'h002F; #100;
A = 16'h00BC; B = 16'h0030; #100;
A = 16'h00BC; B = 16'h0031; #100;
A = 16'h00BC; B = 16'h0032; #100;
A = 16'h00BC; B = 16'h0033; #100;
A = 16'h00BC; B = 16'h0034; #100;
A = 16'h00BC; B = 16'h0035; #100;
A = 16'h00BC; B = 16'h0036; #100;
A = 16'h00BC; B = 16'h0037; #100;
A = 16'h00BC; B = 16'h0038; #100;
A = 16'h00BC; B = 16'h0039; #100;
A = 16'h00BC; B = 16'h003A; #100;
A = 16'h00BC; B = 16'h003B; #100;
A = 16'h00BC; B = 16'h003C; #100;
A = 16'h00BC; B = 16'h003D; #100;
A = 16'h00BC; B = 16'h003E; #100;
A = 16'h00BC; B = 16'h003F; #100;
A = 16'h00BC; B = 16'h0040; #100;
A = 16'h00BC; B = 16'h0041; #100;
A = 16'h00BC; B = 16'h0042; #100;
A = 16'h00BC; B = 16'h0043; #100;
A = 16'h00BC; B = 16'h0044; #100;
A = 16'h00BC; B = 16'h0045; #100;
A = 16'h00BC; B = 16'h0046; #100;
A = 16'h00BC; B = 16'h0047; #100;
A = 16'h00BC; B = 16'h0048; #100;
A = 16'h00BC; B = 16'h0049; #100;
A = 16'h00BC; B = 16'h004A; #100;
A = 16'h00BC; B = 16'h004B; #100;
A = 16'h00BC; B = 16'h004C; #100;
A = 16'h00BC; B = 16'h004D; #100;
A = 16'h00BC; B = 16'h004E; #100;
A = 16'h00BC; B = 16'h004F; #100;
A = 16'h00BC; B = 16'h0050; #100;
A = 16'h00BC; B = 16'h0051; #100;
A = 16'h00BC; B = 16'h0052; #100;
A = 16'h00BC; B = 16'h0053; #100;
A = 16'h00BC; B = 16'h0054; #100;
A = 16'h00BC; B = 16'h0055; #100;
A = 16'h00BC; B = 16'h0056; #100;
A = 16'h00BC; B = 16'h0057; #100;
A = 16'h00BC; B = 16'h0058; #100;
A = 16'h00BC; B = 16'h0059; #100;
A = 16'h00BC; B = 16'h005A; #100;
A = 16'h00BC; B = 16'h005B; #100;
A = 16'h00BC; B = 16'h005C; #100;
A = 16'h00BC; B = 16'h005D; #100;
A = 16'h00BC; B = 16'h005E; #100;
A = 16'h00BC; B = 16'h005F; #100;
A = 16'h00BC; B = 16'h0060; #100;
A = 16'h00BC; B = 16'h0061; #100;
A = 16'h00BC; B = 16'h0062; #100;
A = 16'h00BC; B = 16'h0063; #100;
A = 16'h00BC; B = 16'h0064; #100;
A = 16'h00BC; B = 16'h0065; #100;
A = 16'h00BC; B = 16'h0066; #100;
A = 16'h00BC; B = 16'h0067; #100;
A = 16'h00BC; B = 16'h0068; #100;
A = 16'h00BC; B = 16'h0069; #100;
A = 16'h00BC; B = 16'h006A; #100;
A = 16'h00BC; B = 16'h006B; #100;
A = 16'h00BC; B = 16'h006C; #100;
A = 16'h00BC; B = 16'h006D; #100;
A = 16'h00BC; B = 16'h006E; #100;
A = 16'h00BC; B = 16'h006F; #100;
A = 16'h00BC; B = 16'h0070; #100;
A = 16'h00BC; B = 16'h0071; #100;
A = 16'h00BC; B = 16'h0072; #100;
A = 16'h00BC; B = 16'h0073; #100;
A = 16'h00BC; B = 16'h0074; #100;
A = 16'h00BC; B = 16'h0075; #100;
A = 16'h00BC; B = 16'h0076; #100;
A = 16'h00BC; B = 16'h0077; #100;
A = 16'h00BC; B = 16'h0078; #100;
A = 16'h00BC; B = 16'h0079; #100;
A = 16'h00BC; B = 16'h007A; #100;
A = 16'h00BC; B = 16'h007B; #100;
A = 16'h00BC; B = 16'h007C; #100;
A = 16'h00BC; B = 16'h007D; #100;
A = 16'h00BC; B = 16'h007E; #100;
A = 16'h00BC; B = 16'h007F; #100;
A = 16'h00BC; B = 16'h0080; #100;
A = 16'h00BC; B = 16'h0081; #100;
A = 16'h00BC; B = 16'h0082; #100;
A = 16'h00BC; B = 16'h0083; #100;
A = 16'h00BC; B = 16'h0084; #100;
A = 16'h00BC; B = 16'h0085; #100;
A = 16'h00BC; B = 16'h0086; #100;
A = 16'h00BC; B = 16'h0087; #100;
A = 16'h00BC; B = 16'h0088; #100;
A = 16'h00BC; B = 16'h0089; #100;
A = 16'h00BC; B = 16'h008A; #100;
A = 16'h00BC; B = 16'h008B; #100;
A = 16'h00BC; B = 16'h008C; #100;
A = 16'h00BC; B = 16'h008D; #100;
A = 16'h00BC; B = 16'h008E; #100;
A = 16'h00BC; B = 16'h008F; #100;
A = 16'h00BC; B = 16'h0090; #100;
A = 16'h00BC; B = 16'h0091; #100;
A = 16'h00BC; B = 16'h0092; #100;
A = 16'h00BC; B = 16'h0093; #100;
A = 16'h00BC; B = 16'h0094; #100;
A = 16'h00BC; B = 16'h0095; #100;
A = 16'h00BC; B = 16'h0096; #100;
A = 16'h00BC; B = 16'h0097; #100;
A = 16'h00BC; B = 16'h0098; #100;
A = 16'h00BC; B = 16'h0099; #100;
A = 16'h00BC; B = 16'h009A; #100;
A = 16'h00BC; B = 16'h009B; #100;
A = 16'h00BC; B = 16'h009C; #100;
A = 16'h00BC; B = 16'h009D; #100;
A = 16'h00BC; B = 16'h009E; #100;
A = 16'h00BC; B = 16'h009F; #100;
A = 16'h00BC; B = 16'h00A0; #100;
A = 16'h00BC; B = 16'h00A1; #100;
A = 16'h00BC; B = 16'h00A2; #100;
A = 16'h00BC; B = 16'h00A3; #100;
A = 16'h00BC; B = 16'h00A4; #100;
A = 16'h00BC; B = 16'h00A5; #100;
A = 16'h00BC; B = 16'h00A6; #100;
A = 16'h00BC; B = 16'h00A7; #100;
A = 16'h00BC; B = 16'h00A8; #100;
A = 16'h00BC; B = 16'h00A9; #100;
A = 16'h00BC; B = 16'h00AA; #100;
A = 16'h00BC; B = 16'h00AB; #100;
A = 16'h00BC; B = 16'h00AC; #100;
A = 16'h00BC; B = 16'h00AD; #100;
A = 16'h00BC; B = 16'h00AE; #100;
A = 16'h00BC; B = 16'h00AF; #100;
A = 16'h00BC; B = 16'h00B0; #100;
A = 16'h00BC; B = 16'h00B1; #100;
A = 16'h00BC; B = 16'h00B2; #100;
A = 16'h00BC; B = 16'h00B3; #100;
A = 16'h00BC; B = 16'h00B4; #100;
A = 16'h00BC; B = 16'h00B5; #100;
A = 16'h00BC; B = 16'h00B6; #100;
A = 16'h00BC; B = 16'h00B7; #100;
A = 16'h00BC; B = 16'h00B8; #100;
A = 16'h00BC; B = 16'h00B9; #100;
A = 16'h00BC; B = 16'h00BA; #100;
A = 16'h00BC; B = 16'h00BB; #100;
A = 16'h00BC; B = 16'h00BC; #100;
A = 16'h00BC; B = 16'h00BD; #100;
A = 16'h00BC; B = 16'h00BE; #100;
A = 16'h00BC; B = 16'h00BF; #100;
A = 16'h00BC; B = 16'h00C0; #100;
A = 16'h00BC; B = 16'h00C1; #100;
A = 16'h00BC; B = 16'h00C2; #100;
A = 16'h00BC; B = 16'h00C3; #100;
A = 16'h00BC; B = 16'h00C4; #100;
A = 16'h00BC; B = 16'h00C5; #100;
A = 16'h00BC; B = 16'h00C6; #100;
A = 16'h00BC; B = 16'h00C7; #100;
A = 16'h00BC; B = 16'h00C8; #100;
A = 16'h00BC; B = 16'h00C9; #100;
A = 16'h00BC; B = 16'h00CA; #100;
A = 16'h00BC; B = 16'h00CB; #100;
A = 16'h00BC; B = 16'h00CC; #100;
A = 16'h00BC; B = 16'h00CD; #100;
A = 16'h00BC; B = 16'h00CE; #100;
A = 16'h00BC; B = 16'h00CF; #100;
A = 16'h00BC; B = 16'h00D0; #100;
A = 16'h00BC; B = 16'h00D1; #100;
A = 16'h00BC; B = 16'h00D2; #100;
A = 16'h00BC; B = 16'h00D3; #100;
A = 16'h00BC; B = 16'h00D4; #100;
A = 16'h00BC; B = 16'h00D5; #100;
A = 16'h00BC; B = 16'h00D6; #100;
A = 16'h00BC; B = 16'h00D7; #100;
A = 16'h00BC; B = 16'h00D8; #100;
A = 16'h00BC; B = 16'h00D9; #100;
A = 16'h00BC; B = 16'h00DA; #100;
A = 16'h00BC; B = 16'h00DB; #100;
A = 16'h00BC; B = 16'h00DC; #100;
A = 16'h00BC; B = 16'h00DD; #100;
A = 16'h00BC; B = 16'h00DE; #100;
A = 16'h00BC; B = 16'h00DF; #100;
A = 16'h00BC; B = 16'h00E0; #100;
A = 16'h00BC; B = 16'h00E1; #100;
A = 16'h00BC; B = 16'h00E2; #100;
A = 16'h00BC; B = 16'h00E3; #100;
A = 16'h00BC; B = 16'h00E4; #100;
A = 16'h00BC; B = 16'h00E5; #100;
A = 16'h00BC; B = 16'h00E6; #100;
A = 16'h00BC; B = 16'h00E7; #100;
A = 16'h00BC; B = 16'h00E8; #100;
A = 16'h00BC; B = 16'h00E9; #100;
A = 16'h00BC; B = 16'h00EA; #100;
A = 16'h00BC; B = 16'h00EB; #100;
A = 16'h00BC; B = 16'h00EC; #100;
A = 16'h00BC; B = 16'h00ED; #100;
A = 16'h00BC; B = 16'h00EE; #100;
A = 16'h00BC; B = 16'h00EF; #100;
A = 16'h00BC; B = 16'h00F0; #100;
A = 16'h00BC; B = 16'h00F1; #100;
A = 16'h00BC; B = 16'h00F2; #100;
A = 16'h00BC; B = 16'h00F3; #100;
A = 16'h00BC; B = 16'h00F4; #100;
A = 16'h00BC; B = 16'h00F5; #100;
A = 16'h00BC; B = 16'h00F6; #100;
A = 16'h00BC; B = 16'h00F7; #100;
A = 16'h00BC; B = 16'h00F8; #100;
A = 16'h00BC; B = 16'h00F9; #100;
A = 16'h00BC; B = 16'h00FA; #100;
A = 16'h00BC; B = 16'h00FB; #100;
A = 16'h00BC; B = 16'h00FC; #100;
A = 16'h00BC; B = 16'h00FD; #100;
A = 16'h00BC; B = 16'h00FE; #100;
A = 16'h00BC; B = 16'h00FF; #100;
A = 16'h00BD; B = 16'h000; #100;
A = 16'h00BD; B = 16'h001; #100;
A = 16'h00BD; B = 16'h002; #100;
A = 16'h00BD; B = 16'h003; #100;
A = 16'h00BD; B = 16'h004; #100;
A = 16'h00BD; B = 16'h005; #100;
A = 16'h00BD; B = 16'h006; #100;
A = 16'h00BD; B = 16'h007; #100;
A = 16'h00BD; B = 16'h008; #100;
A = 16'h00BD; B = 16'h009; #100;
A = 16'h00BD; B = 16'h00A; #100;
A = 16'h00BD; B = 16'h00B; #100;
A = 16'h00BD; B = 16'h00C; #100;
A = 16'h00BD; B = 16'h00D; #100;
A = 16'h00BD; B = 16'h00E; #100;
A = 16'h00BD; B = 16'h00F; #100;
A = 16'h00BD; B = 16'h0010; #100;
A = 16'h00BD; B = 16'h0011; #100;
A = 16'h00BD; B = 16'h0012; #100;
A = 16'h00BD; B = 16'h0013; #100;
A = 16'h00BD; B = 16'h0014; #100;
A = 16'h00BD; B = 16'h0015; #100;
A = 16'h00BD; B = 16'h0016; #100;
A = 16'h00BD; B = 16'h0017; #100;
A = 16'h00BD; B = 16'h0018; #100;
A = 16'h00BD; B = 16'h0019; #100;
A = 16'h00BD; B = 16'h001A; #100;
A = 16'h00BD; B = 16'h001B; #100;
A = 16'h00BD; B = 16'h001C; #100;
A = 16'h00BD; B = 16'h001D; #100;
A = 16'h00BD; B = 16'h001E; #100;
A = 16'h00BD; B = 16'h001F; #100;
A = 16'h00BD; B = 16'h0020; #100;
A = 16'h00BD; B = 16'h0021; #100;
A = 16'h00BD; B = 16'h0022; #100;
A = 16'h00BD; B = 16'h0023; #100;
A = 16'h00BD; B = 16'h0024; #100;
A = 16'h00BD; B = 16'h0025; #100;
A = 16'h00BD; B = 16'h0026; #100;
A = 16'h00BD; B = 16'h0027; #100;
A = 16'h00BD; B = 16'h0028; #100;
A = 16'h00BD; B = 16'h0029; #100;
A = 16'h00BD; B = 16'h002A; #100;
A = 16'h00BD; B = 16'h002B; #100;
A = 16'h00BD; B = 16'h002C; #100;
A = 16'h00BD; B = 16'h002D; #100;
A = 16'h00BD; B = 16'h002E; #100;
A = 16'h00BD; B = 16'h002F; #100;
A = 16'h00BD; B = 16'h0030; #100;
A = 16'h00BD; B = 16'h0031; #100;
A = 16'h00BD; B = 16'h0032; #100;
A = 16'h00BD; B = 16'h0033; #100;
A = 16'h00BD; B = 16'h0034; #100;
A = 16'h00BD; B = 16'h0035; #100;
A = 16'h00BD; B = 16'h0036; #100;
A = 16'h00BD; B = 16'h0037; #100;
A = 16'h00BD; B = 16'h0038; #100;
A = 16'h00BD; B = 16'h0039; #100;
A = 16'h00BD; B = 16'h003A; #100;
A = 16'h00BD; B = 16'h003B; #100;
A = 16'h00BD; B = 16'h003C; #100;
A = 16'h00BD; B = 16'h003D; #100;
A = 16'h00BD; B = 16'h003E; #100;
A = 16'h00BD; B = 16'h003F; #100;
A = 16'h00BD; B = 16'h0040; #100;
A = 16'h00BD; B = 16'h0041; #100;
A = 16'h00BD; B = 16'h0042; #100;
A = 16'h00BD; B = 16'h0043; #100;
A = 16'h00BD; B = 16'h0044; #100;
A = 16'h00BD; B = 16'h0045; #100;
A = 16'h00BD; B = 16'h0046; #100;
A = 16'h00BD; B = 16'h0047; #100;
A = 16'h00BD; B = 16'h0048; #100;
A = 16'h00BD; B = 16'h0049; #100;
A = 16'h00BD; B = 16'h004A; #100;
A = 16'h00BD; B = 16'h004B; #100;
A = 16'h00BD; B = 16'h004C; #100;
A = 16'h00BD; B = 16'h004D; #100;
A = 16'h00BD; B = 16'h004E; #100;
A = 16'h00BD; B = 16'h004F; #100;
A = 16'h00BD; B = 16'h0050; #100;
A = 16'h00BD; B = 16'h0051; #100;
A = 16'h00BD; B = 16'h0052; #100;
A = 16'h00BD; B = 16'h0053; #100;
A = 16'h00BD; B = 16'h0054; #100;
A = 16'h00BD; B = 16'h0055; #100;
A = 16'h00BD; B = 16'h0056; #100;
A = 16'h00BD; B = 16'h0057; #100;
A = 16'h00BD; B = 16'h0058; #100;
A = 16'h00BD; B = 16'h0059; #100;
A = 16'h00BD; B = 16'h005A; #100;
A = 16'h00BD; B = 16'h005B; #100;
A = 16'h00BD; B = 16'h005C; #100;
A = 16'h00BD; B = 16'h005D; #100;
A = 16'h00BD; B = 16'h005E; #100;
A = 16'h00BD; B = 16'h005F; #100;
A = 16'h00BD; B = 16'h0060; #100;
A = 16'h00BD; B = 16'h0061; #100;
A = 16'h00BD; B = 16'h0062; #100;
A = 16'h00BD; B = 16'h0063; #100;
A = 16'h00BD; B = 16'h0064; #100;
A = 16'h00BD; B = 16'h0065; #100;
A = 16'h00BD; B = 16'h0066; #100;
A = 16'h00BD; B = 16'h0067; #100;
A = 16'h00BD; B = 16'h0068; #100;
A = 16'h00BD; B = 16'h0069; #100;
A = 16'h00BD; B = 16'h006A; #100;
A = 16'h00BD; B = 16'h006B; #100;
A = 16'h00BD; B = 16'h006C; #100;
A = 16'h00BD; B = 16'h006D; #100;
A = 16'h00BD; B = 16'h006E; #100;
A = 16'h00BD; B = 16'h006F; #100;
A = 16'h00BD; B = 16'h0070; #100;
A = 16'h00BD; B = 16'h0071; #100;
A = 16'h00BD; B = 16'h0072; #100;
A = 16'h00BD; B = 16'h0073; #100;
A = 16'h00BD; B = 16'h0074; #100;
A = 16'h00BD; B = 16'h0075; #100;
A = 16'h00BD; B = 16'h0076; #100;
A = 16'h00BD; B = 16'h0077; #100;
A = 16'h00BD; B = 16'h0078; #100;
A = 16'h00BD; B = 16'h0079; #100;
A = 16'h00BD; B = 16'h007A; #100;
A = 16'h00BD; B = 16'h007B; #100;
A = 16'h00BD; B = 16'h007C; #100;
A = 16'h00BD; B = 16'h007D; #100;
A = 16'h00BD; B = 16'h007E; #100;
A = 16'h00BD; B = 16'h007F; #100;
A = 16'h00BD; B = 16'h0080; #100;
A = 16'h00BD; B = 16'h0081; #100;
A = 16'h00BD; B = 16'h0082; #100;
A = 16'h00BD; B = 16'h0083; #100;
A = 16'h00BD; B = 16'h0084; #100;
A = 16'h00BD; B = 16'h0085; #100;
A = 16'h00BD; B = 16'h0086; #100;
A = 16'h00BD; B = 16'h0087; #100;
A = 16'h00BD; B = 16'h0088; #100;
A = 16'h00BD; B = 16'h0089; #100;
A = 16'h00BD; B = 16'h008A; #100;
A = 16'h00BD; B = 16'h008B; #100;
A = 16'h00BD; B = 16'h008C; #100;
A = 16'h00BD; B = 16'h008D; #100;
A = 16'h00BD; B = 16'h008E; #100;
A = 16'h00BD; B = 16'h008F; #100;
A = 16'h00BD; B = 16'h0090; #100;
A = 16'h00BD; B = 16'h0091; #100;
A = 16'h00BD; B = 16'h0092; #100;
A = 16'h00BD; B = 16'h0093; #100;
A = 16'h00BD; B = 16'h0094; #100;
A = 16'h00BD; B = 16'h0095; #100;
A = 16'h00BD; B = 16'h0096; #100;
A = 16'h00BD; B = 16'h0097; #100;
A = 16'h00BD; B = 16'h0098; #100;
A = 16'h00BD; B = 16'h0099; #100;
A = 16'h00BD; B = 16'h009A; #100;
A = 16'h00BD; B = 16'h009B; #100;
A = 16'h00BD; B = 16'h009C; #100;
A = 16'h00BD; B = 16'h009D; #100;
A = 16'h00BD; B = 16'h009E; #100;
A = 16'h00BD; B = 16'h009F; #100;
A = 16'h00BD; B = 16'h00A0; #100;
A = 16'h00BD; B = 16'h00A1; #100;
A = 16'h00BD; B = 16'h00A2; #100;
A = 16'h00BD; B = 16'h00A3; #100;
A = 16'h00BD; B = 16'h00A4; #100;
A = 16'h00BD; B = 16'h00A5; #100;
A = 16'h00BD; B = 16'h00A6; #100;
A = 16'h00BD; B = 16'h00A7; #100;
A = 16'h00BD; B = 16'h00A8; #100;
A = 16'h00BD; B = 16'h00A9; #100;
A = 16'h00BD; B = 16'h00AA; #100;
A = 16'h00BD; B = 16'h00AB; #100;
A = 16'h00BD; B = 16'h00AC; #100;
A = 16'h00BD; B = 16'h00AD; #100;
A = 16'h00BD; B = 16'h00AE; #100;
A = 16'h00BD; B = 16'h00AF; #100;
A = 16'h00BD; B = 16'h00B0; #100;
A = 16'h00BD; B = 16'h00B1; #100;
A = 16'h00BD; B = 16'h00B2; #100;
A = 16'h00BD; B = 16'h00B3; #100;
A = 16'h00BD; B = 16'h00B4; #100;
A = 16'h00BD; B = 16'h00B5; #100;
A = 16'h00BD; B = 16'h00B6; #100;
A = 16'h00BD; B = 16'h00B7; #100;
A = 16'h00BD; B = 16'h00B8; #100;
A = 16'h00BD; B = 16'h00B9; #100;
A = 16'h00BD; B = 16'h00BA; #100;
A = 16'h00BD; B = 16'h00BB; #100;
A = 16'h00BD; B = 16'h00BC; #100;
A = 16'h00BD; B = 16'h00BD; #100;
A = 16'h00BD; B = 16'h00BE; #100;
A = 16'h00BD; B = 16'h00BF; #100;
A = 16'h00BD; B = 16'h00C0; #100;
A = 16'h00BD; B = 16'h00C1; #100;
A = 16'h00BD; B = 16'h00C2; #100;
A = 16'h00BD; B = 16'h00C3; #100;
A = 16'h00BD; B = 16'h00C4; #100;
A = 16'h00BD; B = 16'h00C5; #100;
A = 16'h00BD; B = 16'h00C6; #100;
A = 16'h00BD; B = 16'h00C7; #100;
A = 16'h00BD; B = 16'h00C8; #100;
A = 16'h00BD; B = 16'h00C9; #100;
A = 16'h00BD; B = 16'h00CA; #100;
A = 16'h00BD; B = 16'h00CB; #100;
A = 16'h00BD; B = 16'h00CC; #100;
A = 16'h00BD; B = 16'h00CD; #100;
A = 16'h00BD; B = 16'h00CE; #100;
A = 16'h00BD; B = 16'h00CF; #100;
A = 16'h00BD; B = 16'h00D0; #100;
A = 16'h00BD; B = 16'h00D1; #100;
A = 16'h00BD; B = 16'h00D2; #100;
A = 16'h00BD; B = 16'h00D3; #100;
A = 16'h00BD; B = 16'h00D4; #100;
A = 16'h00BD; B = 16'h00D5; #100;
A = 16'h00BD; B = 16'h00D6; #100;
A = 16'h00BD; B = 16'h00D7; #100;
A = 16'h00BD; B = 16'h00D8; #100;
A = 16'h00BD; B = 16'h00D9; #100;
A = 16'h00BD; B = 16'h00DA; #100;
A = 16'h00BD; B = 16'h00DB; #100;
A = 16'h00BD; B = 16'h00DC; #100;
A = 16'h00BD; B = 16'h00DD; #100;
A = 16'h00BD; B = 16'h00DE; #100;
A = 16'h00BD; B = 16'h00DF; #100;
A = 16'h00BD; B = 16'h00E0; #100;
A = 16'h00BD; B = 16'h00E1; #100;
A = 16'h00BD; B = 16'h00E2; #100;
A = 16'h00BD; B = 16'h00E3; #100;
A = 16'h00BD; B = 16'h00E4; #100;
A = 16'h00BD; B = 16'h00E5; #100;
A = 16'h00BD; B = 16'h00E6; #100;
A = 16'h00BD; B = 16'h00E7; #100;
A = 16'h00BD; B = 16'h00E8; #100;
A = 16'h00BD; B = 16'h00E9; #100;
A = 16'h00BD; B = 16'h00EA; #100;
A = 16'h00BD; B = 16'h00EB; #100;
A = 16'h00BD; B = 16'h00EC; #100;
A = 16'h00BD; B = 16'h00ED; #100;
A = 16'h00BD; B = 16'h00EE; #100;
A = 16'h00BD; B = 16'h00EF; #100;
A = 16'h00BD; B = 16'h00F0; #100;
A = 16'h00BD; B = 16'h00F1; #100;
A = 16'h00BD; B = 16'h00F2; #100;
A = 16'h00BD; B = 16'h00F3; #100;
A = 16'h00BD; B = 16'h00F4; #100;
A = 16'h00BD; B = 16'h00F5; #100;
A = 16'h00BD; B = 16'h00F6; #100;
A = 16'h00BD; B = 16'h00F7; #100;
A = 16'h00BD; B = 16'h00F8; #100;
A = 16'h00BD; B = 16'h00F9; #100;
A = 16'h00BD; B = 16'h00FA; #100;
A = 16'h00BD; B = 16'h00FB; #100;
A = 16'h00BD; B = 16'h00FC; #100;
A = 16'h00BD; B = 16'h00FD; #100;
A = 16'h00BD; B = 16'h00FE; #100;
A = 16'h00BD; B = 16'h00FF; #100;
A = 16'h00BE; B = 16'h000; #100;
A = 16'h00BE; B = 16'h001; #100;
A = 16'h00BE; B = 16'h002; #100;
A = 16'h00BE; B = 16'h003; #100;
A = 16'h00BE; B = 16'h004; #100;
A = 16'h00BE; B = 16'h005; #100;
A = 16'h00BE; B = 16'h006; #100;
A = 16'h00BE; B = 16'h007; #100;
A = 16'h00BE; B = 16'h008; #100;
A = 16'h00BE; B = 16'h009; #100;
A = 16'h00BE; B = 16'h00A; #100;
A = 16'h00BE; B = 16'h00B; #100;
A = 16'h00BE; B = 16'h00C; #100;
A = 16'h00BE; B = 16'h00D; #100;
A = 16'h00BE; B = 16'h00E; #100;
A = 16'h00BE; B = 16'h00F; #100;
A = 16'h00BE; B = 16'h0010; #100;
A = 16'h00BE; B = 16'h0011; #100;
A = 16'h00BE; B = 16'h0012; #100;
A = 16'h00BE; B = 16'h0013; #100;
A = 16'h00BE; B = 16'h0014; #100;
A = 16'h00BE; B = 16'h0015; #100;
A = 16'h00BE; B = 16'h0016; #100;
A = 16'h00BE; B = 16'h0017; #100;
A = 16'h00BE; B = 16'h0018; #100;
A = 16'h00BE; B = 16'h0019; #100;
A = 16'h00BE; B = 16'h001A; #100;
A = 16'h00BE; B = 16'h001B; #100;
A = 16'h00BE; B = 16'h001C; #100;
A = 16'h00BE; B = 16'h001D; #100;
A = 16'h00BE; B = 16'h001E; #100;
A = 16'h00BE; B = 16'h001F; #100;
A = 16'h00BE; B = 16'h0020; #100;
A = 16'h00BE; B = 16'h0021; #100;
A = 16'h00BE; B = 16'h0022; #100;
A = 16'h00BE; B = 16'h0023; #100;
A = 16'h00BE; B = 16'h0024; #100;
A = 16'h00BE; B = 16'h0025; #100;
A = 16'h00BE; B = 16'h0026; #100;
A = 16'h00BE; B = 16'h0027; #100;
A = 16'h00BE; B = 16'h0028; #100;
A = 16'h00BE; B = 16'h0029; #100;
A = 16'h00BE; B = 16'h002A; #100;
A = 16'h00BE; B = 16'h002B; #100;
A = 16'h00BE; B = 16'h002C; #100;
A = 16'h00BE; B = 16'h002D; #100;
A = 16'h00BE; B = 16'h002E; #100;
A = 16'h00BE; B = 16'h002F; #100;
A = 16'h00BE; B = 16'h0030; #100;
A = 16'h00BE; B = 16'h0031; #100;
A = 16'h00BE; B = 16'h0032; #100;
A = 16'h00BE; B = 16'h0033; #100;
A = 16'h00BE; B = 16'h0034; #100;
A = 16'h00BE; B = 16'h0035; #100;
A = 16'h00BE; B = 16'h0036; #100;
A = 16'h00BE; B = 16'h0037; #100;
A = 16'h00BE; B = 16'h0038; #100;
A = 16'h00BE; B = 16'h0039; #100;
A = 16'h00BE; B = 16'h003A; #100;
A = 16'h00BE; B = 16'h003B; #100;
A = 16'h00BE; B = 16'h003C; #100;
A = 16'h00BE; B = 16'h003D; #100;
A = 16'h00BE; B = 16'h003E; #100;
A = 16'h00BE; B = 16'h003F; #100;
A = 16'h00BE; B = 16'h0040; #100;
A = 16'h00BE; B = 16'h0041; #100;
A = 16'h00BE; B = 16'h0042; #100;
A = 16'h00BE; B = 16'h0043; #100;
A = 16'h00BE; B = 16'h0044; #100;
A = 16'h00BE; B = 16'h0045; #100;
A = 16'h00BE; B = 16'h0046; #100;
A = 16'h00BE; B = 16'h0047; #100;
A = 16'h00BE; B = 16'h0048; #100;
A = 16'h00BE; B = 16'h0049; #100;
A = 16'h00BE; B = 16'h004A; #100;
A = 16'h00BE; B = 16'h004B; #100;
A = 16'h00BE; B = 16'h004C; #100;
A = 16'h00BE; B = 16'h004D; #100;
A = 16'h00BE; B = 16'h004E; #100;
A = 16'h00BE; B = 16'h004F; #100;
A = 16'h00BE; B = 16'h0050; #100;
A = 16'h00BE; B = 16'h0051; #100;
A = 16'h00BE; B = 16'h0052; #100;
A = 16'h00BE; B = 16'h0053; #100;
A = 16'h00BE; B = 16'h0054; #100;
A = 16'h00BE; B = 16'h0055; #100;
A = 16'h00BE; B = 16'h0056; #100;
A = 16'h00BE; B = 16'h0057; #100;
A = 16'h00BE; B = 16'h0058; #100;
A = 16'h00BE; B = 16'h0059; #100;
A = 16'h00BE; B = 16'h005A; #100;
A = 16'h00BE; B = 16'h005B; #100;
A = 16'h00BE; B = 16'h005C; #100;
A = 16'h00BE; B = 16'h005D; #100;
A = 16'h00BE; B = 16'h005E; #100;
A = 16'h00BE; B = 16'h005F; #100;
A = 16'h00BE; B = 16'h0060; #100;
A = 16'h00BE; B = 16'h0061; #100;
A = 16'h00BE; B = 16'h0062; #100;
A = 16'h00BE; B = 16'h0063; #100;
A = 16'h00BE; B = 16'h0064; #100;
A = 16'h00BE; B = 16'h0065; #100;
A = 16'h00BE; B = 16'h0066; #100;
A = 16'h00BE; B = 16'h0067; #100;
A = 16'h00BE; B = 16'h0068; #100;
A = 16'h00BE; B = 16'h0069; #100;
A = 16'h00BE; B = 16'h006A; #100;
A = 16'h00BE; B = 16'h006B; #100;
A = 16'h00BE; B = 16'h006C; #100;
A = 16'h00BE; B = 16'h006D; #100;
A = 16'h00BE; B = 16'h006E; #100;
A = 16'h00BE; B = 16'h006F; #100;
A = 16'h00BE; B = 16'h0070; #100;
A = 16'h00BE; B = 16'h0071; #100;
A = 16'h00BE; B = 16'h0072; #100;
A = 16'h00BE; B = 16'h0073; #100;
A = 16'h00BE; B = 16'h0074; #100;
A = 16'h00BE; B = 16'h0075; #100;
A = 16'h00BE; B = 16'h0076; #100;
A = 16'h00BE; B = 16'h0077; #100;
A = 16'h00BE; B = 16'h0078; #100;
A = 16'h00BE; B = 16'h0079; #100;
A = 16'h00BE; B = 16'h007A; #100;
A = 16'h00BE; B = 16'h007B; #100;
A = 16'h00BE; B = 16'h007C; #100;
A = 16'h00BE; B = 16'h007D; #100;
A = 16'h00BE; B = 16'h007E; #100;
A = 16'h00BE; B = 16'h007F; #100;
A = 16'h00BE; B = 16'h0080; #100;
A = 16'h00BE; B = 16'h0081; #100;
A = 16'h00BE; B = 16'h0082; #100;
A = 16'h00BE; B = 16'h0083; #100;
A = 16'h00BE; B = 16'h0084; #100;
A = 16'h00BE; B = 16'h0085; #100;
A = 16'h00BE; B = 16'h0086; #100;
A = 16'h00BE; B = 16'h0087; #100;
A = 16'h00BE; B = 16'h0088; #100;
A = 16'h00BE; B = 16'h0089; #100;
A = 16'h00BE; B = 16'h008A; #100;
A = 16'h00BE; B = 16'h008B; #100;
A = 16'h00BE; B = 16'h008C; #100;
A = 16'h00BE; B = 16'h008D; #100;
A = 16'h00BE; B = 16'h008E; #100;
A = 16'h00BE; B = 16'h008F; #100;
A = 16'h00BE; B = 16'h0090; #100;
A = 16'h00BE; B = 16'h0091; #100;
A = 16'h00BE; B = 16'h0092; #100;
A = 16'h00BE; B = 16'h0093; #100;
A = 16'h00BE; B = 16'h0094; #100;
A = 16'h00BE; B = 16'h0095; #100;
A = 16'h00BE; B = 16'h0096; #100;
A = 16'h00BE; B = 16'h0097; #100;
A = 16'h00BE; B = 16'h0098; #100;
A = 16'h00BE; B = 16'h0099; #100;
A = 16'h00BE; B = 16'h009A; #100;
A = 16'h00BE; B = 16'h009B; #100;
A = 16'h00BE; B = 16'h009C; #100;
A = 16'h00BE; B = 16'h009D; #100;
A = 16'h00BE; B = 16'h009E; #100;
A = 16'h00BE; B = 16'h009F; #100;
A = 16'h00BE; B = 16'h00A0; #100;
A = 16'h00BE; B = 16'h00A1; #100;
A = 16'h00BE; B = 16'h00A2; #100;
A = 16'h00BE; B = 16'h00A3; #100;
A = 16'h00BE; B = 16'h00A4; #100;
A = 16'h00BE; B = 16'h00A5; #100;
A = 16'h00BE; B = 16'h00A6; #100;
A = 16'h00BE; B = 16'h00A7; #100;
A = 16'h00BE; B = 16'h00A8; #100;
A = 16'h00BE; B = 16'h00A9; #100;
A = 16'h00BE; B = 16'h00AA; #100;
A = 16'h00BE; B = 16'h00AB; #100;
A = 16'h00BE; B = 16'h00AC; #100;
A = 16'h00BE; B = 16'h00AD; #100;
A = 16'h00BE; B = 16'h00AE; #100;
A = 16'h00BE; B = 16'h00AF; #100;
A = 16'h00BE; B = 16'h00B0; #100;
A = 16'h00BE; B = 16'h00B1; #100;
A = 16'h00BE; B = 16'h00B2; #100;
A = 16'h00BE; B = 16'h00B3; #100;
A = 16'h00BE; B = 16'h00B4; #100;
A = 16'h00BE; B = 16'h00B5; #100;
A = 16'h00BE; B = 16'h00B6; #100;
A = 16'h00BE; B = 16'h00B7; #100;
A = 16'h00BE; B = 16'h00B8; #100;
A = 16'h00BE; B = 16'h00B9; #100;
A = 16'h00BE; B = 16'h00BA; #100;
A = 16'h00BE; B = 16'h00BB; #100;
A = 16'h00BE; B = 16'h00BC; #100;
A = 16'h00BE; B = 16'h00BD; #100;
A = 16'h00BE; B = 16'h00BE; #100;
A = 16'h00BE; B = 16'h00BF; #100;
A = 16'h00BE; B = 16'h00C0; #100;
A = 16'h00BE; B = 16'h00C1; #100;
A = 16'h00BE; B = 16'h00C2; #100;
A = 16'h00BE; B = 16'h00C3; #100;
A = 16'h00BE; B = 16'h00C4; #100;
A = 16'h00BE; B = 16'h00C5; #100;
A = 16'h00BE; B = 16'h00C6; #100;
A = 16'h00BE; B = 16'h00C7; #100;
A = 16'h00BE; B = 16'h00C8; #100;
A = 16'h00BE; B = 16'h00C9; #100;
A = 16'h00BE; B = 16'h00CA; #100;
A = 16'h00BE; B = 16'h00CB; #100;
A = 16'h00BE; B = 16'h00CC; #100;
A = 16'h00BE; B = 16'h00CD; #100;
A = 16'h00BE; B = 16'h00CE; #100;
A = 16'h00BE; B = 16'h00CF; #100;
A = 16'h00BE; B = 16'h00D0; #100;
A = 16'h00BE; B = 16'h00D1; #100;
A = 16'h00BE; B = 16'h00D2; #100;
A = 16'h00BE; B = 16'h00D3; #100;
A = 16'h00BE; B = 16'h00D4; #100;
A = 16'h00BE; B = 16'h00D5; #100;
A = 16'h00BE; B = 16'h00D6; #100;
A = 16'h00BE; B = 16'h00D7; #100;
A = 16'h00BE; B = 16'h00D8; #100;
A = 16'h00BE; B = 16'h00D9; #100;
A = 16'h00BE; B = 16'h00DA; #100;
A = 16'h00BE; B = 16'h00DB; #100;
A = 16'h00BE; B = 16'h00DC; #100;
A = 16'h00BE; B = 16'h00DD; #100;
A = 16'h00BE; B = 16'h00DE; #100;
A = 16'h00BE; B = 16'h00DF; #100;
A = 16'h00BE; B = 16'h00E0; #100;
A = 16'h00BE; B = 16'h00E1; #100;
A = 16'h00BE; B = 16'h00E2; #100;
A = 16'h00BE; B = 16'h00E3; #100;
A = 16'h00BE; B = 16'h00E4; #100;
A = 16'h00BE; B = 16'h00E5; #100;
A = 16'h00BE; B = 16'h00E6; #100;
A = 16'h00BE; B = 16'h00E7; #100;
A = 16'h00BE; B = 16'h00E8; #100;
A = 16'h00BE; B = 16'h00E9; #100;
A = 16'h00BE; B = 16'h00EA; #100;
A = 16'h00BE; B = 16'h00EB; #100;
A = 16'h00BE; B = 16'h00EC; #100;
A = 16'h00BE; B = 16'h00ED; #100;
A = 16'h00BE; B = 16'h00EE; #100;
A = 16'h00BE; B = 16'h00EF; #100;
A = 16'h00BE; B = 16'h00F0; #100;
A = 16'h00BE; B = 16'h00F1; #100;
A = 16'h00BE; B = 16'h00F2; #100;
A = 16'h00BE; B = 16'h00F3; #100;
A = 16'h00BE; B = 16'h00F4; #100;
A = 16'h00BE; B = 16'h00F5; #100;
A = 16'h00BE; B = 16'h00F6; #100;
A = 16'h00BE; B = 16'h00F7; #100;
A = 16'h00BE; B = 16'h00F8; #100;
A = 16'h00BE; B = 16'h00F9; #100;
A = 16'h00BE; B = 16'h00FA; #100;
A = 16'h00BE; B = 16'h00FB; #100;
A = 16'h00BE; B = 16'h00FC; #100;
A = 16'h00BE; B = 16'h00FD; #100;
A = 16'h00BE; B = 16'h00FE; #100;
A = 16'h00BE; B = 16'h00FF; #100;
A = 16'h00BF; B = 16'h000; #100;
A = 16'h00BF; B = 16'h001; #100;
A = 16'h00BF; B = 16'h002; #100;
A = 16'h00BF; B = 16'h003; #100;
A = 16'h00BF; B = 16'h004; #100;
A = 16'h00BF; B = 16'h005; #100;
A = 16'h00BF; B = 16'h006; #100;
A = 16'h00BF; B = 16'h007; #100;
A = 16'h00BF; B = 16'h008; #100;
A = 16'h00BF; B = 16'h009; #100;
A = 16'h00BF; B = 16'h00A; #100;
A = 16'h00BF; B = 16'h00B; #100;
A = 16'h00BF; B = 16'h00C; #100;
A = 16'h00BF; B = 16'h00D; #100;
A = 16'h00BF; B = 16'h00E; #100;
A = 16'h00BF; B = 16'h00F; #100;
A = 16'h00BF; B = 16'h0010; #100;
A = 16'h00BF; B = 16'h0011; #100;
A = 16'h00BF; B = 16'h0012; #100;
A = 16'h00BF; B = 16'h0013; #100;
A = 16'h00BF; B = 16'h0014; #100;
A = 16'h00BF; B = 16'h0015; #100;
A = 16'h00BF; B = 16'h0016; #100;
A = 16'h00BF; B = 16'h0017; #100;
A = 16'h00BF; B = 16'h0018; #100;
A = 16'h00BF; B = 16'h0019; #100;
A = 16'h00BF; B = 16'h001A; #100;
A = 16'h00BF; B = 16'h001B; #100;
A = 16'h00BF; B = 16'h001C; #100;
A = 16'h00BF; B = 16'h001D; #100;
A = 16'h00BF; B = 16'h001E; #100;
A = 16'h00BF; B = 16'h001F; #100;
A = 16'h00BF; B = 16'h0020; #100;
A = 16'h00BF; B = 16'h0021; #100;
A = 16'h00BF; B = 16'h0022; #100;
A = 16'h00BF; B = 16'h0023; #100;
A = 16'h00BF; B = 16'h0024; #100;
A = 16'h00BF; B = 16'h0025; #100;
A = 16'h00BF; B = 16'h0026; #100;
A = 16'h00BF; B = 16'h0027; #100;
A = 16'h00BF; B = 16'h0028; #100;
A = 16'h00BF; B = 16'h0029; #100;
A = 16'h00BF; B = 16'h002A; #100;
A = 16'h00BF; B = 16'h002B; #100;
A = 16'h00BF; B = 16'h002C; #100;
A = 16'h00BF; B = 16'h002D; #100;
A = 16'h00BF; B = 16'h002E; #100;
A = 16'h00BF; B = 16'h002F; #100;
A = 16'h00BF; B = 16'h0030; #100;
A = 16'h00BF; B = 16'h0031; #100;
A = 16'h00BF; B = 16'h0032; #100;
A = 16'h00BF; B = 16'h0033; #100;
A = 16'h00BF; B = 16'h0034; #100;
A = 16'h00BF; B = 16'h0035; #100;
A = 16'h00BF; B = 16'h0036; #100;
A = 16'h00BF; B = 16'h0037; #100;
A = 16'h00BF; B = 16'h0038; #100;
A = 16'h00BF; B = 16'h0039; #100;
A = 16'h00BF; B = 16'h003A; #100;
A = 16'h00BF; B = 16'h003B; #100;
A = 16'h00BF; B = 16'h003C; #100;
A = 16'h00BF; B = 16'h003D; #100;
A = 16'h00BF; B = 16'h003E; #100;
A = 16'h00BF; B = 16'h003F; #100;
A = 16'h00BF; B = 16'h0040; #100;
A = 16'h00BF; B = 16'h0041; #100;
A = 16'h00BF; B = 16'h0042; #100;
A = 16'h00BF; B = 16'h0043; #100;
A = 16'h00BF; B = 16'h0044; #100;
A = 16'h00BF; B = 16'h0045; #100;
A = 16'h00BF; B = 16'h0046; #100;
A = 16'h00BF; B = 16'h0047; #100;
A = 16'h00BF; B = 16'h0048; #100;
A = 16'h00BF; B = 16'h0049; #100;
A = 16'h00BF; B = 16'h004A; #100;
A = 16'h00BF; B = 16'h004B; #100;
A = 16'h00BF; B = 16'h004C; #100;
A = 16'h00BF; B = 16'h004D; #100;
A = 16'h00BF; B = 16'h004E; #100;
A = 16'h00BF; B = 16'h004F; #100;
A = 16'h00BF; B = 16'h0050; #100;
A = 16'h00BF; B = 16'h0051; #100;
A = 16'h00BF; B = 16'h0052; #100;
A = 16'h00BF; B = 16'h0053; #100;
A = 16'h00BF; B = 16'h0054; #100;
A = 16'h00BF; B = 16'h0055; #100;
A = 16'h00BF; B = 16'h0056; #100;
A = 16'h00BF; B = 16'h0057; #100;
A = 16'h00BF; B = 16'h0058; #100;
A = 16'h00BF; B = 16'h0059; #100;
A = 16'h00BF; B = 16'h005A; #100;
A = 16'h00BF; B = 16'h005B; #100;
A = 16'h00BF; B = 16'h005C; #100;
A = 16'h00BF; B = 16'h005D; #100;
A = 16'h00BF; B = 16'h005E; #100;
A = 16'h00BF; B = 16'h005F; #100;
A = 16'h00BF; B = 16'h0060; #100;
A = 16'h00BF; B = 16'h0061; #100;
A = 16'h00BF; B = 16'h0062; #100;
A = 16'h00BF; B = 16'h0063; #100;
A = 16'h00BF; B = 16'h0064; #100;
A = 16'h00BF; B = 16'h0065; #100;
A = 16'h00BF; B = 16'h0066; #100;
A = 16'h00BF; B = 16'h0067; #100;
A = 16'h00BF; B = 16'h0068; #100;
A = 16'h00BF; B = 16'h0069; #100;
A = 16'h00BF; B = 16'h006A; #100;
A = 16'h00BF; B = 16'h006B; #100;
A = 16'h00BF; B = 16'h006C; #100;
A = 16'h00BF; B = 16'h006D; #100;
A = 16'h00BF; B = 16'h006E; #100;
A = 16'h00BF; B = 16'h006F; #100;
A = 16'h00BF; B = 16'h0070; #100;
A = 16'h00BF; B = 16'h0071; #100;
A = 16'h00BF; B = 16'h0072; #100;
A = 16'h00BF; B = 16'h0073; #100;
A = 16'h00BF; B = 16'h0074; #100;
A = 16'h00BF; B = 16'h0075; #100;
A = 16'h00BF; B = 16'h0076; #100;
A = 16'h00BF; B = 16'h0077; #100;
A = 16'h00BF; B = 16'h0078; #100;
A = 16'h00BF; B = 16'h0079; #100;
A = 16'h00BF; B = 16'h007A; #100;
A = 16'h00BF; B = 16'h007B; #100;
A = 16'h00BF; B = 16'h007C; #100;
A = 16'h00BF; B = 16'h007D; #100;
A = 16'h00BF; B = 16'h007E; #100;
A = 16'h00BF; B = 16'h007F; #100;
A = 16'h00BF; B = 16'h0080; #100;
A = 16'h00BF; B = 16'h0081; #100;
A = 16'h00BF; B = 16'h0082; #100;
A = 16'h00BF; B = 16'h0083; #100;
A = 16'h00BF; B = 16'h0084; #100;
A = 16'h00BF; B = 16'h0085; #100;
A = 16'h00BF; B = 16'h0086; #100;
A = 16'h00BF; B = 16'h0087; #100;
A = 16'h00BF; B = 16'h0088; #100;
A = 16'h00BF; B = 16'h0089; #100;
A = 16'h00BF; B = 16'h008A; #100;
A = 16'h00BF; B = 16'h008B; #100;
A = 16'h00BF; B = 16'h008C; #100;
A = 16'h00BF; B = 16'h008D; #100;
A = 16'h00BF; B = 16'h008E; #100;
A = 16'h00BF; B = 16'h008F; #100;
A = 16'h00BF; B = 16'h0090; #100;
A = 16'h00BF; B = 16'h0091; #100;
A = 16'h00BF; B = 16'h0092; #100;
A = 16'h00BF; B = 16'h0093; #100;
A = 16'h00BF; B = 16'h0094; #100;
A = 16'h00BF; B = 16'h0095; #100;
A = 16'h00BF; B = 16'h0096; #100;
A = 16'h00BF; B = 16'h0097; #100;
A = 16'h00BF; B = 16'h0098; #100;
A = 16'h00BF; B = 16'h0099; #100;
A = 16'h00BF; B = 16'h009A; #100;
A = 16'h00BF; B = 16'h009B; #100;
A = 16'h00BF; B = 16'h009C; #100;
A = 16'h00BF; B = 16'h009D; #100;
A = 16'h00BF; B = 16'h009E; #100;
A = 16'h00BF; B = 16'h009F; #100;
A = 16'h00BF; B = 16'h00A0; #100;
A = 16'h00BF; B = 16'h00A1; #100;
A = 16'h00BF; B = 16'h00A2; #100;
A = 16'h00BF; B = 16'h00A3; #100;
A = 16'h00BF; B = 16'h00A4; #100;
A = 16'h00BF; B = 16'h00A5; #100;
A = 16'h00BF; B = 16'h00A6; #100;
A = 16'h00BF; B = 16'h00A7; #100;
A = 16'h00BF; B = 16'h00A8; #100;
A = 16'h00BF; B = 16'h00A9; #100;
A = 16'h00BF; B = 16'h00AA; #100;
A = 16'h00BF; B = 16'h00AB; #100;
A = 16'h00BF; B = 16'h00AC; #100;
A = 16'h00BF; B = 16'h00AD; #100;
A = 16'h00BF; B = 16'h00AE; #100;
A = 16'h00BF; B = 16'h00AF; #100;
A = 16'h00BF; B = 16'h00B0; #100;
A = 16'h00BF; B = 16'h00B1; #100;
A = 16'h00BF; B = 16'h00B2; #100;
A = 16'h00BF; B = 16'h00B3; #100;
A = 16'h00BF; B = 16'h00B4; #100;
A = 16'h00BF; B = 16'h00B5; #100;
A = 16'h00BF; B = 16'h00B6; #100;
A = 16'h00BF; B = 16'h00B7; #100;
A = 16'h00BF; B = 16'h00B8; #100;
A = 16'h00BF; B = 16'h00B9; #100;
A = 16'h00BF; B = 16'h00BA; #100;
A = 16'h00BF; B = 16'h00BB; #100;
A = 16'h00BF; B = 16'h00BC; #100;
A = 16'h00BF; B = 16'h00BD; #100;
A = 16'h00BF; B = 16'h00BE; #100;
A = 16'h00BF; B = 16'h00BF; #100;
A = 16'h00BF; B = 16'h00C0; #100;
A = 16'h00BF; B = 16'h00C1; #100;
A = 16'h00BF; B = 16'h00C2; #100;
A = 16'h00BF; B = 16'h00C3; #100;
A = 16'h00BF; B = 16'h00C4; #100;
A = 16'h00BF; B = 16'h00C5; #100;
A = 16'h00BF; B = 16'h00C6; #100;
A = 16'h00BF; B = 16'h00C7; #100;
A = 16'h00BF; B = 16'h00C8; #100;
A = 16'h00BF; B = 16'h00C9; #100;
A = 16'h00BF; B = 16'h00CA; #100;
A = 16'h00BF; B = 16'h00CB; #100;
A = 16'h00BF; B = 16'h00CC; #100;
A = 16'h00BF; B = 16'h00CD; #100;
A = 16'h00BF; B = 16'h00CE; #100;
A = 16'h00BF; B = 16'h00CF; #100;
A = 16'h00BF; B = 16'h00D0; #100;
A = 16'h00BF; B = 16'h00D1; #100;
A = 16'h00BF; B = 16'h00D2; #100;
A = 16'h00BF; B = 16'h00D3; #100;
A = 16'h00BF; B = 16'h00D4; #100;
A = 16'h00BF; B = 16'h00D5; #100;
A = 16'h00BF; B = 16'h00D6; #100;
A = 16'h00BF; B = 16'h00D7; #100;
A = 16'h00BF; B = 16'h00D8; #100;
A = 16'h00BF; B = 16'h00D9; #100;
A = 16'h00BF; B = 16'h00DA; #100;
A = 16'h00BF; B = 16'h00DB; #100;
A = 16'h00BF; B = 16'h00DC; #100;
A = 16'h00BF; B = 16'h00DD; #100;
A = 16'h00BF; B = 16'h00DE; #100;
A = 16'h00BF; B = 16'h00DF; #100;
A = 16'h00BF; B = 16'h00E0; #100;
A = 16'h00BF; B = 16'h00E1; #100;
A = 16'h00BF; B = 16'h00E2; #100;
A = 16'h00BF; B = 16'h00E3; #100;
A = 16'h00BF; B = 16'h00E4; #100;
A = 16'h00BF; B = 16'h00E5; #100;
A = 16'h00BF; B = 16'h00E6; #100;
A = 16'h00BF; B = 16'h00E7; #100;
A = 16'h00BF; B = 16'h00E8; #100;
A = 16'h00BF; B = 16'h00E9; #100;
A = 16'h00BF; B = 16'h00EA; #100;
A = 16'h00BF; B = 16'h00EB; #100;
A = 16'h00BF; B = 16'h00EC; #100;
A = 16'h00BF; B = 16'h00ED; #100;
A = 16'h00BF; B = 16'h00EE; #100;
A = 16'h00BF; B = 16'h00EF; #100;
A = 16'h00BF; B = 16'h00F0; #100;
A = 16'h00BF; B = 16'h00F1; #100;
A = 16'h00BF; B = 16'h00F2; #100;
A = 16'h00BF; B = 16'h00F3; #100;
A = 16'h00BF; B = 16'h00F4; #100;
A = 16'h00BF; B = 16'h00F5; #100;
A = 16'h00BF; B = 16'h00F6; #100;
A = 16'h00BF; B = 16'h00F7; #100;
A = 16'h00BF; B = 16'h00F8; #100;
A = 16'h00BF; B = 16'h00F9; #100;
A = 16'h00BF; B = 16'h00FA; #100;
A = 16'h00BF; B = 16'h00FB; #100;
A = 16'h00BF; B = 16'h00FC; #100;
A = 16'h00BF; B = 16'h00FD; #100;
A = 16'h00BF; B = 16'h00FE; #100;
A = 16'h00BF; B = 16'h00FF; #100;
A = 16'h00C0; B = 16'h000; #100;
A = 16'h00C0; B = 16'h001; #100;
A = 16'h00C0; B = 16'h002; #100;
A = 16'h00C0; B = 16'h003; #100;
A = 16'h00C0; B = 16'h004; #100;
A = 16'h00C0; B = 16'h005; #100;
A = 16'h00C0; B = 16'h006; #100;
A = 16'h00C0; B = 16'h007; #100;
A = 16'h00C0; B = 16'h008; #100;
A = 16'h00C0; B = 16'h009; #100;
A = 16'h00C0; B = 16'h00A; #100;
A = 16'h00C0; B = 16'h00B; #100;
A = 16'h00C0; B = 16'h00C; #100;
A = 16'h00C0; B = 16'h00D; #100;
A = 16'h00C0; B = 16'h00E; #100;
A = 16'h00C0; B = 16'h00F; #100;
A = 16'h00C0; B = 16'h0010; #100;
A = 16'h00C0; B = 16'h0011; #100;
A = 16'h00C0; B = 16'h0012; #100;
A = 16'h00C0; B = 16'h0013; #100;
A = 16'h00C0; B = 16'h0014; #100;
A = 16'h00C0; B = 16'h0015; #100;
A = 16'h00C0; B = 16'h0016; #100;
A = 16'h00C0; B = 16'h0017; #100;
A = 16'h00C0; B = 16'h0018; #100;
A = 16'h00C0; B = 16'h0019; #100;
A = 16'h00C0; B = 16'h001A; #100;
A = 16'h00C0; B = 16'h001B; #100;
A = 16'h00C0; B = 16'h001C; #100;
A = 16'h00C0; B = 16'h001D; #100;
A = 16'h00C0; B = 16'h001E; #100;
A = 16'h00C0; B = 16'h001F; #100;
A = 16'h00C0; B = 16'h0020; #100;
A = 16'h00C0; B = 16'h0021; #100;
A = 16'h00C0; B = 16'h0022; #100;
A = 16'h00C0; B = 16'h0023; #100;
A = 16'h00C0; B = 16'h0024; #100;
A = 16'h00C0; B = 16'h0025; #100;
A = 16'h00C0; B = 16'h0026; #100;
A = 16'h00C0; B = 16'h0027; #100;
A = 16'h00C0; B = 16'h0028; #100;
A = 16'h00C0; B = 16'h0029; #100;
A = 16'h00C0; B = 16'h002A; #100;
A = 16'h00C0; B = 16'h002B; #100;
A = 16'h00C0; B = 16'h002C; #100;
A = 16'h00C0; B = 16'h002D; #100;
A = 16'h00C0; B = 16'h002E; #100;
A = 16'h00C0; B = 16'h002F; #100;
A = 16'h00C0; B = 16'h0030; #100;
A = 16'h00C0; B = 16'h0031; #100;
A = 16'h00C0; B = 16'h0032; #100;
A = 16'h00C0; B = 16'h0033; #100;
A = 16'h00C0; B = 16'h0034; #100;
A = 16'h00C0; B = 16'h0035; #100;
A = 16'h00C0; B = 16'h0036; #100;
A = 16'h00C0; B = 16'h0037; #100;
A = 16'h00C0; B = 16'h0038; #100;
A = 16'h00C0; B = 16'h0039; #100;
A = 16'h00C0; B = 16'h003A; #100;
A = 16'h00C0; B = 16'h003B; #100;
A = 16'h00C0; B = 16'h003C; #100;
A = 16'h00C0; B = 16'h003D; #100;
A = 16'h00C0; B = 16'h003E; #100;
A = 16'h00C0; B = 16'h003F; #100;
A = 16'h00C0; B = 16'h0040; #100;
A = 16'h00C0; B = 16'h0041; #100;
A = 16'h00C0; B = 16'h0042; #100;
A = 16'h00C0; B = 16'h0043; #100;
A = 16'h00C0; B = 16'h0044; #100;
A = 16'h00C0; B = 16'h0045; #100;
A = 16'h00C0; B = 16'h0046; #100;
A = 16'h00C0; B = 16'h0047; #100;
A = 16'h00C0; B = 16'h0048; #100;
A = 16'h00C0; B = 16'h0049; #100;
A = 16'h00C0; B = 16'h004A; #100;
A = 16'h00C0; B = 16'h004B; #100;
A = 16'h00C0; B = 16'h004C; #100;
A = 16'h00C0; B = 16'h004D; #100;
A = 16'h00C0; B = 16'h004E; #100;
A = 16'h00C0; B = 16'h004F; #100;
A = 16'h00C0; B = 16'h0050; #100;
A = 16'h00C0; B = 16'h0051; #100;
A = 16'h00C0; B = 16'h0052; #100;
A = 16'h00C0; B = 16'h0053; #100;
A = 16'h00C0; B = 16'h0054; #100;
A = 16'h00C0; B = 16'h0055; #100;
A = 16'h00C0; B = 16'h0056; #100;
A = 16'h00C0; B = 16'h0057; #100;
A = 16'h00C0; B = 16'h0058; #100;
A = 16'h00C0; B = 16'h0059; #100;
A = 16'h00C0; B = 16'h005A; #100;
A = 16'h00C0; B = 16'h005B; #100;
A = 16'h00C0; B = 16'h005C; #100;
A = 16'h00C0; B = 16'h005D; #100;
A = 16'h00C0; B = 16'h005E; #100;
A = 16'h00C0; B = 16'h005F; #100;
A = 16'h00C0; B = 16'h0060; #100;
A = 16'h00C0; B = 16'h0061; #100;
A = 16'h00C0; B = 16'h0062; #100;
A = 16'h00C0; B = 16'h0063; #100;
A = 16'h00C0; B = 16'h0064; #100;
A = 16'h00C0; B = 16'h0065; #100;
A = 16'h00C0; B = 16'h0066; #100;
A = 16'h00C0; B = 16'h0067; #100;
A = 16'h00C0; B = 16'h0068; #100;
A = 16'h00C0; B = 16'h0069; #100;
A = 16'h00C0; B = 16'h006A; #100;
A = 16'h00C0; B = 16'h006B; #100;
A = 16'h00C0; B = 16'h006C; #100;
A = 16'h00C0; B = 16'h006D; #100;
A = 16'h00C0; B = 16'h006E; #100;
A = 16'h00C0; B = 16'h006F; #100;
A = 16'h00C0; B = 16'h0070; #100;
A = 16'h00C0; B = 16'h0071; #100;
A = 16'h00C0; B = 16'h0072; #100;
A = 16'h00C0; B = 16'h0073; #100;
A = 16'h00C0; B = 16'h0074; #100;
A = 16'h00C0; B = 16'h0075; #100;
A = 16'h00C0; B = 16'h0076; #100;
A = 16'h00C0; B = 16'h0077; #100;
A = 16'h00C0; B = 16'h0078; #100;
A = 16'h00C0; B = 16'h0079; #100;
A = 16'h00C0; B = 16'h007A; #100;
A = 16'h00C0; B = 16'h007B; #100;
A = 16'h00C0; B = 16'h007C; #100;
A = 16'h00C0; B = 16'h007D; #100;
A = 16'h00C0; B = 16'h007E; #100;
A = 16'h00C0; B = 16'h007F; #100;
A = 16'h00C0; B = 16'h0080; #100;
A = 16'h00C0; B = 16'h0081; #100;
A = 16'h00C0; B = 16'h0082; #100;
A = 16'h00C0; B = 16'h0083; #100;
A = 16'h00C0; B = 16'h0084; #100;
A = 16'h00C0; B = 16'h0085; #100;
A = 16'h00C0; B = 16'h0086; #100;
A = 16'h00C0; B = 16'h0087; #100;
A = 16'h00C0; B = 16'h0088; #100;
A = 16'h00C0; B = 16'h0089; #100;
A = 16'h00C0; B = 16'h008A; #100;
A = 16'h00C0; B = 16'h008B; #100;
A = 16'h00C0; B = 16'h008C; #100;
A = 16'h00C0; B = 16'h008D; #100;
A = 16'h00C0; B = 16'h008E; #100;
A = 16'h00C0; B = 16'h008F; #100;
A = 16'h00C0; B = 16'h0090; #100;
A = 16'h00C0; B = 16'h0091; #100;
A = 16'h00C0; B = 16'h0092; #100;
A = 16'h00C0; B = 16'h0093; #100;
A = 16'h00C0; B = 16'h0094; #100;
A = 16'h00C0; B = 16'h0095; #100;
A = 16'h00C0; B = 16'h0096; #100;
A = 16'h00C0; B = 16'h0097; #100;
A = 16'h00C0; B = 16'h0098; #100;
A = 16'h00C0; B = 16'h0099; #100;
A = 16'h00C0; B = 16'h009A; #100;
A = 16'h00C0; B = 16'h009B; #100;
A = 16'h00C0; B = 16'h009C; #100;
A = 16'h00C0; B = 16'h009D; #100;
A = 16'h00C0; B = 16'h009E; #100;
A = 16'h00C0; B = 16'h009F; #100;
A = 16'h00C0; B = 16'h00A0; #100;
A = 16'h00C0; B = 16'h00A1; #100;
A = 16'h00C0; B = 16'h00A2; #100;
A = 16'h00C0; B = 16'h00A3; #100;
A = 16'h00C0; B = 16'h00A4; #100;
A = 16'h00C0; B = 16'h00A5; #100;
A = 16'h00C0; B = 16'h00A6; #100;
A = 16'h00C0; B = 16'h00A7; #100;
A = 16'h00C0; B = 16'h00A8; #100;
A = 16'h00C0; B = 16'h00A9; #100;
A = 16'h00C0; B = 16'h00AA; #100;
A = 16'h00C0; B = 16'h00AB; #100;
A = 16'h00C0; B = 16'h00AC; #100;
A = 16'h00C0; B = 16'h00AD; #100;
A = 16'h00C0; B = 16'h00AE; #100;
A = 16'h00C0; B = 16'h00AF; #100;
A = 16'h00C0; B = 16'h00B0; #100;
A = 16'h00C0; B = 16'h00B1; #100;
A = 16'h00C0; B = 16'h00B2; #100;
A = 16'h00C0; B = 16'h00B3; #100;
A = 16'h00C0; B = 16'h00B4; #100;
A = 16'h00C0; B = 16'h00B5; #100;
A = 16'h00C0; B = 16'h00B6; #100;
A = 16'h00C0; B = 16'h00B7; #100;
A = 16'h00C0; B = 16'h00B8; #100;
A = 16'h00C0; B = 16'h00B9; #100;
A = 16'h00C0; B = 16'h00BA; #100;
A = 16'h00C0; B = 16'h00BB; #100;
A = 16'h00C0; B = 16'h00BC; #100;
A = 16'h00C0; B = 16'h00BD; #100;
A = 16'h00C0; B = 16'h00BE; #100;
A = 16'h00C0; B = 16'h00BF; #100;
A = 16'h00C0; B = 16'h00C0; #100;
A = 16'h00C0; B = 16'h00C1; #100;
A = 16'h00C0; B = 16'h00C2; #100;
A = 16'h00C0; B = 16'h00C3; #100;
A = 16'h00C0; B = 16'h00C4; #100;
A = 16'h00C0; B = 16'h00C5; #100;
A = 16'h00C0; B = 16'h00C6; #100;
A = 16'h00C0; B = 16'h00C7; #100;
A = 16'h00C0; B = 16'h00C8; #100;
A = 16'h00C0; B = 16'h00C9; #100;
A = 16'h00C0; B = 16'h00CA; #100;
A = 16'h00C0; B = 16'h00CB; #100;
A = 16'h00C0; B = 16'h00CC; #100;
A = 16'h00C0; B = 16'h00CD; #100;
A = 16'h00C0; B = 16'h00CE; #100;
A = 16'h00C0; B = 16'h00CF; #100;
A = 16'h00C0; B = 16'h00D0; #100;
A = 16'h00C0; B = 16'h00D1; #100;
A = 16'h00C0; B = 16'h00D2; #100;
A = 16'h00C0; B = 16'h00D3; #100;
A = 16'h00C0; B = 16'h00D4; #100;
A = 16'h00C0; B = 16'h00D5; #100;
A = 16'h00C0; B = 16'h00D6; #100;
A = 16'h00C0; B = 16'h00D7; #100;
A = 16'h00C0; B = 16'h00D8; #100;
A = 16'h00C0; B = 16'h00D9; #100;
A = 16'h00C0; B = 16'h00DA; #100;
A = 16'h00C0; B = 16'h00DB; #100;
A = 16'h00C0; B = 16'h00DC; #100;
A = 16'h00C0; B = 16'h00DD; #100;
A = 16'h00C0; B = 16'h00DE; #100;
A = 16'h00C0; B = 16'h00DF; #100;
A = 16'h00C0; B = 16'h00E0; #100;
A = 16'h00C0; B = 16'h00E1; #100;
A = 16'h00C0; B = 16'h00E2; #100;
A = 16'h00C0; B = 16'h00E3; #100;
A = 16'h00C0; B = 16'h00E4; #100;
A = 16'h00C0; B = 16'h00E5; #100;
A = 16'h00C0; B = 16'h00E6; #100;
A = 16'h00C0; B = 16'h00E7; #100;
A = 16'h00C0; B = 16'h00E8; #100;
A = 16'h00C0; B = 16'h00E9; #100;
A = 16'h00C0; B = 16'h00EA; #100;
A = 16'h00C0; B = 16'h00EB; #100;
A = 16'h00C0; B = 16'h00EC; #100;
A = 16'h00C0; B = 16'h00ED; #100;
A = 16'h00C0; B = 16'h00EE; #100;
A = 16'h00C0; B = 16'h00EF; #100;
A = 16'h00C0; B = 16'h00F0; #100;
A = 16'h00C0; B = 16'h00F1; #100;
A = 16'h00C0; B = 16'h00F2; #100;
A = 16'h00C0; B = 16'h00F3; #100;
A = 16'h00C0; B = 16'h00F4; #100;
A = 16'h00C0; B = 16'h00F5; #100;
A = 16'h00C0; B = 16'h00F6; #100;
A = 16'h00C0; B = 16'h00F7; #100;
A = 16'h00C0; B = 16'h00F8; #100;
A = 16'h00C0; B = 16'h00F9; #100;
A = 16'h00C0; B = 16'h00FA; #100;
A = 16'h00C0; B = 16'h00FB; #100;
A = 16'h00C0; B = 16'h00FC; #100;
A = 16'h00C0; B = 16'h00FD; #100;
A = 16'h00C0; B = 16'h00FE; #100;
A = 16'h00C0; B = 16'h00FF; #100;
A = 16'h00C1; B = 16'h000; #100;
A = 16'h00C1; B = 16'h001; #100;
A = 16'h00C1; B = 16'h002; #100;
A = 16'h00C1; B = 16'h003; #100;
A = 16'h00C1; B = 16'h004; #100;
A = 16'h00C1; B = 16'h005; #100;
A = 16'h00C1; B = 16'h006; #100;
A = 16'h00C1; B = 16'h007; #100;
A = 16'h00C1; B = 16'h008; #100;
A = 16'h00C1; B = 16'h009; #100;
A = 16'h00C1; B = 16'h00A; #100;
A = 16'h00C1; B = 16'h00B; #100;
A = 16'h00C1; B = 16'h00C; #100;
A = 16'h00C1; B = 16'h00D; #100;
A = 16'h00C1; B = 16'h00E; #100;
A = 16'h00C1; B = 16'h00F; #100;
A = 16'h00C1; B = 16'h0010; #100;
A = 16'h00C1; B = 16'h0011; #100;
A = 16'h00C1; B = 16'h0012; #100;
A = 16'h00C1; B = 16'h0013; #100;
A = 16'h00C1; B = 16'h0014; #100;
A = 16'h00C1; B = 16'h0015; #100;
A = 16'h00C1; B = 16'h0016; #100;
A = 16'h00C1; B = 16'h0017; #100;
A = 16'h00C1; B = 16'h0018; #100;
A = 16'h00C1; B = 16'h0019; #100;
A = 16'h00C1; B = 16'h001A; #100;
A = 16'h00C1; B = 16'h001B; #100;
A = 16'h00C1; B = 16'h001C; #100;
A = 16'h00C1; B = 16'h001D; #100;
A = 16'h00C1; B = 16'h001E; #100;
A = 16'h00C1; B = 16'h001F; #100;
A = 16'h00C1; B = 16'h0020; #100;
A = 16'h00C1; B = 16'h0021; #100;
A = 16'h00C1; B = 16'h0022; #100;
A = 16'h00C1; B = 16'h0023; #100;
A = 16'h00C1; B = 16'h0024; #100;
A = 16'h00C1; B = 16'h0025; #100;
A = 16'h00C1; B = 16'h0026; #100;
A = 16'h00C1; B = 16'h0027; #100;
A = 16'h00C1; B = 16'h0028; #100;
A = 16'h00C1; B = 16'h0029; #100;
A = 16'h00C1; B = 16'h002A; #100;
A = 16'h00C1; B = 16'h002B; #100;
A = 16'h00C1; B = 16'h002C; #100;
A = 16'h00C1; B = 16'h002D; #100;
A = 16'h00C1; B = 16'h002E; #100;
A = 16'h00C1; B = 16'h002F; #100;
A = 16'h00C1; B = 16'h0030; #100;
A = 16'h00C1; B = 16'h0031; #100;
A = 16'h00C1; B = 16'h0032; #100;
A = 16'h00C1; B = 16'h0033; #100;
A = 16'h00C1; B = 16'h0034; #100;
A = 16'h00C1; B = 16'h0035; #100;
A = 16'h00C1; B = 16'h0036; #100;
A = 16'h00C1; B = 16'h0037; #100;
A = 16'h00C1; B = 16'h0038; #100;
A = 16'h00C1; B = 16'h0039; #100;
A = 16'h00C1; B = 16'h003A; #100;
A = 16'h00C1; B = 16'h003B; #100;
A = 16'h00C1; B = 16'h003C; #100;
A = 16'h00C1; B = 16'h003D; #100;
A = 16'h00C1; B = 16'h003E; #100;
A = 16'h00C1; B = 16'h003F; #100;
A = 16'h00C1; B = 16'h0040; #100;
A = 16'h00C1; B = 16'h0041; #100;
A = 16'h00C1; B = 16'h0042; #100;
A = 16'h00C1; B = 16'h0043; #100;
A = 16'h00C1; B = 16'h0044; #100;
A = 16'h00C1; B = 16'h0045; #100;
A = 16'h00C1; B = 16'h0046; #100;
A = 16'h00C1; B = 16'h0047; #100;
A = 16'h00C1; B = 16'h0048; #100;
A = 16'h00C1; B = 16'h0049; #100;
A = 16'h00C1; B = 16'h004A; #100;
A = 16'h00C1; B = 16'h004B; #100;
A = 16'h00C1; B = 16'h004C; #100;
A = 16'h00C1; B = 16'h004D; #100;
A = 16'h00C1; B = 16'h004E; #100;
A = 16'h00C1; B = 16'h004F; #100;
A = 16'h00C1; B = 16'h0050; #100;
A = 16'h00C1; B = 16'h0051; #100;
A = 16'h00C1; B = 16'h0052; #100;
A = 16'h00C1; B = 16'h0053; #100;
A = 16'h00C1; B = 16'h0054; #100;
A = 16'h00C1; B = 16'h0055; #100;
A = 16'h00C1; B = 16'h0056; #100;
A = 16'h00C1; B = 16'h0057; #100;
A = 16'h00C1; B = 16'h0058; #100;
A = 16'h00C1; B = 16'h0059; #100;
A = 16'h00C1; B = 16'h005A; #100;
A = 16'h00C1; B = 16'h005B; #100;
A = 16'h00C1; B = 16'h005C; #100;
A = 16'h00C1; B = 16'h005D; #100;
A = 16'h00C1; B = 16'h005E; #100;
A = 16'h00C1; B = 16'h005F; #100;
A = 16'h00C1; B = 16'h0060; #100;
A = 16'h00C1; B = 16'h0061; #100;
A = 16'h00C1; B = 16'h0062; #100;
A = 16'h00C1; B = 16'h0063; #100;
A = 16'h00C1; B = 16'h0064; #100;
A = 16'h00C1; B = 16'h0065; #100;
A = 16'h00C1; B = 16'h0066; #100;
A = 16'h00C1; B = 16'h0067; #100;
A = 16'h00C1; B = 16'h0068; #100;
A = 16'h00C1; B = 16'h0069; #100;
A = 16'h00C1; B = 16'h006A; #100;
A = 16'h00C1; B = 16'h006B; #100;
A = 16'h00C1; B = 16'h006C; #100;
A = 16'h00C1; B = 16'h006D; #100;
A = 16'h00C1; B = 16'h006E; #100;
A = 16'h00C1; B = 16'h006F; #100;
A = 16'h00C1; B = 16'h0070; #100;
A = 16'h00C1; B = 16'h0071; #100;
A = 16'h00C1; B = 16'h0072; #100;
A = 16'h00C1; B = 16'h0073; #100;
A = 16'h00C1; B = 16'h0074; #100;
A = 16'h00C1; B = 16'h0075; #100;
A = 16'h00C1; B = 16'h0076; #100;
A = 16'h00C1; B = 16'h0077; #100;
A = 16'h00C1; B = 16'h0078; #100;
A = 16'h00C1; B = 16'h0079; #100;
A = 16'h00C1; B = 16'h007A; #100;
A = 16'h00C1; B = 16'h007B; #100;
A = 16'h00C1; B = 16'h007C; #100;
A = 16'h00C1; B = 16'h007D; #100;
A = 16'h00C1; B = 16'h007E; #100;
A = 16'h00C1; B = 16'h007F; #100;
A = 16'h00C1; B = 16'h0080; #100;
A = 16'h00C1; B = 16'h0081; #100;
A = 16'h00C1; B = 16'h0082; #100;
A = 16'h00C1; B = 16'h0083; #100;
A = 16'h00C1; B = 16'h0084; #100;
A = 16'h00C1; B = 16'h0085; #100;
A = 16'h00C1; B = 16'h0086; #100;
A = 16'h00C1; B = 16'h0087; #100;
A = 16'h00C1; B = 16'h0088; #100;
A = 16'h00C1; B = 16'h0089; #100;
A = 16'h00C1; B = 16'h008A; #100;
A = 16'h00C1; B = 16'h008B; #100;
A = 16'h00C1; B = 16'h008C; #100;
A = 16'h00C1; B = 16'h008D; #100;
A = 16'h00C1; B = 16'h008E; #100;
A = 16'h00C1; B = 16'h008F; #100;
A = 16'h00C1; B = 16'h0090; #100;
A = 16'h00C1; B = 16'h0091; #100;
A = 16'h00C1; B = 16'h0092; #100;
A = 16'h00C1; B = 16'h0093; #100;
A = 16'h00C1; B = 16'h0094; #100;
A = 16'h00C1; B = 16'h0095; #100;
A = 16'h00C1; B = 16'h0096; #100;
A = 16'h00C1; B = 16'h0097; #100;
A = 16'h00C1; B = 16'h0098; #100;
A = 16'h00C1; B = 16'h0099; #100;
A = 16'h00C1; B = 16'h009A; #100;
A = 16'h00C1; B = 16'h009B; #100;
A = 16'h00C1; B = 16'h009C; #100;
A = 16'h00C1; B = 16'h009D; #100;
A = 16'h00C1; B = 16'h009E; #100;
A = 16'h00C1; B = 16'h009F; #100;
A = 16'h00C1; B = 16'h00A0; #100;
A = 16'h00C1; B = 16'h00A1; #100;
A = 16'h00C1; B = 16'h00A2; #100;
A = 16'h00C1; B = 16'h00A3; #100;
A = 16'h00C1; B = 16'h00A4; #100;
A = 16'h00C1; B = 16'h00A5; #100;
A = 16'h00C1; B = 16'h00A6; #100;
A = 16'h00C1; B = 16'h00A7; #100;
A = 16'h00C1; B = 16'h00A8; #100;
A = 16'h00C1; B = 16'h00A9; #100;
A = 16'h00C1; B = 16'h00AA; #100;
A = 16'h00C1; B = 16'h00AB; #100;
A = 16'h00C1; B = 16'h00AC; #100;
A = 16'h00C1; B = 16'h00AD; #100;
A = 16'h00C1; B = 16'h00AE; #100;
A = 16'h00C1; B = 16'h00AF; #100;
A = 16'h00C1; B = 16'h00B0; #100;
A = 16'h00C1; B = 16'h00B1; #100;
A = 16'h00C1; B = 16'h00B2; #100;
A = 16'h00C1; B = 16'h00B3; #100;
A = 16'h00C1; B = 16'h00B4; #100;
A = 16'h00C1; B = 16'h00B5; #100;
A = 16'h00C1; B = 16'h00B6; #100;
A = 16'h00C1; B = 16'h00B7; #100;
A = 16'h00C1; B = 16'h00B8; #100;
A = 16'h00C1; B = 16'h00B9; #100;
A = 16'h00C1; B = 16'h00BA; #100;
A = 16'h00C1; B = 16'h00BB; #100;
A = 16'h00C1; B = 16'h00BC; #100;
A = 16'h00C1; B = 16'h00BD; #100;
A = 16'h00C1; B = 16'h00BE; #100;
A = 16'h00C1; B = 16'h00BF; #100;
A = 16'h00C1; B = 16'h00C0; #100;
A = 16'h00C1; B = 16'h00C1; #100;
A = 16'h00C1; B = 16'h00C2; #100;
A = 16'h00C1; B = 16'h00C3; #100;
A = 16'h00C1; B = 16'h00C4; #100;
A = 16'h00C1; B = 16'h00C5; #100;
A = 16'h00C1; B = 16'h00C6; #100;
A = 16'h00C1; B = 16'h00C7; #100;
A = 16'h00C1; B = 16'h00C8; #100;
A = 16'h00C1; B = 16'h00C9; #100;
A = 16'h00C1; B = 16'h00CA; #100;
A = 16'h00C1; B = 16'h00CB; #100;
A = 16'h00C1; B = 16'h00CC; #100;
A = 16'h00C1; B = 16'h00CD; #100;
A = 16'h00C1; B = 16'h00CE; #100;
A = 16'h00C1; B = 16'h00CF; #100;
A = 16'h00C1; B = 16'h00D0; #100;
A = 16'h00C1; B = 16'h00D1; #100;
A = 16'h00C1; B = 16'h00D2; #100;
A = 16'h00C1; B = 16'h00D3; #100;
A = 16'h00C1; B = 16'h00D4; #100;
A = 16'h00C1; B = 16'h00D5; #100;
A = 16'h00C1; B = 16'h00D6; #100;
A = 16'h00C1; B = 16'h00D7; #100;
A = 16'h00C1; B = 16'h00D8; #100;
A = 16'h00C1; B = 16'h00D9; #100;
A = 16'h00C1; B = 16'h00DA; #100;
A = 16'h00C1; B = 16'h00DB; #100;
A = 16'h00C1; B = 16'h00DC; #100;
A = 16'h00C1; B = 16'h00DD; #100;
A = 16'h00C1; B = 16'h00DE; #100;
A = 16'h00C1; B = 16'h00DF; #100;
A = 16'h00C1; B = 16'h00E0; #100;
A = 16'h00C1; B = 16'h00E1; #100;
A = 16'h00C1; B = 16'h00E2; #100;
A = 16'h00C1; B = 16'h00E3; #100;
A = 16'h00C1; B = 16'h00E4; #100;
A = 16'h00C1; B = 16'h00E5; #100;
A = 16'h00C1; B = 16'h00E6; #100;
A = 16'h00C1; B = 16'h00E7; #100;
A = 16'h00C1; B = 16'h00E8; #100;
A = 16'h00C1; B = 16'h00E9; #100;
A = 16'h00C1; B = 16'h00EA; #100;
A = 16'h00C1; B = 16'h00EB; #100;
A = 16'h00C1; B = 16'h00EC; #100;
A = 16'h00C1; B = 16'h00ED; #100;
A = 16'h00C1; B = 16'h00EE; #100;
A = 16'h00C1; B = 16'h00EF; #100;
A = 16'h00C1; B = 16'h00F0; #100;
A = 16'h00C1; B = 16'h00F1; #100;
A = 16'h00C1; B = 16'h00F2; #100;
A = 16'h00C1; B = 16'h00F3; #100;
A = 16'h00C1; B = 16'h00F4; #100;
A = 16'h00C1; B = 16'h00F5; #100;
A = 16'h00C1; B = 16'h00F6; #100;
A = 16'h00C1; B = 16'h00F7; #100;
A = 16'h00C1; B = 16'h00F8; #100;
A = 16'h00C1; B = 16'h00F9; #100;
A = 16'h00C1; B = 16'h00FA; #100;
A = 16'h00C1; B = 16'h00FB; #100;
A = 16'h00C1; B = 16'h00FC; #100;
A = 16'h00C1; B = 16'h00FD; #100;
A = 16'h00C1; B = 16'h00FE; #100;
A = 16'h00C1; B = 16'h00FF; #100;
A = 16'h00C2; B = 16'h000; #100;
A = 16'h00C2; B = 16'h001; #100;
A = 16'h00C2; B = 16'h002; #100;
A = 16'h00C2; B = 16'h003; #100;
A = 16'h00C2; B = 16'h004; #100;
A = 16'h00C2; B = 16'h005; #100;
A = 16'h00C2; B = 16'h006; #100;
A = 16'h00C2; B = 16'h007; #100;
A = 16'h00C2; B = 16'h008; #100;
A = 16'h00C2; B = 16'h009; #100;
A = 16'h00C2; B = 16'h00A; #100;
A = 16'h00C2; B = 16'h00B; #100;
A = 16'h00C2; B = 16'h00C; #100;
A = 16'h00C2; B = 16'h00D; #100;
A = 16'h00C2; B = 16'h00E; #100;
A = 16'h00C2; B = 16'h00F; #100;
A = 16'h00C2; B = 16'h0010; #100;
A = 16'h00C2; B = 16'h0011; #100;
A = 16'h00C2; B = 16'h0012; #100;
A = 16'h00C2; B = 16'h0013; #100;
A = 16'h00C2; B = 16'h0014; #100;
A = 16'h00C2; B = 16'h0015; #100;
A = 16'h00C2; B = 16'h0016; #100;
A = 16'h00C2; B = 16'h0017; #100;
A = 16'h00C2; B = 16'h0018; #100;
A = 16'h00C2; B = 16'h0019; #100;
A = 16'h00C2; B = 16'h001A; #100;
A = 16'h00C2; B = 16'h001B; #100;
A = 16'h00C2; B = 16'h001C; #100;
A = 16'h00C2; B = 16'h001D; #100;
A = 16'h00C2; B = 16'h001E; #100;
A = 16'h00C2; B = 16'h001F; #100;
A = 16'h00C2; B = 16'h0020; #100;
A = 16'h00C2; B = 16'h0021; #100;
A = 16'h00C2; B = 16'h0022; #100;
A = 16'h00C2; B = 16'h0023; #100;
A = 16'h00C2; B = 16'h0024; #100;
A = 16'h00C2; B = 16'h0025; #100;
A = 16'h00C2; B = 16'h0026; #100;
A = 16'h00C2; B = 16'h0027; #100;
A = 16'h00C2; B = 16'h0028; #100;
A = 16'h00C2; B = 16'h0029; #100;
A = 16'h00C2; B = 16'h002A; #100;
A = 16'h00C2; B = 16'h002B; #100;
A = 16'h00C2; B = 16'h002C; #100;
A = 16'h00C2; B = 16'h002D; #100;
A = 16'h00C2; B = 16'h002E; #100;
A = 16'h00C2; B = 16'h002F; #100;
A = 16'h00C2; B = 16'h0030; #100;
A = 16'h00C2; B = 16'h0031; #100;
A = 16'h00C2; B = 16'h0032; #100;
A = 16'h00C2; B = 16'h0033; #100;
A = 16'h00C2; B = 16'h0034; #100;
A = 16'h00C2; B = 16'h0035; #100;
A = 16'h00C2; B = 16'h0036; #100;
A = 16'h00C2; B = 16'h0037; #100;
A = 16'h00C2; B = 16'h0038; #100;
A = 16'h00C2; B = 16'h0039; #100;
A = 16'h00C2; B = 16'h003A; #100;
A = 16'h00C2; B = 16'h003B; #100;
A = 16'h00C2; B = 16'h003C; #100;
A = 16'h00C2; B = 16'h003D; #100;
A = 16'h00C2; B = 16'h003E; #100;
A = 16'h00C2; B = 16'h003F; #100;
A = 16'h00C2; B = 16'h0040; #100;
A = 16'h00C2; B = 16'h0041; #100;
A = 16'h00C2; B = 16'h0042; #100;
A = 16'h00C2; B = 16'h0043; #100;
A = 16'h00C2; B = 16'h0044; #100;
A = 16'h00C2; B = 16'h0045; #100;
A = 16'h00C2; B = 16'h0046; #100;
A = 16'h00C2; B = 16'h0047; #100;
A = 16'h00C2; B = 16'h0048; #100;
A = 16'h00C2; B = 16'h0049; #100;
A = 16'h00C2; B = 16'h004A; #100;
A = 16'h00C2; B = 16'h004B; #100;
A = 16'h00C2; B = 16'h004C; #100;
A = 16'h00C2; B = 16'h004D; #100;
A = 16'h00C2; B = 16'h004E; #100;
A = 16'h00C2; B = 16'h004F; #100;
A = 16'h00C2; B = 16'h0050; #100;
A = 16'h00C2; B = 16'h0051; #100;
A = 16'h00C2; B = 16'h0052; #100;
A = 16'h00C2; B = 16'h0053; #100;
A = 16'h00C2; B = 16'h0054; #100;
A = 16'h00C2; B = 16'h0055; #100;
A = 16'h00C2; B = 16'h0056; #100;
A = 16'h00C2; B = 16'h0057; #100;
A = 16'h00C2; B = 16'h0058; #100;
A = 16'h00C2; B = 16'h0059; #100;
A = 16'h00C2; B = 16'h005A; #100;
A = 16'h00C2; B = 16'h005B; #100;
A = 16'h00C2; B = 16'h005C; #100;
A = 16'h00C2; B = 16'h005D; #100;
A = 16'h00C2; B = 16'h005E; #100;
A = 16'h00C2; B = 16'h005F; #100;
A = 16'h00C2; B = 16'h0060; #100;
A = 16'h00C2; B = 16'h0061; #100;
A = 16'h00C2; B = 16'h0062; #100;
A = 16'h00C2; B = 16'h0063; #100;
A = 16'h00C2; B = 16'h0064; #100;
A = 16'h00C2; B = 16'h0065; #100;
A = 16'h00C2; B = 16'h0066; #100;
A = 16'h00C2; B = 16'h0067; #100;
A = 16'h00C2; B = 16'h0068; #100;
A = 16'h00C2; B = 16'h0069; #100;
A = 16'h00C2; B = 16'h006A; #100;
A = 16'h00C2; B = 16'h006B; #100;
A = 16'h00C2; B = 16'h006C; #100;
A = 16'h00C2; B = 16'h006D; #100;
A = 16'h00C2; B = 16'h006E; #100;
A = 16'h00C2; B = 16'h006F; #100;
A = 16'h00C2; B = 16'h0070; #100;
A = 16'h00C2; B = 16'h0071; #100;
A = 16'h00C2; B = 16'h0072; #100;
A = 16'h00C2; B = 16'h0073; #100;
A = 16'h00C2; B = 16'h0074; #100;
A = 16'h00C2; B = 16'h0075; #100;
A = 16'h00C2; B = 16'h0076; #100;
A = 16'h00C2; B = 16'h0077; #100;
A = 16'h00C2; B = 16'h0078; #100;
A = 16'h00C2; B = 16'h0079; #100;
A = 16'h00C2; B = 16'h007A; #100;
A = 16'h00C2; B = 16'h007B; #100;
A = 16'h00C2; B = 16'h007C; #100;
A = 16'h00C2; B = 16'h007D; #100;
A = 16'h00C2; B = 16'h007E; #100;
A = 16'h00C2; B = 16'h007F; #100;
A = 16'h00C2; B = 16'h0080; #100;
A = 16'h00C2; B = 16'h0081; #100;
A = 16'h00C2; B = 16'h0082; #100;
A = 16'h00C2; B = 16'h0083; #100;
A = 16'h00C2; B = 16'h0084; #100;
A = 16'h00C2; B = 16'h0085; #100;
A = 16'h00C2; B = 16'h0086; #100;
A = 16'h00C2; B = 16'h0087; #100;
A = 16'h00C2; B = 16'h0088; #100;
A = 16'h00C2; B = 16'h0089; #100;
A = 16'h00C2; B = 16'h008A; #100;
A = 16'h00C2; B = 16'h008B; #100;
A = 16'h00C2; B = 16'h008C; #100;
A = 16'h00C2; B = 16'h008D; #100;
A = 16'h00C2; B = 16'h008E; #100;
A = 16'h00C2; B = 16'h008F; #100;
A = 16'h00C2; B = 16'h0090; #100;
A = 16'h00C2; B = 16'h0091; #100;
A = 16'h00C2; B = 16'h0092; #100;
A = 16'h00C2; B = 16'h0093; #100;
A = 16'h00C2; B = 16'h0094; #100;
A = 16'h00C2; B = 16'h0095; #100;
A = 16'h00C2; B = 16'h0096; #100;
A = 16'h00C2; B = 16'h0097; #100;
A = 16'h00C2; B = 16'h0098; #100;
A = 16'h00C2; B = 16'h0099; #100;
A = 16'h00C2; B = 16'h009A; #100;
A = 16'h00C2; B = 16'h009B; #100;
A = 16'h00C2; B = 16'h009C; #100;
A = 16'h00C2; B = 16'h009D; #100;
A = 16'h00C2; B = 16'h009E; #100;
A = 16'h00C2; B = 16'h009F; #100;
A = 16'h00C2; B = 16'h00A0; #100;
A = 16'h00C2; B = 16'h00A1; #100;
A = 16'h00C2; B = 16'h00A2; #100;
A = 16'h00C2; B = 16'h00A3; #100;
A = 16'h00C2; B = 16'h00A4; #100;
A = 16'h00C2; B = 16'h00A5; #100;
A = 16'h00C2; B = 16'h00A6; #100;
A = 16'h00C2; B = 16'h00A7; #100;
A = 16'h00C2; B = 16'h00A8; #100;
A = 16'h00C2; B = 16'h00A9; #100;
A = 16'h00C2; B = 16'h00AA; #100;
A = 16'h00C2; B = 16'h00AB; #100;
A = 16'h00C2; B = 16'h00AC; #100;
A = 16'h00C2; B = 16'h00AD; #100;
A = 16'h00C2; B = 16'h00AE; #100;
A = 16'h00C2; B = 16'h00AF; #100;
A = 16'h00C2; B = 16'h00B0; #100;
A = 16'h00C2; B = 16'h00B1; #100;
A = 16'h00C2; B = 16'h00B2; #100;
A = 16'h00C2; B = 16'h00B3; #100;
A = 16'h00C2; B = 16'h00B4; #100;
A = 16'h00C2; B = 16'h00B5; #100;
A = 16'h00C2; B = 16'h00B6; #100;
A = 16'h00C2; B = 16'h00B7; #100;
A = 16'h00C2; B = 16'h00B8; #100;
A = 16'h00C2; B = 16'h00B9; #100;
A = 16'h00C2; B = 16'h00BA; #100;
A = 16'h00C2; B = 16'h00BB; #100;
A = 16'h00C2; B = 16'h00BC; #100;
A = 16'h00C2; B = 16'h00BD; #100;
A = 16'h00C2; B = 16'h00BE; #100;
A = 16'h00C2; B = 16'h00BF; #100;
A = 16'h00C2; B = 16'h00C0; #100;
A = 16'h00C2; B = 16'h00C1; #100;
A = 16'h00C2; B = 16'h00C2; #100;
A = 16'h00C2; B = 16'h00C3; #100;
A = 16'h00C2; B = 16'h00C4; #100;
A = 16'h00C2; B = 16'h00C5; #100;
A = 16'h00C2; B = 16'h00C6; #100;
A = 16'h00C2; B = 16'h00C7; #100;
A = 16'h00C2; B = 16'h00C8; #100;
A = 16'h00C2; B = 16'h00C9; #100;
A = 16'h00C2; B = 16'h00CA; #100;
A = 16'h00C2; B = 16'h00CB; #100;
A = 16'h00C2; B = 16'h00CC; #100;
A = 16'h00C2; B = 16'h00CD; #100;
A = 16'h00C2; B = 16'h00CE; #100;
A = 16'h00C2; B = 16'h00CF; #100;
A = 16'h00C2; B = 16'h00D0; #100;
A = 16'h00C2; B = 16'h00D1; #100;
A = 16'h00C2; B = 16'h00D2; #100;
A = 16'h00C2; B = 16'h00D3; #100;
A = 16'h00C2; B = 16'h00D4; #100;
A = 16'h00C2; B = 16'h00D5; #100;
A = 16'h00C2; B = 16'h00D6; #100;
A = 16'h00C2; B = 16'h00D7; #100;
A = 16'h00C2; B = 16'h00D8; #100;
A = 16'h00C2; B = 16'h00D9; #100;
A = 16'h00C2; B = 16'h00DA; #100;
A = 16'h00C2; B = 16'h00DB; #100;
A = 16'h00C2; B = 16'h00DC; #100;
A = 16'h00C2; B = 16'h00DD; #100;
A = 16'h00C2; B = 16'h00DE; #100;
A = 16'h00C2; B = 16'h00DF; #100;
A = 16'h00C2; B = 16'h00E0; #100;
A = 16'h00C2; B = 16'h00E1; #100;
A = 16'h00C2; B = 16'h00E2; #100;
A = 16'h00C2; B = 16'h00E3; #100;
A = 16'h00C2; B = 16'h00E4; #100;
A = 16'h00C2; B = 16'h00E5; #100;
A = 16'h00C2; B = 16'h00E6; #100;
A = 16'h00C2; B = 16'h00E7; #100;
A = 16'h00C2; B = 16'h00E8; #100;
A = 16'h00C2; B = 16'h00E9; #100;
A = 16'h00C2; B = 16'h00EA; #100;
A = 16'h00C2; B = 16'h00EB; #100;
A = 16'h00C2; B = 16'h00EC; #100;
A = 16'h00C2; B = 16'h00ED; #100;
A = 16'h00C2; B = 16'h00EE; #100;
A = 16'h00C2; B = 16'h00EF; #100;
A = 16'h00C2; B = 16'h00F0; #100;
A = 16'h00C2; B = 16'h00F1; #100;
A = 16'h00C2; B = 16'h00F2; #100;
A = 16'h00C2; B = 16'h00F3; #100;
A = 16'h00C2; B = 16'h00F4; #100;
A = 16'h00C2; B = 16'h00F5; #100;
A = 16'h00C2; B = 16'h00F6; #100;
A = 16'h00C2; B = 16'h00F7; #100;
A = 16'h00C2; B = 16'h00F8; #100;
A = 16'h00C2; B = 16'h00F9; #100;
A = 16'h00C2; B = 16'h00FA; #100;
A = 16'h00C2; B = 16'h00FB; #100;
A = 16'h00C2; B = 16'h00FC; #100;
A = 16'h00C2; B = 16'h00FD; #100;
A = 16'h00C2; B = 16'h00FE; #100;
A = 16'h00C2; B = 16'h00FF; #100;
A = 16'h00C3; B = 16'h000; #100;
A = 16'h00C3; B = 16'h001; #100;
A = 16'h00C3; B = 16'h002; #100;
A = 16'h00C3; B = 16'h003; #100;
A = 16'h00C3; B = 16'h004; #100;
A = 16'h00C3; B = 16'h005; #100;
A = 16'h00C3; B = 16'h006; #100;
A = 16'h00C3; B = 16'h007; #100;
A = 16'h00C3; B = 16'h008; #100;
A = 16'h00C3; B = 16'h009; #100;
A = 16'h00C3; B = 16'h00A; #100;
A = 16'h00C3; B = 16'h00B; #100;
A = 16'h00C3; B = 16'h00C; #100;
A = 16'h00C3; B = 16'h00D; #100;
A = 16'h00C3; B = 16'h00E; #100;
A = 16'h00C3; B = 16'h00F; #100;
A = 16'h00C3; B = 16'h0010; #100;
A = 16'h00C3; B = 16'h0011; #100;
A = 16'h00C3; B = 16'h0012; #100;
A = 16'h00C3; B = 16'h0013; #100;
A = 16'h00C3; B = 16'h0014; #100;
A = 16'h00C3; B = 16'h0015; #100;
A = 16'h00C3; B = 16'h0016; #100;
A = 16'h00C3; B = 16'h0017; #100;
A = 16'h00C3; B = 16'h0018; #100;
A = 16'h00C3; B = 16'h0019; #100;
A = 16'h00C3; B = 16'h001A; #100;
A = 16'h00C3; B = 16'h001B; #100;
A = 16'h00C3; B = 16'h001C; #100;
A = 16'h00C3; B = 16'h001D; #100;
A = 16'h00C3; B = 16'h001E; #100;
A = 16'h00C3; B = 16'h001F; #100;
A = 16'h00C3; B = 16'h0020; #100;
A = 16'h00C3; B = 16'h0021; #100;
A = 16'h00C3; B = 16'h0022; #100;
A = 16'h00C3; B = 16'h0023; #100;
A = 16'h00C3; B = 16'h0024; #100;
A = 16'h00C3; B = 16'h0025; #100;
A = 16'h00C3; B = 16'h0026; #100;
A = 16'h00C3; B = 16'h0027; #100;
A = 16'h00C3; B = 16'h0028; #100;
A = 16'h00C3; B = 16'h0029; #100;
A = 16'h00C3; B = 16'h002A; #100;
A = 16'h00C3; B = 16'h002B; #100;
A = 16'h00C3; B = 16'h002C; #100;
A = 16'h00C3; B = 16'h002D; #100;
A = 16'h00C3; B = 16'h002E; #100;
A = 16'h00C3; B = 16'h002F; #100;
A = 16'h00C3; B = 16'h0030; #100;
A = 16'h00C3; B = 16'h0031; #100;
A = 16'h00C3; B = 16'h0032; #100;
A = 16'h00C3; B = 16'h0033; #100;
A = 16'h00C3; B = 16'h0034; #100;
A = 16'h00C3; B = 16'h0035; #100;
A = 16'h00C3; B = 16'h0036; #100;
A = 16'h00C3; B = 16'h0037; #100;
A = 16'h00C3; B = 16'h0038; #100;
A = 16'h00C3; B = 16'h0039; #100;
A = 16'h00C3; B = 16'h003A; #100;
A = 16'h00C3; B = 16'h003B; #100;
A = 16'h00C3; B = 16'h003C; #100;
A = 16'h00C3; B = 16'h003D; #100;
A = 16'h00C3; B = 16'h003E; #100;
A = 16'h00C3; B = 16'h003F; #100;
A = 16'h00C3; B = 16'h0040; #100;
A = 16'h00C3; B = 16'h0041; #100;
A = 16'h00C3; B = 16'h0042; #100;
A = 16'h00C3; B = 16'h0043; #100;
A = 16'h00C3; B = 16'h0044; #100;
A = 16'h00C3; B = 16'h0045; #100;
A = 16'h00C3; B = 16'h0046; #100;
A = 16'h00C3; B = 16'h0047; #100;
A = 16'h00C3; B = 16'h0048; #100;
A = 16'h00C3; B = 16'h0049; #100;
A = 16'h00C3; B = 16'h004A; #100;
A = 16'h00C3; B = 16'h004B; #100;
A = 16'h00C3; B = 16'h004C; #100;
A = 16'h00C3; B = 16'h004D; #100;
A = 16'h00C3; B = 16'h004E; #100;
A = 16'h00C3; B = 16'h004F; #100;
A = 16'h00C3; B = 16'h0050; #100;
A = 16'h00C3; B = 16'h0051; #100;
A = 16'h00C3; B = 16'h0052; #100;
A = 16'h00C3; B = 16'h0053; #100;
A = 16'h00C3; B = 16'h0054; #100;
A = 16'h00C3; B = 16'h0055; #100;
A = 16'h00C3; B = 16'h0056; #100;
A = 16'h00C3; B = 16'h0057; #100;
A = 16'h00C3; B = 16'h0058; #100;
A = 16'h00C3; B = 16'h0059; #100;
A = 16'h00C3; B = 16'h005A; #100;
A = 16'h00C3; B = 16'h005B; #100;
A = 16'h00C3; B = 16'h005C; #100;
A = 16'h00C3; B = 16'h005D; #100;
A = 16'h00C3; B = 16'h005E; #100;
A = 16'h00C3; B = 16'h005F; #100;
A = 16'h00C3; B = 16'h0060; #100;
A = 16'h00C3; B = 16'h0061; #100;
A = 16'h00C3; B = 16'h0062; #100;
A = 16'h00C3; B = 16'h0063; #100;
A = 16'h00C3; B = 16'h0064; #100;
A = 16'h00C3; B = 16'h0065; #100;
A = 16'h00C3; B = 16'h0066; #100;
A = 16'h00C3; B = 16'h0067; #100;
A = 16'h00C3; B = 16'h0068; #100;
A = 16'h00C3; B = 16'h0069; #100;
A = 16'h00C3; B = 16'h006A; #100;
A = 16'h00C3; B = 16'h006B; #100;
A = 16'h00C3; B = 16'h006C; #100;
A = 16'h00C3; B = 16'h006D; #100;
A = 16'h00C3; B = 16'h006E; #100;
A = 16'h00C3; B = 16'h006F; #100;
A = 16'h00C3; B = 16'h0070; #100;
A = 16'h00C3; B = 16'h0071; #100;
A = 16'h00C3; B = 16'h0072; #100;
A = 16'h00C3; B = 16'h0073; #100;
A = 16'h00C3; B = 16'h0074; #100;
A = 16'h00C3; B = 16'h0075; #100;
A = 16'h00C3; B = 16'h0076; #100;
A = 16'h00C3; B = 16'h0077; #100;
A = 16'h00C3; B = 16'h0078; #100;
A = 16'h00C3; B = 16'h0079; #100;
A = 16'h00C3; B = 16'h007A; #100;
A = 16'h00C3; B = 16'h007B; #100;
A = 16'h00C3; B = 16'h007C; #100;
A = 16'h00C3; B = 16'h007D; #100;
A = 16'h00C3; B = 16'h007E; #100;
A = 16'h00C3; B = 16'h007F; #100;
A = 16'h00C3; B = 16'h0080; #100;
A = 16'h00C3; B = 16'h0081; #100;
A = 16'h00C3; B = 16'h0082; #100;
A = 16'h00C3; B = 16'h0083; #100;
A = 16'h00C3; B = 16'h0084; #100;
A = 16'h00C3; B = 16'h0085; #100;
A = 16'h00C3; B = 16'h0086; #100;
A = 16'h00C3; B = 16'h0087; #100;
A = 16'h00C3; B = 16'h0088; #100;
A = 16'h00C3; B = 16'h0089; #100;
A = 16'h00C3; B = 16'h008A; #100;
A = 16'h00C3; B = 16'h008B; #100;
A = 16'h00C3; B = 16'h008C; #100;
A = 16'h00C3; B = 16'h008D; #100;
A = 16'h00C3; B = 16'h008E; #100;
A = 16'h00C3; B = 16'h008F; #100;
A = 16'h00C3; B = 16'h0090; #100;
A = 16'h00C3; B = 16'h0091; #100;
A = 16'h00C3; B = 16'h0092; #100;
A = 16'h00C3; B = 16'h0093; #100;
A = 16'h00C3; B = 16'h0094; #100;
A = 16'h00C3; B = 16'h0095; #100;
A = 16'h00C3; B = 16'h0096; #100;
A = 16'h00C3; B = 16'h0097; #100;
A = 16'h00C3; B = 16'h0098; #100;
A = 16'h00C3; B = 16'h0099; #100;
A = 16'h00C3; B = 16'h009A; #100;
A = 16'h00C3; B = 16'h009B; #100;
A = 16'h00C3; B = 16'h009C; #100;
A = 16'h00C3; B = 16'h009D; #100;
A = 16'h00C3; B = 16'h009E; #100;
A = 16'h00C3; B = 16'h009F; #100;
A = 16'h00C3; B = 16'h00A0; #100;
A = 16'h00C3; B = 16'h00A1; #100;
A = 16'h00C3; B = 16'h00A2; #100;
A = 16'h00C3; B = 16'h00A3; #100;
A = 16'h00C3; B = 16'h00A4; #100;
A = 16'h00C3; B = 16'h00A5; #100;
A = 16'h00C3; B = 16'h00A6; #100;
A = 16'h00C3; B = 16'h00A7; #100;
A = 16'h00C3; B = 16'h00A8; #100;
A = 16'h00C3; B = 16'h00A9; #100;
A = 16'h00C3; B = 16'h00AA; #100;
A = 16'h00C3; B = 16'h00AB; #100;
A = 16'h00C3; B = 16'h00AC; #100;
A = 16'h00C3; B = 16'h00AD; #100;
A = 16'h00C3; B = 16'h00AE; #100;
A = 16'h00C3; B = 16'h00AF; #100;
A = 16'h00C3; B = 16'h00B0; #100;
A = 16'h00C3; B = 16'h00B1; #100;
A = 16'h00C3; B = 16'h00B2; #100;
A = 16'h00C3; B = 16'h00B3; #100;
A = 16'h00C3; B = 16'h00B4; #100;
A = 16'h00C3; B = 16'h00B5; #100;
A = 16'h00C3; B = 16'h00B6; #100;
A = 16'h00C3; B = 16'h00B7; #100;
A = 16'h00C3; B = 16'h00B8; #100;
A = 16'h00C3; B = 16'h00B9; #100;
A = 16'h00C3; B = 16'h00BA; #100;
A = 16'h00C3; B = 16'h00BB; #100;
A = 16'h00C3; B = 16'h00BC; #100;
A = 16'h00C3; B = 16'h00BD; #100;
A = 16'h00C3; B = 16'h00BE; #100;
A = 16'h00C3; B = 16'h00BF; #100;
A = 16'h00C3; B = 16'h00C0; #100;
A = 16'h00C3; B = 16'h00C1; #100;
A = 16'h00C3; B = 16'h00C2; #100;
A = 16'h00C3; B = 16'h00C3; #100;
A = 16'h00C3; B = 16'h00C4; #100;
A = 16'h00C3; B = 16'h00C5; #100;
A = 16'h00C3; B = 16'h00C6; #100;
A = 16'h00C3; B = 16'h00C7; #100;
A = 16'h00C3; B = 16'h00C8; #100;
A = 16'h00C3; B = 16'h00C9; #100;
A = 16'h00C3; B = 16'h00CA; #100;
A = 16'h00C3; B = 16'h00CB; #100;
A = 16'h00C3; B = 16'h00CC; #100;
A = 16'h00C3; B = 16'h00CD; #100;
A = 16'h00C3; B = 16'h00CE; #100;
A = 16'h00C3; B = 16'h00CF; #100;
A = 16'h00C3; B = 16'h00D0; #100;
A = 16'h00C3; B = 16'h00D1; #100;
A = 16'h00C3; B = 16'h00D2; #100;
A = 16'h00C3; B = 16'h00D3; #100;
A = 16'h00C3; B = 16'h00D4; #100;
A = 16'h00C3; B = 16'h00D5; #100;
A = 16'h00C3; B = 16'h00D6; #100;
A = 16'h00C3; B = 16'h00D7; #100;
A = 16'h00C3; B = 16'h00D8; #100;
A = 16'h00C3; B = 16'h00D9; #100;
A = 16'h00C3; B = 16'h00DA; #100;
A = 16'h00C3; B = 16'h00DB; #100;
A = 16'h00C3; B = 16'h00DC; #100;
A = 16'h00C3; B = 16'h00DD; #100;
A = 16'h00C3; B = 16'h00DE; #100;
A = 16'h00C3; B = 16'h00DF; #100;
A = 16'h00C3; B = 16'h00E0; #100;
A = 16'h00C3; B = 16'h00E1; #100;
A = 16'h00C3; B = 16'h00E2; #100;
A = 16'h00C3; B = 16'h00E3; #100;
A = 16'h00C3; B = 16'h00E4; #100;
A = 16'h00C3; B = 16'h00E5; #100;
A = 16'h00C3; B = 16'h00E6; #100;
A = 16'h00C3; B = 16'h00E7; #100;
A = 16'h00C3; B = 16'h00E8; #100;
A = 16'h00C3; B = 16'h00E9; #100;
A = 16'h00C3; B = 16'h00EA; #100;
A = 16'h00C3; B = 16'h00EB; #100;
A = 16'h00C3; B = 16'h00EC; #100;
A = 16'h00C3; B = 16'h00ED; #100;
A = 16'h00C3; B = 16'h00EE; #100;
A = 16'h00C3; B = 16'h00EF; #100;
A = 16'h00C3; B = 16'h00F0; #100;
A = 16'h00C3; B = 16'h00F1; #100;
A = 16'h00C3; B = 16'h00F2; #100;
A = 16'h00C3; B = 16'h00F3; #100;
A = 16'h00C3; B = 16'h00F4; #100;
A = 16'h00C3; B = 16'h00F5; #100;
A = 16'h00C3; B = 16'h00F6; #100;
A = 16'h00C3; B = 16'h00F7; #100;
A = 16'h00C3; B = 16'h00F8; #100;
A = 16'h00C3; B = 16'h00F9; #100;
A = 16'h00C3; B = 16'h00FA; #100;
A = 16'h00C3; B = 16'h00FB; #100;
A = 16'h00C3; B = 16'h00FC; #100;
A = 16'h00C3; B = 16'h00FD; #100;
A = 16'h00C3; B = 16'h00FE; #100;
A = 16'h00C3; B = 16'h00FF; #100;
A = 16'h00C4; B = 16'h000; #100;
A = 16'h00C4; B = 16'h001; #100;
A = 16'h00C4; B = 16'h002; #100;
A = 16'h00C4; B = 16'h003; #100;
A = 16'h00C4; B = 16'h004; #100;
A = 16'h00C4; B = 16'h005; #100;
A = 16'h00C4; B = 16'h006; #100;
A = 16'h00C4; B = 16'h007; #100;
A = 16'h00C4; B = 16'h008; #100;
A = 16'h00C4; B = 16'h009; #100;
A = 16'h00C4; B = 16'h00A; #100;
A = 16'h00C4; B = 16'h00B; #100;
A = 16'h00C4; B = 16'h00C; #100;
A = 16'h00C4; B = 16'h00D; #100;
A = 16'h00C4; B = 16'h00E; #100;
A = 16'h00C4; B = 16'h00F; #100;
A = 16'h00C4; B = 16'h0010; #100;
A = 16'h00C4; B = 16'h0011; #100;
A = 16'h00C4; B = 16'h0012; #100;
A = 16'h00C4; B = 16'h0013; #100;
A = 16'h00C4; B = 16'h0014; #100;
A = 16'h00C4; B = 16'h0015; #100;
A = 16'h00C4; B = 16'h0016; #100;
A = 16'h00C4; B = 16'h0017; #100;
A = 16'h00C4; B = 16'h0018; #100;
A = 16'h00C4; B = 16'h0019; #100;
A = 16'h00C4; B = 16'h001A; #100;
A = 16'h00C4; B = 16'h001B; #100;
A = 16'h00C4; B = 16'h001C; #100;
A = 16'h00C4; B = 16'h001D; #100;
A = 16'h00C4; B = 16'h001E; #100;
A = 16'h00C4; B = 16'h001F; #100;
A = 16'h00C4; B = 16'h0020; #100;
A = 16'h00C4; B = 16'h0021; #100;
A = 16'h00C4; B = 16'h0022; #100;
A = 16'h00C4; B = 16'h0023; #100;
A = 16'h00C4; B = 16'h0024; #100;
A = 16'h00C4; B = 16'h0025; #100;
A = 16'h00C4; B = 16'h0026; #100;
A = 16'h00C4; B = 16'h0027; #100;
A = 16'h00C4; B = 16'h0028; #100;
A = 16'h00C4; B = 16'h0029; #100;
A = 16'h00C4; B = 16'h002A; #100;
A = 16'h00C4; B = 16'h002B; #100;
A = 16'h00C4; B = 16'h002C; #100;
A = 16'h00C4; B = 16'h002D; #100;
A = 16'h00C4; B = 16'h002E; #100;
A = 16'h00C4; B = 16'h002F; #100;
A = 16'h00C4; B = 16'h0030; #100;
A = 16'h00C4; B = 16'h0031; #100;
A = 16'h00C4; B = 16'h0032; #100;
A = 16'h00C4; B = 16'h0033; #100;
A = 16'h00C4; B = 16'h0034; #100;
A = 16'h00C4; B = 16'h0035; #100;
A = 16'h00C4; B = 16'h0036; #100;
A = 16'h00C4; B = 16'h0037; #100;
A = 16'h00C4; B = 16'h0038; #100;
A = 16'h00C4; B = 16'h0039; #100;
A = 16'h00C4; B = 16'h003A; #100;
A = 16'h00C4; B = 16'h003B; #100;
A = 16'h00C4; B = 16'h003C; #100;
A = 16'h00C4; B = 16'h003D; #100;
A = 16'h00C4; B = 16'h003E; #100;
A = 16'h00C4; B = 16'h003F; #100;
A = 16'h00C4; B = 16'h0040; #100;
A = 16'h00C4; B = 16'h0041; #100;
A = 16'h00C4; B = 16'h0042; #100;
A = 16'h00C4; B = 16'h0043; #100;
A = 16'h00C4; B = 16'h0044; #100;
A = 16'h00C4; B = 16'h0045; #100;
A = 16'h00C4; B = 16'h0046; #100;
A = 16'h00C4; B = 16'h0047; #100;
A = 16'h00C4; B = 16'h0048; #100;
A = 16'h00C4; B = 16'h0049; #100;
A = 16'h00C4; B = 16'h004A; #100;
A = 16'h00C4; B = 16'h004B; #100;
A = 16'h00C4; B = 16'h004C; #100;
A = 16'h00C4; B = 16'h004D; #100;
A = 16'h00C4; B = 16'h004E; #100;
A = 16'h00C4; B = 16'h004F; #100;
A = 16'h00C4; B = 16'h0050; #100;
A = 16'h00C4; B = 16'h0051; #100;
A = 16'h00C4; B = 16'h0052; #100;
A = 16'h00C4; B = 16'h0053; #100;
A = 16'h00C4; B = 16'h0054; #100;
A = 16'h00C4; B = 16'h0055; #100;
A = 16'h00C4; B = 16'h0056; #100;
A = 16'h00C4; B = 16'h0057; #100;
A = 16'h00C4; B = 16'h0058; #100;
A = 16'h00C4; B = 16'h0059; #100;
A = 16'h00C4; B = 16'h005A; #100;
A = 16'h00C4; B = 16'h005B; #100;
A = 16'h00C4; B = 16'h005C; #100;
A = 16'h00C4; B = 16'h005D; #100;
A = 16'h00C4; B = 16'h005E; #100;
A = 16'h00C4; B = 16'h005F; #100;
A = 16'h00C4; B = 16'h0060; #100;
A = 16'h00C4; B = 16'h0061; #100;
A = 16'h00C4; B = 16'h0062; #100;
A = 16'h00C4; B = 16'h0063; #100;
A = 16'h00C4; B = 16'h0064; #100;
A = 16'h00C4; B = 16'h0065; #100;
A = 16'h00C4; B = 16'h0066; #100;
A = 16'h00C4; B = 16'h0067; #100;
A = 16'h00C4; B = 16'h0068; #100;
A = 16'h00C4; B = 16'h0069; #100;
A = 16'h00C4; B = 16'h006A; #100;
A = 16'h00C4; B = 16'h006B; #100;
A = 16'h00C4; B = 16'h006C; #100;
A = 16'h00C4; B = 16'h006D; #100;
A = 16'h00C4; B = 16'h006E; #100;
A = 16'h00C4; B = 16'h006F; #100;
A = 16'h00C4; B = 16'h0070; #100;
A = 16'h00C4; B = 16'h0071; #100;
A = 16'h00C4; B = 16'h0072; #100;
A = 16'h00C4; B = 16'h0073; #100;
A = 16'h00C4; B = 16'h0074; #100;
A = 16'h00C4; B = 16'h0075; #100;
A = 16'h00C4; B = 16'h0076; #100;
A = 16'h00C4; B = 16'h0077; #100;
A = 16'h00C4; B = 16'h0078; #100;
A = 16'h00C4; B = 16'h0079; #100;
A = 16'h00C4; B = 16'h007A; #100;
A = 16'h00C4; B = 16'h007B; #100;
A = 16'h00C4; B = 16'h007C; #100;
A = 16'h00C4; B = 16'h007D; #100;
A = 16'h00C4; B = 16'h007E; #100;
A = 16'h00C4; B = 16'h007F; #100;
A = 16'h00C4; B = 16'h0080; #100;
A = 16'h00C4; B = 16'h0081; #100;
A = 16'h00C4; B = 16'h0082; #100;
A = 16'h00C4; B = 16'h0083; #100;
A = 16'h00C4; B = 16'h0084; #100;
A = 16'h00C4; B = 16'h0085; #100;
A = 16'h00C4; B = 16'h0086; #100;
A = 16'h00C4; B = 16'h0087; #100;
A = 16'h00C4; B = 16'h0088; #100;
A = 16'h00C4; B = 16'h0089; #100;
A = 16'h00C4; B = 16'h008A; #100;
A = 16'h00C4; B = 16'h008B; #100;
A = 16'h00C4; B = 16'h008C; #100;
A = 16'h00C4; B = 16'h008D; #100;
A = 16'h00C4; B = 16'h008E; #100;
A = 16'h00C4; B = 16'h008F; #100;
A = 16'h00C4; B = 16'h0090; #100;
A = 16'h00C4; B = 16'h0091; #100;
A = 16'h00C4; B = 16'h0092; #100;
A = 16'h00C4; B = 16'h0093; #100;
A = 16'h00C4; B = 16'h0094; #100;
A = 16'h00C4; B = 16'h0095; #100;
A = 16'h00C4; B = 16'h0096; #100;
A = 16'h00C4; B = 16'h0097; #100;
A = 16'h00C4; B = 16'h0098; #100;
A = 16'h00C4; B = 16'h0099; #100;
A = 16'h00C4; B = 16'h009A; #100;
A = 16'h00C4; B = 16'h009B; #100;
A = 16'h00C4; B = 16'h009C; #100;
A = 16'h00C4; B = 16'h009D; #100;
A = 16'h00C4; B = 16'h009E; #100;
A = 16'h00C4; B = 16'h009F; #100;
A = 16'h00C4; B = 16'h00A0; #100;
A = 16'h00C4; B = 16'h00A1; #100;
A = 16'h00C4; B = 16'h00A2; #100;
A = 16'h00C4; B = 16'h00A3; #100;
A = 16'h00C4; B = 16'h00A4; #100;
A = 16'h00C4; B = 16'h00A5; #100;
A = 16'h00C4; B = 16'h00A6; #100;
A = 16'h00C4; B = 16'h00A7; #100;
A = 16'h00C4; B = 16'h00A8; #100;
A = 16'h00C4; B = 16'h00A9; #100;
A = 16'h00C4; B = 16'h00AA; #100;
A = 16'h00C4; B = 16'h00AB; #100;
A = 16'h00C4; B = 16'h00AC; #100;
A = 16'h00C4; B = 16'h00AD; #100;
A = 16'h00C4; B = 16'h00AE; #100;
A = 16'h00C4; B = 16'h00AF; #100;
A = 16'h00C4; B = 16'h00B0; #100;
A = 16'h00C4; B = 16'h00B1; #100;
A = 16'h00C4; B = 16'h00B2; #100;
A = 16'h00C4; B = 16'h00B3; #100;
A = 16'h00C4; B = 16'h00B4; #100;
A = 16'h00C4; B = 16'h00B5; #100;
A = 16'h00C4; B = 16'h00B6; #100;
A = 16'h00C4; B = 16'h00B7; #100;
A = 16'h00C4; B = 16'h00B8; #100;
A = 16'h00C4; B = 16'h00B9; #100;
A = 16'h00C4; B = 16'h00BA; #100;
A = 16'h00C4; B = 16'h00BB; #100;
A = 16'h00C4; B = 16'h00BC; #100;
A = 16'h00C4; B = 16'h00BD; #100;
A = 16'h00C4; B = 16'h00BE; #100;
A = 16'h00C4; B = 16'h00BF; #100;
A = 16'h00C4; B = 16'h00C0; #100;
A = 16'h00C4; B = 16'h00C1; #100;
A = 16'h00C4; B = 16'h00C2; #100;
A = 16'h00C4; B = 16'h00C3; #100;
A = 16'h00C4; B = 16'h00C4; #100;
A = 16'h00C4; B = 16'h00C5; #100;
A = 16'h00C4; B = 16'h00C6; #100;
A = 16'h00C4; B = 16'h00C7; #100;
A = 16'h00C4; B = 16'h00C8; #100;
A = 16'h00C4; B = 16'h00C9; #100;
A = 16'h00C4; B = 16'h00CA; #100;
A = 16'h00C4; B = 16'h00CB; #100;
A = 16'h00C4; B = 16'h00CC; #100;
A = 16'h00C4; B = 16'h00CD; #100;
A = 16'h00C4; B = 16'h00CE; #100;
A = 16'h00C4; B = 16'h00CF; #100;
A = 16'h00C4; B = 16'h00D0; #100;
A = 16'h00C4; B = 16'h00D1; #100;
A = 16'h00C4; B = 16'h00D2; #100;
A = 16'h00C4; B = 16'h00D3; #100;
A = 16'h00C4; B = 16'h00D4; #100;
A = 16'h00C4; B = 16'h00D5; #100;
A = 16'h00C4; B = 16'h00D6; #100;
A = 16'h00C4; B = 16'h00D7; #100;
A = 16'h00C4; B = 16'h00D8; #100;
A = 16'h00C4; B = 16'h00D9; #100;
A = 16'h00C4; B = 16'h00DA; #100;
A = 16'h00C4; B = 16'h00DB; #100;
A = 16'h00C4; B = 16'h00DC; #100;
A = 16'h00C4; B = 16'h00DD; #100;
A = 16'h00C4; B = 16'h00DE; #100;
A = 16'h00C4; B = 16'h00DF; #100;
A = 16'h00C4; B = 16'h00E0; #100;
A = 16'h00C4; B = 16'h00E1; #100;
A = 16'h00C4; B = 16'h00E2; #100;
A = 16'h00C4; B = 16'h00E3; #100;
A = 16'h00C4; B = 16'h00E4; #100;
A = 16'h00C4; B = 16'h00E5; #100;
A = 16'h00C4; B = 16'h00E6; #100;
A = 16'h00C4; B = 16'h00E7; #100;
A = 16'h00C4; B = 16'h00E8; #100;
A = 16'h00C4; B = 16'h00E9; #100;
A = 16'h00C4; B = 16'h00EA; #100;
A = 16'h00C4; B = 16'h00EB; #100;
A = 16'h00C4; B = 16'h00EC; #100;
A = 16'h00C4; B = 16'h00ED; #100;
A = 16'h00C4; B = 16'h00EE; #100;
A = 16'h00C4; B = 16'h00EF; #100;
A = 16'h00C4; B = 16'h00F0; #100;
A = 16'h00C4; B = 16'h00F1; #100;
A = 16'h00C4; B = 16'h00F2; #100;
A = 16'h00C4; B = 16'h00F3; #100;
A = 16'h00C4; B = 16'h00F4; #100;
A = 16'h00C4; B = 16'h00F5; #100;
A = 16'h00C4; B = 16'h00F6; #100;
A = 16'h00C4; B = 16'h00F7; #100;
A = 16'h00C4; B = 16'h00F8; #100;
A = 16'h00C4; B = 16'h00F9; #100;
A = 16'h00C4; B = 16'h00FA; #100;
A = 16'h00C4; B = 16'h00FB; #100;
A = 16'h00C4; B = 16'h00FC; #100;
A = 16'h00C4; B = 16'h00FD; #100;
A = 16'h00C4; B = 16'h00FE; #100;
A = 16'h00C4; B = 16'h00FF; #100;
A = 16'h00C5; B = 16'h000; #100;
A = 16'h00C5; B = 16'h001; #100;
A = 16'h00C5; B = 16'h002; #100;
A = 16'h00C5; B = 16'h003; #100;
A = 16'h00C5; B = 16'h004; #100;
A = 16'h00C5; B = 16'h005; #100;
A = 16'h00C5; B = 16'h006; #100;
A = 16'h00C5; B = 16'h007; #100;
A = 16'h00C5; B = 16'h008; #100;
A = 16'h00C5; B = 16'h009; #100;
A = 16'h00C5; B = 16'h00A; #100;
A = 16'h00C5; B = 16'h00B; #100;
A = 16'h00C5; B = 16'h00C; #100;
A = 16'h00C5; B = 16'h00D; #100;
A = 16'h00C5; B = 16'h00E; #100;
A = 16'h00C5; B = 16'h00F; #100;
A = 16'h00C5; B = 16'h0010; #100;
A = 16'h00C5; B = 16'h0011; #100;
A = 16'h00C5; B = 16'h0012; #100;
A = 16'h00C5; B = 16'h0013; #100;
A = 16'h00C5; B = 16'h0014; #100;
A = 16'h00C5; B = 16'h0015; #100;
A = 16'h00C5; B = 16'h0016; #100;
A = 16'h00C5; B = 16'h0017; #100;
A = 16'h00C5; B = 16'h0018; #100;
A = 16'h00C5; B = 16'h0019; #100;
A = 16'h00C5; B = 16'h001A; #100;
A = 16'h00C5; B = 16'h001B; #100;
A = 16'h00C5; B = 16'h001C; #100;
A = 16'h00C5; B = 16'h001D; #100;
A = 16'h00C5; B = 16'h001E; #100;
A = 16'h00C5; B = 16'h001F; #100;
A = 16'h00C5; B = 16'h0020; #100;
A = 16'h00C5; B = 16'h0021; #100;
A = 16'h00C5; B = 16'h0022; #100;
A = 16'h00C5; B = 16'h0023; #100;
A = 16'h00C5; B = 16'h0024; #100;
A = 16'h00C5; B = 16'h0025; #100;
A = 16'h00C5; B = 16'h0026; #100;
A = 16'h00C5; B = 16'h0027; #100;
A = 16'h00C5; B = 16'h0028; #100;
A = 16'h00C5; B = 16'h0029; #100;
A = 16'h00C5; B = 16'h002A; #100;
A = 16'h00C5; B = 16'h002B; #100;
A = 16'h00C5; B = 16'h002C; #100;
A = 16'h00C5; B = 16'h002D; #100;
A = 16'h00C5; B = 16'h002E; #100;
A = 16'h00C5; B = 16'h002F; #100;
A = 16'h00C5; B = 16'h0030; #100;
A = 16'h00C5; B = 16'h0031; #100;
A = 16'h00C5; B = 16'h0032; #100;
A = 16'h00C5; B = 16'h0033; #100;
A = 16'h00C5; B = 16'h0034; #100;
A = 16'h00C5; B = 16'h0035; #100;
A = 16'h00C5; B = 16'h0036; #100;
A = 16'h00C5; B = 16'h0037; #100;
A = 16'h00C5; B = 16'h0038; #100;
A = 16'h00C5; B = 16'h0039; #100;
A = 16'h00C5; B = 16'h003A; #100;
A = 16'h00C5; B = 16'h003B; #100;
A = 16'h00C5; B = 16'h003C; #100;
A = 16'h00C5; B = 16'h003D; #100;
A = 16'h00C5; B = 16'h003E; #100;
A = 16'h00C5; B = 16'h003F; #100;
A = 16'h00C5; B = 16'h0040; #100;
A = 16'h00C5; B = 16'h0041; #100;
A = 16'h00C5; B = 16'h0042; #100;
A = 16'h00C5; B = 16'h0043; #100;
A = 16'h00C5; B = 16'h0044; #100;
A = 16'h00C5; B = 16'h0045; #100;
A = 16'h00C5; B = 16'h0046; #100;
A = 16'h00C5; B = 16'h0047; #100;
A = 16'h00C5; B = 16'h0048; #100;
A = 16'h00C5; B = 16'h0049; #100;
A = 16'h00C5; B = 16'h004A; #100;
A = 16'h00C5; B = 16'h004B; #100;
A = 16'h00C5; B = 16'h004C; #100;
A = 16'h00C5; B = 16'h004D; #100;
A = 16'h00C5; B = 16'h004E; #100;
A = 16'h00C5; B = 16'h004F; #100;
A = 16'h00C5; B = 16'h0050; #100;
A = 16'h00C5; B = 16'h0051; #100;
A = 16'h00C5; B = 16'h0052; #100;
A = 16'h00C5; B = 16'h0053; #100;
A = 16'h00C5; B = 16'h0054; #100;
A = 16'h00C5; B = 16'h0055; #100;
A = 16'h00C5; B = 16'h0056; #100;
A = 16'h00C5; B = 16'h0057; #100;
A = 16'h00C5; B = 16'h0058; #100;
A = 16'h00C5; B = 16'h0059; #100;
A = 16'h00C5; B = 16'h005A; #100;
A = 16'h00C5; B = 16'h005B; #100;
A = 16'h00C5; B = 16'h005C; #100;
A = 16'h00C5; B = 16'h005D; #100;
A = 16'h00C5; B = 16'h005E; #100;
A = 16'h00C5; B = 16'h005F; #100;
A = 16'h00C5; B = 16'h0060; #100;
A = 16'h00C5; B = 16'h0061; #100;
A = 16'h00C5; B = 16'h0062; #100;
A = 16'h00C5; B = 16'h0063; #100;
A = 16'h00C5; B = 16'h0064; #100;
A = 16'h00C5; B = 16'h0065; #100;
A = 16'h00C5; B = 16'h0066; #100;
A = 16'h00C5; B = 16'h0067; #100;
A = 16'h00C5; B = 16'h0068; #100;
A = 16'h00C5; B = 16'h0069; #100;
A = 16'h00C5; B = 16'h006A; #100;
A = 16'h00C5; B = 16'h006B; #100;
A = 16'h00C5; B = 16'h006C; #100;
A = 16'h00C5; B = 16'h006D; #100;
A = 16'h00C5; B = 16'h006E; #100;
A = 16'h00C5; B = 16'h006F; #100;
A = 16'h00C5; B = 16'h0070; #100;
A = 16'h00C5; B = 16'h0071; #100;
A = 16'h00C5; B = 16'h0072; #100;
A = 16'h00C5; B = 16'h0073; #100;
A = 16'h00C5; B = 16'h0074; #100;
A = 16'h00C5; B = 16'h0075; #100;
A = 16'h00C5; B = 16'h0076; #100;
A = 16'h00C5; B = 16'h0077; #100;
A = 16'h00C5; B = 16'h0078; #100;
A = 16'h00C5; B = 16'h0079; #100;
A = 16'h00C5; B = 16'h007A; #100;
A = 16'h00C5; B = 16'h007B; #100;
A = 16'h00C5; B = 16'h007C; #100;
A = 16'h00C5; B = 16'h007D; #100;
A = 16'h00C5; B = 16'h007E; #100;
A = 16'h00C5; B = 16'h007F; #100;
A = 16'h00C5; B = 16'h0080; #100;
A = 16'h00C5; B = 16'h0081; #100;
A = 16'h00C5; B = 16'h0082; #100;
A = 16'h00C5; B = 16'h0083; #100;
A = 16'h00C5; B = 16'h0084; #100;
A = 16'h00C5; B = 16'h0085; #100;
A = 16'h00C5; B = 16'h0086; #100;
A = 16'h00C5; B = 16'h0087; #100;
A = 16'h00C5; B = 16'h0088; #100;
A = 16'h00C5; B = 16'h0089; #100;
A = 16'h00C5; B = 16'h008A; #100;
A = 16'h00C5; B = 16'h008B; #100;
A = 16'h00C5; B = 16'h008C; #100;
A = 16'h00C5; B = 16'h008D; #100;
A = 16'h00C5; B = 16'h008E; #100;
A = 16'h00C5; B = 16'h008F; #100;
A = 16'h00C5; B = 16'h0090; #100;
A = 16'h00C5; B = 16'h0091; #100;
A = 16'h00C5; B = 16'h0092; #100;
A = 16'h00C5; B = 16'h0093; #100;
A = 16'h00C5; B = 16'h0094; #100;
A = 16'h00C5; B = 16'h0095; #100;
A = 16'h00C5; B = 16'h0096; #100;
A = 16'h00C5; B = 16'h0097; #100;
A = 16'h00C5; B = 16'h0098; #100;
A = 16'h00C5; B = 16'h0099; #100;
A = 16'h00C5; B = 16'h009A; #100;
A = 16'h00C5; B = 16'h009B; #100;
A = 16'h00C5; B = 16'h009C; #100;
A = 16'h00C5; B = 16'h009D; #100;
A = 16'h00C5; B = 16'h009E; #100;
A = 16'h00C5; B = 16'h009F; #100;
A = 16'h00C5; B = 16'h00A0; #100;
A = 16'h00C5; B = 16'h00A1; #100;
A = 16'h00C5; B = 16'h00A2; #100;
A = 16'h00C5; B = 16'h00A3; #100;
A = 16'h00C5; B = 16'h00A4; #100;
A = 16'h00C5; B = 16'h00A5; #100;
A = 16'h00C5; B = 16'h00A6; #100;
A = 16'h00C5; B = 16'h00A7; #100;
A = 16'h00C5; B = 16'h00A8; #100;
A = 16'h00C5; B = 16'h00A9; #100;
A = 16'h00C5; B = 16'h00AA; #100;
A = 16'h00C5; B = 16'h00AB; #100;
A = 16'h00C5; B = 16'h00AC; #100;
A = 16'h00C5; B = 16'h00AD; #100;
A = 16'h00C5; B = 16'h00AE; #100;
A = 16'h00C5; B = 16'h00AF; #100;
A = 16'h00C5; B = 16'h00B0; #100;
A = 16'h00C5; B = 16'h00B1; #100;
A = 16'h00C5; B = 16'h00B2; #100;
A = 16'h00C5; B = 16'h00B3; #100;
A = 16'h00C5; B = 16'h00B4; #100;
A = 16'h00C5; B = 16'h00B5; #100;
A = 16'h00C5; B = 16'h00B6; #100;
A = 16'h00C5; B = 16'h00B7; #100;
A = 16'h00C5; B = 16'h00B8; #100;
A = 16'h00C5; B = 16'h00B9; #100;
A = 16'h00C5; B = 16'h00BA; #100;
A = 16'h00C5; B = 16'h00BB; #100;
A = 16'h00C5; B = 16'h00BC; #100;
A = 16'h00C5; B = 16'h00BD; #100;
A = 16'h00C5; B = 16'h00BE; #100;
A = 16'h00C5; B = 16'h00BF; #100;
A = 16'h00C5; B = 16'h00C0; #100;
A = 16'h00C5; B = 16'h00C1; #100;
A = 16'h00C5; B = 16'h00C2; #100;
A = 16'h00C5; B = 16'h00C3; #100;
A = 16'h00C5; B = 16'h00C4; #100;
A = 16'h00C5; B = 16'h00C5; #100;
A = 16'h00C5; B = 16'h00C6; #100;
A = 16'h00C5; B = 16'h00C7; #100;
A = 16'h00C5; B = 16'h00C8; #100;
A = 16'h00C5; B = 16'h00C9; #100;
A = 16'h00C5; B = 16'h00CA; #100;
A = 16'h00C5; B = 16'h00CB; #100;
A = 16'h00C5; B = 16'h00CC; #100;
A = 16'h00C5; B = 16'h00CD; #100;
A = 16'h00C5; B = 16'h00CE; #100;
A = 16'h00C5; B = 16'h00CF; #100;
A = 16'h00C5; B = 16'h00D0; #100;
A = 16'h00C5; B = 16'h00D1; #100;
A = 16'h00C5; B = 16'h00D2; #100;
A = 16'h00C5; B = 16'h00D3; #100;
A = 16'h00C5; B = 16'h00D4; #100;
A = 16'h00C5; B = 16'h00D5; #100;
A = 16'h00C5; B = 16'h00D6; #100;
A = 16'h00C5; B = 16'h00D7; #100;
A = 16'h00C5; B = 16'h00D8; #100;
A = 16'h00C5; B = 16'h00D9; #100;
A = 16'h00C5; B = 16'h00DA; #100;
A = 16'h00C5; B = 16'h00DB; #100;
A = 16'h00C5; B = 16'h00DC; #100;
A = 16'h00C5; B = 16'h00DD; #100;
A = 16'h00C5; B = 16'h00DE; #100;
A = 16'h00C5; B = 16'h00DF; #100;
A = 16'h00C5; B = 16'h00E0; #100;
A = 16'h00C5; B = 16'h00E1; #100;
A = 16'h00C5; B = 16'h00E2; #100;
A = 16'h00C5; B = 16'h00E3; #100;
A = 16'h00C5; B = 16'h00E4; #100;
A = 16'h00C5; B = 16'h00E5; #100;
A = 16'h00C5; B = 16'h00E6; #100;
A = 16'h00C5; B = 16'h00E7; #100;
A = 16'h00C5; B = 16'h00E8; #100;
A = 16'h00C5; B = 16'h00E9; #100;
A = 16'h00C5; B = 16'h00EA; #100;
A = 16'h00C5; B = 16'h00EB; #100;
A = 16'h00C5; B = 16'h00EC; #100;
A = 16'h00C5; B = 16'h00ED; #100;
A = 16'h00C5; B = 16'h00EE; #100;
A = 16'h00C5; B = 16'h00EF; #100;
A = 16'h00C5; B = 16'h00F0; #100;
A = 16'h00C5; B = 16'h00F1; #100;
A = 16'h00C5; B = 16'h00F2; #100;
A = 16'h00C5; B = 16'h00F3; #100;
A = 16'h00C5; B = 16'h00F4; #100;
A = 16'h00C5; B = 16'h00F5; #100;
A = 16'h00C5; B = 16'h00F6; #100;
A = 16'h00C5; B = 16'h00F7; #100;
A = 16'h00C5; B = 16'h00F8; #100;
A = 16'h00C5; B = 16'h00F9; #100;
A = 16'h00C5; B = 16'h00FA; #100;
A = 16'h00C5; B = 16'h00FB; #100;
A = 16'h00C5; B = 16'h00FC; #100;
A = 16'h00C5; B = 16'h00FD; #100;
A = 16'h00C5; B = 16'h00FE; #100;
A = 16'h00C5; B = 16'h00FF; #100;
A = 16'h00C6; B = 16'h000; #100;
A = 16'h00C6; B = 16'h001; #100;
A = 16'h00C6; B = 16'h002; #100;
A = 16'h00C6; B = 16'h003; #100;
A = 16'h00C6; B = 16'h004; #100;
A = 16'h00C6; B = 16'h005; #100;
A = 16'h00C6; B = 16'h006; #100;
A = 16'h00C6; B = 16'h007; #100;
A = 16'h00C6; B = 16'h008; #100;
A = 16'h00C6; B = 16'h009; #100;
A = 16'h00C6; B = 16'h00A; #100;
A = 16'h00C6; B = 16'h00B; #100;
A = 16'h00C6; B = 16'h00C; #100;
A = 16'h00C6; B = 16'h00D; #100;
A = 16'h00C6; B = 16'h00E; #100;
A = 16'h00C6; B = 16'h00F; #100;
A = 16'h00C6; B = 16'h0010; #100;
A = 16'h00C6; B = 16'h0011; #100;
A = 16'h00C6; B = 16'h0012; #100;
A = 16'h00C6; B = 16'h0013; #100;
A = 16'h00C6; B = 16'h0014; #100;
A = 16'h00C6; B = 16'h0015; #100;
A = 16'h00C6; B = 16'h0016; #100;
A = 16'h00C6; B = 16'h0017; #100;
A = 16'h00C6; B = 16'h0018; #100;
A = 16'h00C6; B = 16'h0019; #100;
A = 16'h00C6; B = 16'h001A; #100;
A = 16'h00C6; B = 16'h001B; #100;
A = 16'h00C6; B = 16'h001C; #100;
A = 16'h00C6; B = 16'h001D; #100;
A = 16'h00C6; B = 16'h001E; #100;
A = 16'h00C6; B = 16'h001F; #100;
A = 16'h00C6; B = 16'h0020; #100;
A = 16'h00C6; B = 16'h0021; #100;
A = 16'h00C6; B = 16'h0022; #100;
A = 16'h00C6; B = 16'h0023; #100;
A = 16'h00C6; B = 16'h0024; #100;
A = 16'h00C6; B = 16'h0025; #100;
A = 16'h00C6; B = 16'h0026; #100;
A = 16'h00C6; B = 16'h0027; #100;
A = 16'h00C6; B = 16'h0028; #100;
A = 16'h00C6; B = 16'h0029; #100;
A = 16'h00C6; B = 16'h002A; #100;
A = 16'h00C6; B = 16'h002B; #100;
A = 16'h00C6; B = 16'h002C; #100;
A = 16'h00C6; B = 16'h002D; #100;
A = 16'h00C6; B = 16'h002E; #100;
A = 16'h00C6; B = 16'h002F; #100;
A = 16'h00C6; B = 16'h0030; #100;
A = 16'h00C6; B = 16'h0031; #100;
A = 16'h00C6; B = 16'h0032; #100;
A = 16'h00C6; B = 16'h0033; #100;
A = 16'h00C6; B = 16'h0034; #100;
A = 16'h00C6; B = 16'h0035; #100;
A = 16'h00C6; B = 16'h0036; #100;
A = 16'h00C6; B = 16'h0037; #100;
A = 16'h00C6; B = 16'h0038; #100;
A = 16'h00C6; B = 16'h0039; #100;
A = 16'h00C6; B = 16'h003A; #100;
A = 16'h00C6; B = 16'h003B; #100;
A = 16'h00C6; B = 16'h003C; #100;
A = 16'h00C6; B = 16'h003D; #100;
A = 16'h00C6; B = 16'h003E; #100;
A = 16'h00C6; B = 16'h003F; #100;
A = 16'h00C6; B = 16'h0040; #100;
A = 16'h00C6; B = 16'h0041; #100;
A = 16'h00C6; B = 16'h0042; #100;
A = 16'h00C6; B = 16'h0043; #100;
A = 16'h00C6; B = 16'h0044; #100;
A = 16'h00C6; B = 16'h0045; #100;
A = 16'h00C6; B = 16'h0046; #100;
A = 16'h00C6; B = 16'h0047; #100;
A = 16'h00C6; B = 16'h0048; #100;
A = 16'h00C6; B = 16'h0049; #100;
A = 16'h00C6; B = 16'h004A; #100;
A = 16'h00C6; B = 16'h004B; #100;
A = 16'h00C6; B = 16'h004C; #100;
A = 16'h00C6; B = 16'h004D; #100;
A = 16'h00C6; B = 16'h004E; #100;
A = 16'h00C6; B = 16'h004F; #100;
A = 16'h00C6; B = 16'h0050; #100;
A = 16'h00C6; B = 16'h0051; #100;
A = 16'h00C6; B = 16'h0052; #100;
A = 16'h00C6; B = 16'h0053; #100;
A = 16'h00C6; B = 16'h0054; #100;
A = 16'h00C6; B = 16'h0055; #100;
A = 16'h00C6; B = 16'h0056; #100;
A = 16'h00C6; B = 16'h0057; #100;
A = 16'h00C6; B = 16'h0058; #100;
A = 16'h00C6; B = 16'h0059; #100;
A = 16'h00C6; B = 16'h005A; #100;
A = 16'h00C6; B = 16'h005B; #100;
A = 16'h00C6; B = 16'h005C; #100;
A = 16'h00C6; B = 16'h005D; #100;
A = 16'h00C6; B = 16'h005E; #100;
A = 16'h00C6; B = 16'h005F; #100;
A = 16'h00C6; B = 16'h0060; #100;
A = 16'h00C6; B = 16'h0061; #100;
A = 16'h00C6; B = 16'h0062; #100;
A = 16'h00C6; B = 16'h0063; #100;
A = 16'h00C6; B = 16'h0064; #100;
A = 16'h00C6; B = 16'h0065; #100;
A = 16'h00C6; B = 16'h0066; #100;
A = 16'h00C6; B = 16'h0067; #100;
A = 16'h00C6; B = 16'h0068; #100;
A = 16'h00C6; B = 16'h0069; #100;
A = 16'h00C6; B = 16'h006A; #100;
A = 16'h00C6; B = 16'h006B; #100;
A = 16'h00C6; B = 16'h006C; #100;
A = 16'h00C6; B = 16'h006D; #100;
A = 16'h00C6; B = 16'h006E; #100;
A = 16'h00C6; B = 16'h006F; #100;
A = 16'h00C6; B = 16'h0070; #100;
A = 16'h00C6; B = 16'h0071; #100;
A = 16'h00C6; B = 16'h0072; #100;
A = 16'h00C6; B = 16'h0073; #100;
A = 16'h00C6; B = 16'h0074; #100;
A = 16'h00C6; B = 16'h0075; #100;
A = 16'h00C6; B = 16'h0076; #100;
A = 16'h00C6; B = 16'h0077; #100;
A = 16'h00C6; B = 16'h0078; #100;
A = 16'h00C6; B = 16'h0079; #100;
A = 16'h00C6; B = 16'h007A; #100;
A = 16'h00C6; B = 16'h007B; #100;
A = 16'h00C6; B = 16'h007C; #100;
A = 16'h00C6; B = 16'h007D; #100;
A = 16'h00C6; B = 16'h007E; #100;
A = 16'h00C6; B = 16'h007F; #100;
A = 16'h00C6; B = 16'h0080; #100;
A = 16'h00C6; B = 16'h0081; #100;
A = 16'h00C6; B = 16'h0082; #100;
A = 16'h00C6; B = 16'h0083; #100;
A = 16'h00C6; B = 16'h0084; #100;
A = 16'h00C6; B = 16'h0085; #100;
A = 16'h00C6; B = 16'h0086; #100;
A = 16'h00C6; B = 16'h0087; #100;
A = 16'h00C6; B = 16'h0088; #100;
A = 16'h00C6; B = 16'h0089; #100;
A = 16'h00C6; B = 16'h008A; #100;
A = 16'h00C6; B = 16'h008B; #100;
A = 16'h00C6; B = 16'h008C; #100;
A = 16'h00C6; B = 16'h008D; #100;
A = 16'h00C6; B = 16'h008E; #100;
A = 16'h00C6; B = 16'h008F; #100;
A = 16'h00C6; B = 16'h0090; #100;
A = 16'h00C6; B = 16'h0091; #100;
A = 16'h00C6; B = 16'h0092; #100;
A = 16'h00C6; B = 16'h0093; #100;
A = 16'h00C6; B = 16'h0094; #100;
A = 16'h00C6; B = 16'h0095; #100;
A = 16'h00C6; B = 16'h0096; #100;
A = 16'h00C6; B = 16'h0097; #100;
A = 16'h00C6; B = 16'h0098; #100;
A = 16'h00C6; B = 16'h0099; #100;
A = 16'h00C6; B = 16'h009A; #100;
A = 16'h00C6; B = 16'h009B; #100;
A = 16'h00C6; B = 16'h009C; #100;
A = 16'h00C6; B = 16'h009D; #100;
A = 16'h00C6; B = 16'h009E; #100;
A = 16'h00C6; B = 16'h009F; #100;
A = 16'h00C6; B = 16'h00A0; #100;
A = 16'h00C6; B = 16'h00A1; #100;
A = 16'h00C6; B = 16'h00A2; #100;
A = 16'h00C6; B = 16'h00A3; #100;
A = 16'h00C6; B = 16'h00A4; #100;
A = 16'h00C6; B = 16'h00A5; #100;
A = 16'h00C6; B = 16'h00A6; #100;
A = 16'h00C6; B = 16'h00A7; #100;
A = 16'h00C6; B = 16'h00A8; #100;
A = 16'h00C6; B = 16'h00A9; #100;
A = 16'h00C6; B = 16'h00AA; #100;
A = 16'h00C6; B = 16'h00AB; #100;
A = 16'h00C6; B = 16'h00AC; #100;
A = 16'h00C6; B = 16'h00AD; #100;
A = 16'h00C6; B = 16'h00AE; #100;
A = 16'h00C6; B = 16'h00AF; #100;
A = 16'h00C6; B = 16'h00B0; #100;
A = 16'h00C6; B = 16'h00B1; #100;
A = 16'h00C6; B = 16'h00B2; #100;
A = 16'h00C6; B = 16'h00B3; #100;
A = 16'h00C6; B = 16'h00B4; #100;
A = 16'h00C6; B = 16'h00B5; #100;
A = 16'h00C6; B = 16'h00B6; #100;
A = 16'h00C6; B = 16'h00B7; #100;
A = 16'h00C6; B = 16'h00B8; #100;
A = 16'h00C6; B = 16'h00B9; #100;
A = 16'h00C6; B = 16'h00BA; #100;
A = 16'h00C6; B = 16'h00BB; #100;
A = 16'h00C6; B = 16'h00BC; #100;
A = 16'h00C6; B = 16'h00BD; #100;
A = 16'h00C6; B = 16'h00BE; #100;
A = 16'h00C6; B = 16'h00BF; #100;
A = 16'h00C6; B = 16'h00C0; #100;
A = 16'h00C6; B = 16'h00C1; #100;
A = 16'h00C6; B = 16'h00C2; #100;
A = 16'h00C6; B = 16'h00C3; #100;
A = 16'h00C6; B = 16'h00C4; #100;
A = 16'h00C6; B = 16'h00C5; #100;
A = 16'h00C6; B = 16'h00C6; #100;
A = 16'h00C6; B = 16'h00C7; #100;
A = 16'h00C6; B = 16'h00C8; #100;
A = 16'h00C6; B = 16'h00C9; #100;
A = 16'h00C6; B = 16'h00CA; #100;
A = 16'h00C6; B = 16'h00CB; #100;
A = 16'h00C6; B = 16'h00CC; #100;
A = 16'h00C6; B = 16'h00CD; #100;
A = 16'h00C6; B = 16'h00CE; #100;
A = 16'h00C6; B = 16'h00CF; #100;
A = 16'h00C6; B = 16'h00D0; #100;
A = 16'h00C6; B = 16'h00D1; #100;
A = 16'h00C6; B = 16'h00D2; #100;
A = 16'h00C6; B = 16'h00D3; #100;
A = 16'h00C6; B = 16'h00D4; #100;
A = 16'h00C6; B = 16'h00D5; #100;
A = 16'h00C6; B = 16'h00D6; #100;
A = 16'h00C6; B = 16'h00D7; #100;
A = 16'h00C6; B = 16'h00D8; #100;
A = 16'h00C6; B = 16'h00D9; #100;
A = 16'h00C6; B = 16'h00DA; #100;
A = 16'h00C6; B = 16'h00DB; #100;
A = 16'h00C6; B = 16'h00DC; #100;
A = 16'h00C6; B = 16'h00DD; #100;
A = 16'h00C6; B = 16'h00DE; #100;
A = 16'h00C6; B = 16'h00DF; #100;
A = 16'h00C6; B = 16'h00E0; #100;
A = 16'h00C6; B = 16'h00E1; #100;
A = 16'h00C6; B = 16'h00E2; #100;
A = 16'h00C6; B = 16'h00E3; #100;
A = 16'h00C6; B = 16'h00E4; #100;
A = 16'h00C6; B = 16'h00E5; #100;
A = 16'h00C6; B = 16'h00E6; #100;
A = 16'h00C6; B = 16'h00E7; #100;
A = 16'h00C6; B = 16'h00E8; #100;
A = 16'h00C6; B = 16'h00E9; #100;
A = 16'h00C6; B = 16'h00EA; #100;
A = 16'h00C6; B = 16'h00EB; #100;
A = 16'h00C6; B = 16'h00EC; #100;
A = 16'h00C6; B = 16'h00ED; #100;
A = 16'h00C6; B = 16'h00EE; #100;
A = 16'h00C6; B = 16'h00EF; #100;
A = 16'h00C6; B = 16'h00F0; #100;
A = 16'h00C6; B = 16'h00F1; #100;
A = 16'h00C6; B = 16'h00F2; #100;
A = 16'h00C6; B = 16'h00F3; #100;
A = 16'h00C6; B = 16'h00F4; #100;
A = 16'h00C6; B = 16'h00F5; #100;
A = 16'h00C6; B = 16'h00F6; #100;
A = 16'h00C6; B = 16'h00F7; #100;
A = 16'h00C6; B = 16'h00F8; #100;
A = 16'h00C6; B = 16'h00F9; #100;
A = 16'h00C6; B = 16'h00FA; #100;
A = 16'h00C6; B = 16'h00FB; #100;
A = 16'h00C6; B = 16'h00FC; #100;
A = 16'h00C6; B = 16'h00FD; #100;
A = 16'h00C6; B = 16'h00FE; #100;
A = 16'h00C6; B = 16'h00FF; #100;
A = 16'h00C7; B = 16'h000; #100;
A = 16'h00C7; B = 16'h001; #100;
A = 16'h00C7; B = 16'h002; #100;
A = 16'h00C7; B = 16'h003; #100;
A = 16'h00C7; B = 16'h004; #100;
A = 16'h00C7; B = 16'h005; #100;
A = 16'h00C7; B = 16'h006; #100;
A = 16'h00C7; B = 16'h007; #100;
A = 16'h00C7; B = 16'h008; #100;
A = 16'h00C7; B = 16'h009; #100;
A = 16'h00C7; B = 16'h00A; #100;
A = 16'h00C7; B = 16'h00B; #100;
A = 16'h00C7; B = 16'h00C; #100;
A = 16'h00C7; B = 16'h00D; #100;
A = 16'h00C7; B = 16'h00E; #100;
A = 16'h00C7; B = 16'h00F; #100;
A = 16'h00C7; B = 16'h0010; #100;
A = 16'h00C7; B = 16'h0011; #100;
A = 16'h00C7; B = 16'h0012; #100;
A = 16'h00C7; B = 16'h0013; #100;
A = 16'h00C7; B = 16'h0014; #100;
A = 16'h00C7; B = 16'h0015; #100;
A = 16'h00C7; B = 16'h0016; #100;
A = 16'h00C7; B = 16'h0017; #100;
A = 16'h00C7; B = 16'h0018; #100;
A = 16'h00C7; B = 16'h0019; #100;
A = 16'h00C7; B = 16'h001A; #100;
A = 16'h00C7; B = 16'h001B; #100;
A = 16'h00C7; B = 16'h001C; #100;
A = 16'h00C7; B = 16'h001D; #100;
A = 16'h00C7; B = 16'h001E; #100;
A = 16'h00C7; B = 16'h001F; #100;
A = 16'h00C7; B = 16'h0020; #100;
A = 16'h00C7; B = 16'h0021; #100;
A = 16'h00C7; B = 16'h0022; #100;
A = 16'h00C7; B = 16'h0023; #100;
A = 16'h00C7; B = 16'h0024; #100;
A = 16'h00C7; B = 16'h0025; #100;
A = 16'h00C7; B = 16'h0026; #100;
A = 16'h00C7; B = 16'h0027; #100;
A = 16'h00C7; B = 16'h0028; #100;
A = 16'h00C7; B = 16'h0029; #100;
A = 16'h00C7; B = 16'h002A; #100;
A = 16'h00C7; B = 16'h002B; #100;
A = 16'h00C7; B = 16'h002C; #100;
A = 16'h00C7; B = 16'h002D; #100;
A = 16'h00C7; B = 16'h002E; #100;
A = 16'h00C7; B = 16'h002F; #100;
A = 16'h00C7; B = 16'h0030; #100;
A = 16'h00C7; B = 16'h0031; #100;
A = 16'h00C7; B = 16'h0032; #100;
A = 16'h00C7; B = 16'h0033; #100;
A = 16'h00C7; B = 16'h0034; #100;
A = 16'h00C7; B = 16'h0035; #100;
A = 16'h00C7; B = 16'h0036; #100;
A = 16'h00C7; B = 16'h0037; #100;
A = 16'h00C7; B = 16'h0038; #100;
A = 16'h00C7; B = 16'h0039; #100;
A = 16'h00C7; B = 16'h003A; #100;
A = 16'h00C7; B = 16'h003B; #100;
A = 16'h00C7; B = 16'h003C; #100;
A = 16'h00C7; B = 16'h003D; #100;
A = 16'h00C7; B = 16'h003E; #100;
A = 16'h00C7; B = 16'h003F; #100;
A = 16'h00C7; B = 16'h0040; #100;
A = 16'h00C7; B = 16'h0041; #100;
A = 16'h00C7; B = 16'h0042; #100;
A = 16'h00C7; B = 16'h0043; #100;
A = 16'h00C7; B = 16'h0044; #100;
A = 16'h00C7; B = 16'h0045; #100;
A = 16'h00C7; B = 16'h0046; #100;
A = 16'h00C7; B = 16'h0047; #100;
A = 16'h00C7; B = 16'h0048; #100;
A = 16'h00C7; B = 16'h0049; #100;
A = 16'h00C7; B = 16'h004A; #100;
A = 16'h00C7; B = 16'h004B; #100;
A = 16'h00C7; B = 16'h004C; #100;
A = 16'h00C7; B = 16'h004D; #100;
A = 16'h00C7; B = 16'h004E; #100;
A = 16'h00C7; B = 16'h004F; #100;
A = 16'h00C7; B = 16'h0050; #100;
A = 16'h00C7; B = 16'h0051; #100;
A = 16'h00C7; B = 16'h0052; #100;
A = 16'h00C7; B = 16'h0053; #100;
A = 16'h00C7; B = 16'h0054; #100;
A = 16'h00C7; B = 16'h0055; #100;
A = 16'h00C7; B = 16'h0056; #100;
A = 16'h00C7; B = 16'h0057; #100;
A = 16'h00C7; B = 16'h0058; #100;
A = 16'h00C7; B = 16'h0059; #100;
A = 16'h00C7; B = 16'h005A; #100;
A = 16'h00C7; B = 16'h005B; #100;
A = 16'h00C7; B = 16'h005C; #100;
A = 16'h00C7; B = 16'h005D; #100;
A = 16'h00C7; B = 16'h005E; #100;
A = 16'h00C7; B = 16'h005F; #100;
A = 16'h00C7; B = 16'h0060; #100;
A = 16'h00C7; B = 16'h0061; #100;
A = 16'h00C7; B = 16'h0062; #100;
A = 16'h00C7; B = 16'h0063; #100;
A = 16'h00C7; B = 16'h0064; #100;
A = 16'h00C7; B = 16'h0065; #100;
A = 16'h00C7; B = 16'h0066; #100;
A = 16'h00C7; B = 16'h0067; #100;
A = 16'h00C7; B = 16'h0068; #100;
A = 16'h00C7; B = 16'h0069; #100;
A = 16'h00C7; B = 16'h006A; #100;
A = 16'h00C7; B = 16'h006B; #100;
A = 16'h00C7; B = 16'h006C; #100;
A = 16'h00C7; B = 16'h006D; #100;
A = 16'h00C7; B = 16'h006E; #100;
A = 16'h00C7; B = 16'h006F; #100;
A = 16'h00C7; B = 16'h0070; #100;
A = 16'h00C7; B = 16'h0071; #100;
A = 16'h00C7; B = 16'h0072; #100;
A = 16'h00C7; B = 16'h0073; #100;
A = 16'h00C7; B = 16'h0074; #100;
A = 16'h00C7; B = 16'h0075; #100;
A = 16'h00C7; B = 16'h0076; #100;
A = 16'h00C7; B = 16'h0077; #100;
A = 16'h00C7; B = 16'h0078; #100;
A = 16'h00C7; B = 16'h0079; #100;
A = 16'h00C7; B = 16'h007A; #100;
A = 16'h00C7; B = 16'h007B; #100;
A = 16'h00C7; B = 16'h007C; #100;
A = 16'h00C7; B = 16'h007D; #100;
A = 16'h00C7; B = 16'h007E; #100;
A = 16'h00C7; B = 16'h007F; #100;
A = 16'h00C7; B = 16'h0080; #100;
A = 16'h00C7; B = 16'h0081; #100;
A = 16'h00C7; B = 16'h0082; #100;
A = 16'h00C7; B = 16'h0083; #100;
A = 16'h00C7; B = 16'h0084; #100;
A = 16'h00C7; B = 16'h0085; #100;
A = 16'h00C7; B = 16'h0086; #100;
A = 16'h00C7; B = 16'h0087; #100;
A = 16'h00C7; B = 16'h0088; #100;
A = 16'h00C7; B = 16'h0089; #100;
A = 16'h00C7; B = 16'h008A; #100;
A = 16'h00C7; B = 16'h008B; #100;
A = 16'h00C7; B = 16'h008C; #100;
A = 16'h00C7; B = 16'h008D; #100;
A = 16'h00C7; B = 16'h008E; #100;
A = 16'h00C7; B = 16'h008F; #100;
A = 16'h00C7; B = 16'h0090; #100;
A = 16'h00C7; B = 16'h0091; #100;
A = 16'h00C7; B = 16'h0092; #100;
A = 16'h00C7; B = 16'h0093; #100;
A = 16'h00C7; B = 16'h0094; #100;
A = 16'h00C7; B = 16'h0095; #100;
A = 16'h00C7; B = 16'h0096; #100;
A = 16'h00C7; B = 16'h0097; #100;
A = 16'h00C7; B = 16'h0098; #100;
A = 16'h00C7; B = 16'h0099; #100;
A = 16'h00C7; B = 16'h009A; #100;
A = 16'h00C7; B = 16'h009B; #100;
A = 16'h00C7; B = 16'h009C; #100;
A = 16'h00C7; B = 16'h009D; #100;
A = 16'h00C7; B = 16'h009E; #100;
A = 16'h00C7; B = 16'h009F; #100;
A = 16'h00C7; B = 16'h00A0; #100;
A = 16'h00C7; B = 16'h00A1; #100;
A = 16'h00C7; B = 16'h00A2; #100;
A = 16'h00C7; B = 16'h00A3; #100;
A = 16'h00C7; B = 16'h00A4; #100;
A = 16'h00C7; B = 16'h00A5; #100;
A = 16'h00C7; B = 16'h00A6; #100;
A = 16'h00C7; B = 16'h00A7; #100;
A = 16'h00C7; B = 16'h00A8; #100;
A = 16'h00C7; B = 16'h00A9; #100;
A = 16'h00C7; B = 16'h00AA; #100;
A = 16'h00C7; B = 16'h00AB; #100;
A = 16'h00C7; B = 16'h00AC; #100;
A = 16'h00C7; B = 16'h00AD; #100;
A = 16'h00C7; B = 16'h00AE; #100;
A = 16'h00C7; B = 16'h00AF; #100;
A = 16'h00C7; B = 16'h00B0; #100;
A = 16'h00C7; B = 16'h00B1; #100;
A = 16'h00C7; B = 16'h00B2; #100;
A = 16'h00C7; B = 16'h00B3; #100;
A = 16'h00C7; B = 16'h00B4; #100;
A = 16'h00C7; B = 16'h00B5; #100;
A = 16'h00C7; B = 16'h00B6; #100;
A = 16'h00C7; B = 16'h00B7; #100;
A = 16'h00C7; B = 16'h00B8; #100;
A = 16'h00C7; B = 16'h00B9; #100;
A = 16'h00C7; B = 16'h00BA; #100;
A = 16'h00C7; B = 16'h00BB; #100;
A = 16'h00C7; B = 16'h00BC; #100;
A = 16'h00C7; B = 16'h00BD; #100;
A = 16'h00C7; B = 16'h00BE; #100;
A = 16'h00C7; B = 16'h00BF; #100;
A = 16'h00C7; B = 16'h00C0; #100;
A = 16'h00C7; B = 16'h00C1; #100;
A = 16'h00C7; B = 16'h00C2; #100;
A = 16'h00C7; B = 16'h00C3; #100;
A = 16'h00C7; B = 16'h00C4; #100;
A = 16'h00C7; B = 16'h00C5; #100;
A = 16'h00C7; B = 16'h00C6; #100;
A = 16'h00C7; B = 16'h00C7; #100;
A = 16'h00C7; B = 16'h00C8; #100;
A = 16'h00C7; B = 16'h00C9; #100;
A = 16'h00C7; B = 16'h00CA; #100;
A = 16'h00C7; B = 16'h00CB; #100;
A = 16'h00C7; B = 16'h00CC; #100;
A = 16'h00C7; B = 16'h00CD; #100;
A = 16'h00C7; B = 16'h00CE; #100;
A = 16'h00C7; B = 16'h00CF; #100;
A = 16'h00C7; B = 16'h00D0; #100;
A = 16'h00C7; B = 16'h00D1; #100;
A = 16'h00C7; B = 16'h00D2; #100;
A = 16'h00C7; B = 16'h00D3; #100;
A = 16'h00C7; B = 16'h00D4; #100;
A = 16'h00C7; B = 16'h00D5; #100;
A = 16'h00C7; B = 16'h00D6; #100;
A = 16'h00C7; B = 16'h00D7; #100;
A = 16'h00C7; B = 16'h00D8; #100;
A = 16'h00C7; B = 16'h00D9; #100;
A = 16'h00C7; B = 16'h00DA; #100;
A = 16'h00C7; B = 16'h00DB; #100;
A = 16'h00C7; B = 16'h00DC; #100;
A = 16'h00C7; B = 16'h00DD; #100;
A = 16'h00C7; B = 16'h00DE; #100;
A = 16'h00C7; B = 16'h00DF; #100;
A = 16'h00C7; B = 16'h00E0; #100;
A = 16'h00C7; B = 16'h00E1; #100;
A = 16'h00C7; B = 16'h00E2; #100;
A = 16'h00C7; B = 16'h00E3; #100;
A = 16'h00C7; B = 16'h00E4; #100;
A = 16'h00C7; B = 16'h00E5; #100;
A = 16'h00C7; B = 16'h00E6; #100;
A = 16'h00C7; B = 16'h00E7; #100;
A = 16'h00C7; B = 16'h00E8; #100;
A = 16'h00C7; B = 16'h00E9; #100;
A = 16'h00C7; B = 16'h00EA; #100;
A = 16'h00C7; B = 16'h00EB; #100;
A = 16'h00C7; B = 16'h00EC; #100;
A = 16'h00C7; B = 16'h00ED; #100;
A = 16'h00C7; B = 16'h00EE; #100;
A = 16'h00C7; B = 16'h00EF; #100;
A = 16'h00C7; B = 16'h00F0; #100;
A = 16'h00C7; B = 16'h00F1; #100;
A = 16'h00C7; B = 16'h00F2; #100;
A = 16'h00C7; B = 16'h00F3; #100;
A = 16'h00C7; B = 16'h00F4; #100;
A = 16'h00C7; B = 16'h00F5; #100;
A = 16'h00C7; B = 16'h00F6; #100;
A = 16'h00C7; B = 16'h00F7; #100;
A = 16'h00C7; B = 16'h00F8; #100;
A = 16'h00C7; B = 16'h00F9; #100;
A = 16'h00C7; B = 16'h00FA; #100;
A = 16'h00C7; B = 16'h00FB; #100;
A = 16'h00C7; B = 16'h00FC; #100;
A = 16'h00C7; B = 16'h00FD; #100;
A = 16'h00C7; B = 16'h00FE; #100;
A = 16'h00C7; B = 16'h00FF; #100;
A = 16'h00C8; B = 16'h000; #100;
A = 16'h00C8; B = 16'h001; #100;
A = 16'h00C8; B = 16'h002; #100;
A = 16'h00C8; B = 16'h003; #100;
A = 16'h00C8; B = 16'h004; #100;
A = 16'h00C8; B = 16'h005; #100;
A = 16'h00C8; B = 16'h006; #100;
A = 16'h00C8; B = 16'h007; #100;
A = 16'h00C8; B = 16'h008; #100;
A = 16'h00C8; B = 16'h009; #100;
A = 16'h00C8; B = 16'h00A; #100;
A = 16'h00C8; B = 16'h00B; #100;
A = 16'h00C8; B = 16'h00C; #100;
A = 16'h00C8; B = 16'h00D; #100;
A = 16'h00C8; B = 16'h00E; #100;
A = 16'h00C8; B = 16'h00F; #100;
A = 16'h00C8; B = 16'h0010; #100;
A = 16'h00C8; B = 16'h0011; #100;
A = 16'h00C8; B = 16'h0012; #100;
A = 16'h00C8; B = 16'h0013; #100;
A = 16'h00C8; B = 16'h0014; #100;
A = 16'h00C8; B = 16'h0015; #100;
A = 16'h00C8; B = 16'h0016; #100;
A = 16'h00C8; B = 16'h0017; #100;
A = 16'h00C8; B = 16'h0018; #100;
A = 16'h00C8; B = 16'h0019; #100;
A = 16'h00C8; B = 16'h001A; #100;
A = 16'h00C8; B = 16'h001B; #100;
A = 16'h00C8; B = 16'h001C; #100;
A = 16'h00C8; B = 16'h001D; #100;
A = 16'h00C8; B = 16'h001E; #100;
A = 16'h00C8; B = 16'h001F; #100;
A = 16'h00C8; B = 16'h0020; #100;
A = 16'h00C8; B = 16'h0021; #100;
A = 16'h00C8; B = 16'h0022; #100;
A = 16'h00C8; B = 16'h0023; #100;
A = 16'h00C8; B = 16'h0024; #100;
A = 16'h00C8; B = 16'h0025; #100;
A = 16'h00C8; B = 16'h0026; #100;
A = 16'h00C8; B = 16'h0027; #100;
A = 16'h00C8; B = 16'h0028; #100;
A = 16'h00C8; B = 16'h0029; #100;
A = 16'h00C8; B = 16'h002A; #100;
A = 16'h00C8; B = 16'h002B; #100;
A = 16'h00C8; B = 16'h002C; #100;
A = 16'h00C8; B = 16'h002D; #100;
A = 16'h00C8; B = 16'h002E; #100;
A = 16'h00C8; B = 16'h002F; #100;
A = 16'h00C8; B = 16'h0030; #100;
A = 16'h00C8; B = 16'h0031; #100;
A = 16'h00C8; B = 16'h0032; #100;
A = 16'h00C8; B = 16'h0033; #100;
A = 16'h00C8; B = 16'h0034; #100;
A = 16'h00C8; B = 16'h0035; #100;
A = 16'h00C8; B = 16'h0036; #100;
A = 16'h00C8; B = 16'h0037; #100;
A = 16'h00C8; B = 16'h0038; #100;
A = 16'h00C8; B = 16'h0039; #100;
A = 16'h00C8; B = 16'h003A; #100;
A = 16'h00C8; B = 16'h003B; #100;
A = 16'h00C8; B = 16'h003C; #100;
A = 16'h00C8; B = 16'h003D; #100;
A = 16'h00C8; B = 16'h003E; #100;
A = 16'h00C8; B = 16'h003F; #100;
A = 16'h00C8; B = 16'h0040; #100;
A = 16'h00C8; B = 16'h0041; #100;
A = 16'h00C8; B = 16'h0042; #100;
A = 16'h00C8; B = 16'h0043; #100;
A = 16'h00C8; B = 16'h0044; #100;
A = 16'h00C8; B = 16'h0045; #100;
A = 16'h00C8; B = 16'h0046; #100;
A = 16'h00C8; B = 16'h0047; #100;
A = 16'h00C8; B = 16'h0048; #100;
A = 16'h00C8; B = 16'h0049; #100;
A = 16'h00C8; B = 16'h004A; #100;
A = 16'h00C8; B = 16'h004B; #100;
A = 16'h00C8; B = 16'h004C; #100;
A = 16'h00C8; B = 16'h004D; #100;
A = 16'h00C8; B = 16'h004E; #100;
A = 16'h00C8; B = 16'h004F; #100;
A = 16'h00C8; B = 16'h0050; #100;
A = 16'h00C8; B = 16'h0051; #100;
A = 16'h00C8; B = 16'h0052; #100;
A = 16'h00C8; B = 16'h0053; #100;
A = 16'h00C8; B = 16'h0054; #100;
A = 16'h00C8; B = 16'h0055; #100;
A = 16'h00C8; B = 16'h0056; #100;
A = 16'h00C8; B = 16'h0057; #100;
A = 16'h00C8; B = 16'h0058; #100;
A = 16'h00C8; B = 16'h0059; #100;
A = 16'h00C8; B = 16'h005A; #100;
A = 16'h00C8; B = 16'h005B; #100;
A = 16'h00C8; B = 16'h005C; #100;
A = 16'h00C8; B = 16'h005D; #100;
A = 16'h00C8; B = 16'h005E; #100;
A = 16'h00C8; B = 16'h005F; #100;
A = 16'h00C8; B = 16'h0060; #100;
A = 16'h00C8; B = 16'h0061; #100;
A = 16'h00C8; B = 16'h0062; #100;
A = 16'h00C8; B = 16'h0063; #100;
A = 16'h00C8; B = 16'h0064; #100;
A = 16'h00C8; B = 16'h0065; #100;
A = 16'h00C8; B = 16'h0066; #100;
A = 16'h00C8; B = 16'h0067; #100;
A = 16'h00C8; B = 16'h0068; #100;
A = 16'h00C8; B = 16'h0069; #100;
A = 16'h00C8; B = 16'h006A; #100;
A = 16'h00C8; B = 16'h006B; #100;
A = 16'h00C8; B = 16'h006C; #100;
A = 16'h00C8; B = 16'h006D; #100;
A = 16'h00C8; B = 16'h006E; #100;
A = 16'h00C8; B = 16'h006F; #100;
A = 16'h00C8; B = 16'h0070; #100;
A = 16'h00C8; B = 16'h0071; #100;
A = 16'h00C8; B = 16'h0072; #100;
A = 16'h00C8; B = 16'h0073; #100;
A = 16'h00C8; B = 16'h0074; #100;
A = 16'h00C8; B = 16'h0075; #100;
A = 16'h00C8; B = 16'h0076; #100;
A = 16'h00C8; B = 16'h0077; #100;
A = 16'h00C8; B = 16'h0078; #100;
A = 16'h00C8; B = 16'h0079; #100;
A = 16'h00C8; B = 16'h007A; #100;
A = 16'h00C8; B = 16'h007B; #100;
A = 16'h00C8; B = 16'h007C; #100;
A = 16'h00C8; B = 16'h007D; #100;
A = 16'h00C8; B = 16'h007E; #100;
A = 16'h00C8; B = 16'h007F; #100;
A = 16'h00C8; B = 16'h0080; #100;
A = 16'h00C8; B = 16'h0081; #100;
A = 16'h00C8; B = 16'h0082; #100;
A = 16'h00C8; B = 16'h0083; #100;
A = 16'h00C8; B = 16'h0084; #100;
A = 16'h00C8; B = 16'h0085; #100;
A = 16'h00C8; B = 16'h0086; #100;
A = 16'h00C8; B = 16'h0087; #100;
A = 16'h00C8; B = 16'h0088; #100;
A = 16'h00C8; B = 16'h0089; #100;
A = 16'h00C8; B = 16'h008A; #100;
A = 16'h00C8; B = 16'h008B; #100;
A = 16'h00C8; B = 16'h008C; #100;
A = 16'h00C8; B = 16'h008D; #100;
A = 16'h00C8; B = 16'h008E; #100;
A = 16'h00C8; B = 16'h008F; #100;
A = 16'h00C8; B = 16'h0090; #100;
A = 16'h00C8; B = 16'h0091; #100;
A = 16'h00C8; B = 16'h0092; #100;
A = 16'h00C8; B = 16'h0093; #100;
A = 16'h00C8; B = 16'h0094; #100;
A = 16'h00C8; B = 16'h0095; #100;
A = 16'h00C8; B = 16'h0096; #100;
A = 16'h00C8; B = 16'h0097; #100;
A = 16'h00C8; B = 16'h0098; #100;
A = 16'h00C8; B = 16'h0099; #100;
A = 16'h00C8; B = 16'h009A; #100;
A = 16'h00C8; B = 16'h009B; #100;
A = 16'h00C8; B = 16'h009C; #100;
A = 16'h00C8; B = 16'h009D; #100;
A = 16'h00C8; B = 16'h009E; #100;
A = 16'h00C8; B = 16'h009F; #100;
A = 16'h00C8; B = 16'h00A0; #100;
A = 16'h00C8; B = 16'h00A1; #100;
A = 16'h00C8; B = 16'h00A2; #100;
A = 16'h00C8; B = 16'h00A3; #100;
A = 16'h00C8; B = 16'h00A4; #100;
A = 16'h00C8; B = 16'h00A5; #100;
A = 16'h00C8; B = 16'h00A6; #100;
A = 16'h00C8; B = 16'h00A7; #100;
A = 16'h00C8; B = 16'h00A8; #100;
A = 16'h00C8; B = 16'h00A9; #100;
A = 16'h00C8; B = 16'h00AA; #100;
A = 16'h00C8; B = 16'h00AB; #100;
A = 16'h00C8; B = 16'h00AC; #100;
A = 16'h00C8; B = 16'h00AD; #100;
A = 16'h00C8; B = 16'h00AE; #100;
A = 16'h00C8; B = 16'h00AF; #100;
A = 16'h00C8; B = 16'h00B0; #100;
A = 16'h00C8; B = 16'h00B1; #100;
A = 16'h00C8; B = 16'h00B2; #100;
A = 16'h00C8; B = 16'h00B3; #100;
A = 16'h00C8; B = 16'h00B4; #100;
A = 16'h00C8; B = 16'h00B5; #100;
A = 16'h00C8; B = 16'h00B6; #100;
A = 16'h00C8; B = 16'h00B7; #100;
A = 16'h00C8; B = 16'h00B8; #100;
A = 16'h00C8; B = 16'h00B9; #100;
A = 16'h00C8; B = 16'h00BA; #100;
A = 16'h00C8; B = 16'h00BB; #100;
A = 16'h00C8; B = 16'h00BC; #100;
A = 16'h00C8; B = 16'h00BD; #100;
A = 16'h00C8; B = 16'h00BE; #100;
A = 16'h00C8; B = 16'h00BF; #100;
A = 16'h00C8; B = 16'h00C0; #100;
A = 16'h00C8; B = 16'h00C1; #100;
A = 16'h00C8; B = 16'h00C2; #100;
A = 16'h00C8; B = 16'h00C3; #100;
A = 16'h00C8; B = 16'h00C4; #100;
A = 16'h00C8; B = 16'h00C5; #100;
A = 16'h00C8; B = 16'h00C6; #100;
A = 16'h00C8; B = 16'h00C7; #100;
A = 16'h00C8; B = 16'h00C8; #100;
A = 16'h00C8; B = 16'h00C9; #100;
A = 16'h00C8; B = 16'h00CA; #100;
A = 16'h00C8; B = 16'h00CB; #100;
A = 16'h00C8; B = 16'h00CC; #100;
A = 16'h00C8; B = 16'h00CD; #100;
A = 16'h00C8; B = 16'h00CE; #100;
A = 16'h00C8; B = 16'h00CF; #100;
A = 16'h00C8; B = 16'h00D0; #100;
A = 16'h00C8; B = 16'h00D1; #100;
A = 16'h00C8; B = 16'h00D2; #100;
A = 16'h00C8; B = 16'h00D3; #100;
A = 16'h00C8; B = 16'h00D4; #100;
A = 16'h00C8; B = 16'h00D5; #100;
A = 16'h00C8; B = 16'h00D6; #100;
A = 16'h00C8; B = 16'h00D7; #100;
A = 16'h00C8; B = 16'h00D8; #100;
A = 16'h00C8; B = 16'h00D9; #100;
A = 16'h00C8; B = 16'h00DA; #100;
A = 16'h00C8; B = 16'h00DB; #100;
A = 16'h00C8; B = 16'h00DC; #100;
A = 16'h00C8; B = 16'h00DD; #100;
A = 16'h00C8; B = 16'h00DE; #100;
A = 16'h00C8; B = 16'h00DF; #100;
A = 16'h00C8; B = 16'h00E0; #100;
A = 16'h00C8; B = 16'h00E1; #100;
A = 16'h00C8; B = 16'h00E2; #100;
A = 16'h00C8; B = 16'h00E3; #100;
A = 16'h00C8; B = 16'h00E4; #100;
A = 16'h00C8; B = 16'h00E5; #100;
A = 16'h00C8; B = 16'h00E6; #100;
A = 16'h00C8; B = 16'h00E7; #100;
A = 16'h00C8; B = 16'h00E8; #100;
A = 16'h00C8; B = 16'h00E9; #100;
A = 16'h00C8; B = 16'h00EA; #100;
A = 16'h00C8; B = 16'h00EB; #100;
A = 16'h00C8; B = 16'h00EC; #100;
A = 16'h00C8; B = 16'h00ED; #100;
A = 16'h00C8; B = 16'h00EE; #100;
A = 16'h00C8; B = 16'h00EF; #100;
A = 16'h00C8; B = 16'h00F0; #100;
A = 16'h00C8; B = 16'h00F1; #100;
A = 16'h00C8; B = 16'h00F2; #100;
A = 16'h00C8; B = 16'h00F3; #100;
A = 16'h00C8; B = 16'h00F4; #100;
A = 16'h00C8; B = 16'h00F5; #100;
A = 16'h00C8; B = 16'h00F6; #100;
A = 16'h00C8; B = 16'h00F7; #100;
A = 16'h00C8; B = 16'h00F8; #100;
A = 16'h00C8; B = 16'h00F9; #100;
A = 16'h00C8; B = 16'h00FA; #100;
A = 16'h00C8; B = 16'h00FB; #100;
A = 16'h00C8; B = 16'h00FC; #100;
A = 16'h00C8; B = 16'h00FD; #100;
A = 16'h00C8; B = 16'h00FE; #100;
A = 16'h00C8; B = 16'h00FF; #100;
A = 16'h00C9; B = 16'h000; #100;
A = 16'h00C9; B = 16'h001; #100;
A = 16'h00C9; B = 16'h002; #100;
A = 16'h00C9; B = 16'h003; #100;
A = 16'h00C9; B = 16'h004; #100;
A = 16'h00C9; B = 16'h005; #100;
A = 16'h00C9; B = 16'h006; #100;
A = 16'h00C9; B = 16'h007; #100;
A = 16'h00C9; B = 16'h008; #100;
A = 16'h00C9; B = 16'h009; #100;
A = 16'h00C9; B = 16'h00A; #100;
A = 16'h00C9; B = 16'h00B; #100;
A = 16'h00C9; B = 16'h00C; #100;
A = 16'h00C9; B = 16'h00D; #100;
A = 16'h00C9; B = 16'h00E; #100;
A = 16'h00C9; B = 16'h00F; #100;
A = 16'h00C9; B = 16'h0010; #100;
A = 16'h00C9; B = 16'h0011; #100;
A = 16'h00C9; B = 16'h0012; #100;
A = 16'h00C9; B = 16'h0013; #100;
A = 16'h00C9; B = 16'h0014; #100;
A = 16'h00C9; B = 16'h0015; #100;
A = 16'h00C9; B = 16'h0016; #100;
A = 16'h00C9; B = 16'h0017; #100;
A = 16'h00C9; B = 16'h0018; #100;
A = 16'h00C9; B = 16'h0019; #100;
A = 16'h00C9; B = 16'h001A; #100;
A = 16'h00C9; B = 16'h001B; #100;
A = 16'h00C9; B = 16'h001C; #100;
A = 16'h00C9; B = 16'h001D; #100;
A = 16'h00C9; B = 16'h001E; #100;
A = 16'h00C9; B = 16'h001F; #100;
A = 16'h00C9; B = 16'h0020; #100;
A = 16'h00C9; B = 16'h0021; #100;
A = 16'h00C9; B = 16'h0022; #100;
A = 16'h00C9; B = 16'h0023; #100;
A = 16'h00C9; B = 16'h0024; #100;
A = 16'h00C9; B = 16'h0025; #100;
A = 16'h00C9; B = 16'h0026; #100;
A = 16'h00C9; B = 16'h0027; #100;
A = 16'h00C9; B = 16'h0028; #100;
A = 16'h00C9; B = 16'h0029; #100;
A = 16'h00C9; B = 16'h002A; #100;
A = 16'h00C9; B = 16'h002B; #100;
A = 16'h00C9; B = 16'h002C; #100;
A = 16'h00C9; B = 16'h002D; #100;
A = 16'h00C9; B = 16'h002E; #100;
A = 16'h00C9; B = 16'h002F; #100;
A = 16'h00C9; B = 16'h0030; #100;
A = 16'h00C9; B = 16'h0031; #100;
A = 16'h00C9; B = 16'h0032; #100;
A = 16'h00C9; B = 16'h0033; #100;
A = 16'h00C9; B = 16'h0034; #100;
A = 16'h00C9; B = 16'h0035; #100;
A = 16'h00C9; B = 16'h0036; #100;
A = 16'h00C9; B = 16'h0037; #100;
A = 16'h00C9; B = 16'h0038; #100;
A = 16'h00C9; B = 16'h0039; #100;
A = 16'h00C9; B = 16'h003A; #100;
A = 16'h00C9; B = 16'h003B; #100;
A = 16'h00C9; B = 16'h003C; #100;
A = 16'h00C9; B = 16'h003D; #100;
A = 16'h00C9; B = 16'h003E; #100;
A = 16'h00C9; B = 16'h003F; #100;
A = 16'h00C9; B = 16'h0040; #100;
A = 16'h00C9; B = 16'h0041; #100;
A = 16'h00C9; B = 16'h0042; #100;
A = 16'h00C9; B = 16'h0043; #100;
A = 16'h00C9; B = 16'h0044; #100;
A = 16'h00C9; B = 16'h0045; #100;
A = 16'h00C9; B = 16'h0046; #100;
A = 16'h00C9; B = 16'h0047; #100;
A = 16'h00C9; B = 16'h0048; #100;
A = 16'h00C9; B = 16'h0049; #100;
A = 16'h00C9; B = 16'h004A; #100;
A = 16'h00C9; B = 16'h004B; #100;
A = 16'h00C9; B = 16'h004C; #100;
A = 16'h00C9; B = 16'h004D; #100;
A = 16'h00C9; B = 16'h004E; #100;
A = 16'h00C9; B = 16'h004F; #100;
A = 16'h00C9; B = 16'h0050; #100;
A = 16'h00C9; B = 16'h0051; #100;
A = 16'h00C9; B = 16'h0052; #100;
A = 16'h00C9; B = 16'h0053; #100;
A = 16'h00C9; B = 16'h0054; #100;
A = 16'h00C9; B = 16'h0055; #100;
A = 16'h00C9; B = 16'h0056; #100;
A = 16'h00C9; B = 16'h0057; #100;
A = 16'h00C9; B = 16'h0058; #100;
A = 16'h00C9; B = 16'h0059; #100;
A = 16'h00C9; B = 16'h005A; #100;
A = 16'h00C9; B = 16'h005B; #100;
A = 16'h00C9; B = 16'h005C; #100;
A = 16'h00C9; B = 16'h005D; #100;
A = 16'h00C9; B = 16'h005E; #100;
A = 16'h00C9; B = 16'h005F; #100;
A = 16'h00C9; B = 16'h0060; #100;
A = 16'h00C9; B = 16'h0061; #100;
A = 16'h00C9; B = 16'h0062; #100;
A = 16'h00C9; B = 16'h0063; #100;
A = 16'h00C9; B = 16'h0064; #100;
A = 16'h00C9; B = 16'h0065; #100;
A = 16'h00C9; B = 16'h0066; #100;
A = 16'h00C9; B = 16'h0067; #100;
A = 16'h00C9; B = 16'h0068; #100;
A = 16'h00C9; B = 16'h0069; #100;
A = 16'h00C9; B = 16'h006A; #100;
A = 16'h00C9; B = 16'h006B; #100;
A = 16'h00C9; B = 16'h006C; #100;
A = 16'h00C9; B = 16'h006D; #100;
A = 16'h00C9; B = 16'h006E; #100;
A = 16'h00C9; B = 16'h006F; #100;
A = 16'h00C9; B = 16'h0070; #100;
A = 16'h00C9; B = 16'h0071; #100;
A = 16'h00C9; B = 16'h0072; #100;
A = 16'h00C9; B = 16'h0073; #100;
A = 16'h00C9; B = 16'h0074; #100;
A = 16'h00C9; B = 16'h0075; #100;
A = 16'h00C9; B = 16'h0076; #100;
A = 16'h00C9; B = 16'h0077; #100;
A = 16'h00C9; B = 16'h0078; #100;
A = 16'h00C9; B = 16'h0079; #100;
A = 16'h00C9; B = 16'h007A; #100;
A = 16'h00C9; B = 16'h007B; #100;
A = 16'h00C9; B = 16'h007C; #100;
A = 16'h00C9; B = 16'h007D; #100;
A = 16'h00C9; B = 16'h007E; #100;
A = 16'h00C9; B = 16'h007F; #100;
A = 16'h00C9; B = 16'h0080; #100;
A = 16'h00C9; B = 16'h0081; #100;
A = 16'h00C9; B = 16'h0082; #100;
A = 16'h00C9; B = 16'h0083; #100;
A = 16'h00C9; B = 16'h0084; #100;
A = 16'h00C9; B = 16'h0085; #100;
A = 16'h00C9; B = 16'h0086; #100;
A = 16'h00C9; B = 16'h0087; #100;
A = 16'h00C9; B = 16'h0088; #100;
A = 16'h00C9; B = 16'h0089; #100;
A = 16'h00C9; B = 16'h008A; #100;
A = 16'h00C9; B = 16'h008B; #100;
A = 16'h00C9; B = 16'h008C; #100;
A = 16'h00C9; B = 16'h008D; #100;
A = 16'h00C9; B = 16'h008E; #100;
A = 16'h00C9; B = 16'h008F; #100;
A = 16'h00C9; B = 16'h0090; #100;
A = 16'h00C9; B = 16'h0091; #100;
A = 16'h00C9; B = 16'h0092; #100;
A = 16'h00C9; B = 16'h0093; #100;
A = 16'h00C9; B = 16'h0094; #100;
A = 16'h00C9; B = 16'h0095; #100;
A = 16'h00C9; B = 16'h0096; #100;
A = 16'h00C9; B = 16'h0097; #100;
A = 16'h00C9; B = 16'h0098; #100;
A = 16'h00C9; B = 16'h0099; #100;
A = 16'h00C9; B = 16'h009A; #100;
A = 16'h00C9; B = 16'h009B; #100;
A = 16'h00C9; B = 16'h009C; #100;
A = 16'h00C9; B = 16'h009D; #100;
A = 16'h00C9; B = 16'h009E; #100;
A = 16'h00C9; B = 16'h009F; #100;
A = 16'h00C9; B = 16'h00A0; #100;
A = 16'h00C9; B = 16'h00A1; #100;
A = 16'h00C9; B = 16'h00A2; #100;
A = 16'h00C9; B = 16'h00A3; #100;
A = 16'h00C9; B = 16'h00A4; #100;
A = 16'h00C9; B = 16'h00A5; #100;
A = 16'h00C9; B = 16'h00A6; #100;
A = 16'h00C9; B = 16'h00A7; #100;
A = 16'h00C9; B = 16'h00A8; #100;
A = 16'h00C9; B = 16'h00A9; #100;
A = 16'h00C9; B = 16'h00AA; #100;
A = 16'h00C9; B = 16'h00AB; #100;
A = 16'h00C9; B = 16'h00AC; #100;
A = 16'h00C9; B = 16'h00AD; #100;
A = 16'h00C9; B = 16'h00AE; #100;
A = 16'h00C9; B = 16'h00AF; #100;
A = 16'h00C9; B = 16'h00B0; #100;
A = 16'h00C9; B = 16'h00B1; #100;
A = 16'h00C9; B = 16'h00B2; #100;
A = 16'h00C9; B = 16'h00B3; #100;
A = 16'h00C9; B = 16'h00B4; #100;
A = 16'h00C9; B = 16'h00B5; #100;
A = 16'h00C9; B = 16'h00B6; #100;
A = 16'h00C9; B = 16'h00B7; #100;
A = 16'h00C9; B = 16'h00B8; #100;
A = 16'h00C9; B = 16'h00B9; #100;
A = 16'h00C9; B = 16'h00BA; #100;
A = 16'h00C9; B = 16'h00BB; #100;
A = 16'h00C9; B = 16'h00BC; #100;
A = 16'h00C9; B = 16'h00BD; #100;
A = 16'h00C9; B = 16'h00BE; #100;
A = 16'h00C9; B = 16'h00BF; #100;
A = 16'h00C9; B = 16'h00C0; #100;
A = 16'h00C9; B = 16'h00C1; #100;
A = 16'h00C9; B = 16'h00C2; #100;
A = 16'h00C9; B = 16'h00C3; #100;
A = 16'h00C9; B = 16'h00C4; #100;
A = 16'h00C9; B = 16'h00C5; #100;
A = 16'h00C9; B = 16'h00C6; #100;
A = 16'h00C9; B = 16'h00C7; #100;
A = 16'h00C9; B = 16'h00C8; #100;
A = 16'h00C9; B = 16'h00C9; #100;
A = 16'h00C9; B = 16'h00CA; #100;
A = 16'h00C9; B = 16'h00CB; #100;
A = 16'h00C9; B = 16'h00CC; #100;
A = 16'h00C9; B = 16'h00CD; #100;
A = 16'h00C9; B = 16'h00CE; #100;
A = 16'h00C9; B = 16'h00CF; #100;
A = 16'h00C9; B = 16'h00D0; #100;
A = 16'h00C9; B = 16'h00D1; #100;
A = 16'h00C9; B = 16'h00D2; #100;
A = 16'h00C9; B = 16'h00D3; #100;
A = 16'h00C9; B = 16'h00D4; #100;
A = 16'h00C9; B = 16'h00D5; #100;
A = 16'h00C9; B = 16'h00D6; #100;
A = 16'h00C9; B = 16'h00D7; #100;
A = 16'h00C9; B = 16'h00D8; #100;
A = 16'h00C9; B = 16'h00D9; #100;
A = 16'h00C9; B = 16'h00DA; #100;
A = 16'h00C9; B = 16'h00DB; #100;
A = 16'h00C9; B = 16'h00DC; #100;
A = 16'h00C9; B = 16'h00DD; #100;
A = 16'h00C9; B = 16'h00DE; #100;
A = 16'h00C9; B = 16'h00DF; #100;
A = 16'h00C9; B = 16'h00E0; #100;
A = 16'h00C9; B = 16'h00E1; #100;
A = 16'h00C9; B = 16'h00E2; #100;
A = 16'h00C9; B = 16'h00E3; #100;
A = 16'h00C9; B = 16'h00E4; #100;
A = 16'h00C9; B = 16'h00E5; #100;
A = 16'h00C9; B = 16'h00E6; #100;
A = 16'h00C9; B = 16'h00E7; #100;
A = 16'h00C9; B = 16'h00E8; #100;
A = 16'h00C9; B = 16'h00E9; #100;
A = 16'h00C9; B = 16'h00EA; #100;
A = 16'h00C9; B = 16'h00EB; #100;
A = 16'h00C9; B = 16'h00EC; #100;
A = 16'h00C9; B = 16'h00ED; #100;
A = 16'h00C9; B = 16'h00EE; #100;
A = 16'h00C9; B = 16'h00EF; #100;
A = 16'h00C9; B = 16'h00F0; #100;
A = 16'h00C9; B = 16'h00F1; #100;
A = 16'h00C9; B = 16'h00F2; #100;
A = 16'h00C9; B = 16'h00F3; #100;
A = 16'h00C9; B = 16'h00F4; #100;
A = 16'h00C9; B = 16'h00F5; #100;
A = 16'h00C9; B = 16'h00F6; #100;
A = 16'h00C9; B = 16'h00F7; #100;
A = 16'h00C9; B = 16'h00F8; #100;
A = 16'h00C9; B = 16'h00F9; #100;
A = 16'h00C9; B = 16'h00FA; #100;
A = 16'h00C9; B = 16'h00FB; #100;
A = 16'h00C9; B = 16'h00FC; #100;
A = 16'h00C9; B = 16'h00FD; #100;
A = 16'h00C9; B = 16'h00FE; #100;
A = 16'h00C9; B = 16'h00FF; #100;
A = 16'h00CA; B = 16'h000; #100;
A = 16'h00CA; B = 16'h001; #100;
A = 16'h00CA; B = 16'h002; #100;
A = 16'h00CA; B = 16'h003; #100;
A = 16'h00CA; B = 16'h004; #100;
A = 16'h00CA; B = 16'h005; #100;
A = 16'h00CA; B = 16'h006; #100;
A = 16'h00CA; B = 16'h007; #100;
A = 16'h00CA; B = 16'h008; #100;
A = 16'h00CA; B = 16'h009; #100;
A = 16'h00CA; B = 16'h00A; #100;
A = 16'h00CA; B = 16'h00B; #100;
A = 16'h00CA; B = 16'h00C; #100;
A = 16'h00CA; B = 16'h00D; #100;
A = 16'h00CA; B = 16'h00E; #100;
A = 16'h00CA; B = 16'h00F; #100;
A = 16'h00CA; B = 16'h0010; #100;
A = 16'h00CA; B = 16'h0011; #100;
A = 16'h00CA; B = 16'h0012; #100;
A = 16'h00CA; B = 16'h0013; #100;
A = 16'h00CA; B = 16'h0014; #100;
A = 16'h00CA; B = 16'h0015; #100;
A = 16'h00CA; B = 16'h0016; #100;
A = 16'h00CA; B = 16'h0017; #100;
A = 16'h00CA; B = 16'h0018; #100;
A = 16'h00CA; B = 16'h0019; #100;
A = 16'h00CA; B = 16'h001A; #100;
A = 16'h00CA; B = 16'h001B; #100;
A = 16'h00CA; B = 16'h001C; #100;
A = 16'h00CA; B = 16'h001D; #100;
A = 16'h00CA; B = 16'h001E; #100;
A = 16'h00CA; B = 16'h001F; #100;
A = 16'h00CA; B = 16'h0020; #100;
A = 16'h00CA; B = 16'h0021; #100;
A = 16'h00CA; B = 16'h0022; #100;
A = 16'h00CA; B = 16'h0023; #100;
A = 16'h00CA; B = 16'h0024; #100;
A = 16'h00CA; B = 16'h0025; #100;
A = 16'h00CA; B = 16'h0026; #100;
A = 16'h00CA; B = 16'h0027; #100;
A = 16'h00CA; B = 16'h0028; #100;
A = 16'h00CA; B = 16'h0029; #100;
A = 16'h00CA; B = 16'h002A; #100;
A = 16'h00CA; B = 16'h002B; #100;
A = 16'h00CA; B = 16'h002C; #100;
A = 16'h00CA; B = 16'h002D; #100;
A = 16'h00CA; B = 16'h002E; #100;
A = 16'h00CA; B = 16'h002F; #100;
A = 16'h00CA; B = 16'h0030; #100;
A = 16'h00CA; B = 16'h0031; #100;
A = 16'h00CA; B = 16'h0032; #100;
A = 16'h00CA; B = 16'h0033; #100;
A = 16'h00CA; B = 16'h0034; #100;
A = 16'h00CA; B = 16'h0035; #100;
A = 16'h00CA; B = 16'h0036; #100;
A = 16'h00CA; B = 16'h0037; #100;
A = 16'h00CA; B = 16'h0038; #100;
A = 16'h00CA; B = 16'h0039; #100;
A = 16'h00CA; B = 16'h003A; #100;
A = 16'h00CA; B = 16'h003B; #100;
A = 16'h00CA; B = 16'h003C; #100;
A = 16'h00CA; B = 16'h003D; #100;
A = 16'h00CA; B = 16'h003E; #100;
A = 16'h00CA; B = 16'h003F; #100;
A = 16'h00CA; B = 16'h0040; #100;
A = 16'h00CA; B = 16'h0041; #100;
A = 16'h00CA; B = 16'h0042; #100;
A = 16'h00CA; B = 16'h0043; #100;
A = 16'h00CA; B = 16'h0044; #100;
A = 16'h00CA; B = 16'h0045; #100;
A = 16'h00CA; B = 16'h0046; #100;
A = 16'h00CA; B = 16'h0047; #100;
A = 16'h00CA; B = 16'h0048; #100;
A = 16'h00CA; B = 16'h0049; #100;
A = 16'h00CA; B = 16'h004A; #100;
A = 16'h00CA; B = 16'h004B; #100;
A = 16'h00CA; B = 16'h004C; #100;
A = 16'h00CA; B = 16'h004D; #100;
A = 16'h00CA; B = 16'h004E; #100;
A = 16'h00CA; B = 16'h004F; #100;
A = 16'h00CA; B = 16'h0050; #100;
A = 16'h00CA; B = 16'h0051; #100;
A = 16'h00CA; B = 16'h0052; #100;
A = 16'h00CA; B = 16'h0053; #100;
A = 16'h00CA; B = 16'h0054; #100;
A = 16'h00CA; B = 16'h0055; #100;
A = 16'h00CA; B = 16'h0056; #100;
A = 16'h00CA; B = 16'h0057; #100;
A = 16'h00CA; B = 16'h0058; #100;
A = 16'h00CA; B = 16'h0059; #100;
A = 16'h00CA; B = 16'h005A; #100;
A = 16'h00CA; B = 16'h005B; #100;
A = 16'h00CA; B = 16'h005C; #100;
A = 16'h00CA; B = 16'h005D; #100;
A = 16'h00CA; B = 16'h005E; #100;
A = 16'h00CA; B = 16'h005F; #100;
A = 16'h00CA; B = 16'h0060; #100;
A = 16'h00CA; B = 16'h0061; #100;
A = 16'h00CA; B = 16'h0062; #100;
A = 16'h00CA; B = 16'h0063; #100;
A = 16'h00CA; B = 16'h0064; #100;
A = 16'h00CA; B = 16'h0065; #100;
A = 16'h00CA; B = 16'h0066; #100;
A = 16'h00CA; B = 16'h0067; #100;
A = 16'h00CA; B = 16'h0068; #100;
A = 16'h00CA; B = 16'h0069; #100;
A = 16'h00CA; B = 16'h006A; #100;
A = 16'h00CA; B = 16'h006B; #100;
A = 16'h00CA; B = 16'h006C; #100;
A = 16'h00CA; B = 16'h006D; #100;
A = 16'h00CA; B = 16'h006E; #100;
A = 16'h00CA; B = 16'h006F; #100;
A = 16'h00CA; B = 16'h0070; #100;
A = 16'h00CA; B = 16'h0071; #100;
A = 16'h00CA; B = 16'h0072; #100;
A = 16'h00CA; B = 16'h0073; #100;
A = 16'h00CA; B = 16'h0074; #100;
A = 16'h00CA; B = 16'h0075; #100;
A = 16'h00CA; B = 16'h0076; #100;
A = 16'h00CA; B = 16'h0077; #100;
A = 16'h00CA; B = 16'h0078; #100;
A = 16'h00CA; B = 16'h0079; #100;
A = 16'h00CA; B = 16'h007A; #100;
A = 16'h00CA; B = 16'h007B; #100;
A = 16'h00CA; B = 16'h007C; #100;
A = 16'h00CA; B = 16'h007D; #100;
A = 16'h00CA; B = 16'h007E; #100;
A = 16'h00CA; B = 16'h007F; #100;
A = 16'h00CA; B = 16'h0080; #100;
A = 16'h00CA; B = 16'h0081; #100;
A = 16'h00CA; B = 16'h0082; #100;
A = 16'h00CA; B = 16'h0083; #100;
A = 16'h00CA; B = 16'h0084; #100;
A = 16'h00CA; B = 16'h0085; #100;
A = 16'h00CA; B = 16'h0086; #100;
A = 16'h00CA; B = 16'h0087; #100;
A = 16'h00CA; B = 16'h0088; #100;
A = 16'h00CA; B = 16'h0089; #100;
A = 16'h00CA; B = 16'h008A; #100;
A = 16'h00CA; B = 16'h008B; #100;
A = 16'h00CA; B = 16'h008C; #100;
A = 16'h00CA; B = 16'h008D; #100;
A = 16'h00CA; B = 16'h008E; #100;
A = 16'h00CA; B = 16'h008F; #100;
A = 16'h00CA; B = 16'h0090; #100;
A = 16'h00CA; B = 16'h0091; #100;
A = 16'h00CA; B = 16'h0092; #100;
A = 16'h00CA; B = 16'h0093; #100;
A = 16'h00CA; B = 16'h0094; #100;
A = 16'h00CA; B = 16'h0095; #100;
A = 16'h00CA; B = 16'h0096; #100;
A = 16'h00CA; B = 16'h0097; #100;
A = 16'h00CA; B = 16'h0098; #100;
A = 16'h00CA; B = 16'h0099; #100;
A = 16'h00CA; B = 16'h009A; #100;
A = 16'h00CA; B = 16'h009B; #100;
A = 16'h00CA; B = 16'h009C; #100;
A = 16'h00CA; B = 16'h009D; #100;
A = 16'h00CA; B = 16'h009E; #100;
A = 16'h00CA; B = 16'h009F; #100;
A = 16'h00CA; B = 16'h00A0; #100;
A = 16'h00CA; B = 16'h00A1; #100;
A = 16'h00CA; B = 16'h00A2; #100;
A = 16'h00CA; B = 16'h00A3; #100;
A = 16'h00CA; B = 16'h00A4; #100;
A = 16'h00CA; B = 16'h00A5; #100;
A = 16'h00CA; B = 16'h00A6; #100;
A = 16'h00CA; B = 16'h00A7; #100;
A = 16'h00CA; B = 16'h00A8; #100;
A = 16'h00CA; B = 16'h00A9; #100;
A = 16'h00CA; B = 16'h00AA; #100;
A = 16'h00CA; B = 16'h00AB; #100;
A = 16'h00CA; B = 16'h00AC; #100;
A = 16'h00CA; B = 16'h00AD; #100;
A = 16'h00CA; B = 16'h00AE; #100;
A = 16'h00CA; B = 16'h00AF; #100;
A = 16'h00CA; B = 16'h00B0; #100;
A = 16'h00CA; B = 16'h00B1; #100;
A = 16'h00CA; B = 16'h00B2; #100;
A = 16'h00CA; B = 16'h00B3; #100;
A = 16'h00CA; B = 16'h00B4; #100;
A = 16'h00CA; B = 16'h00B5; #100;
A = 16'h00CA; B = 16'h00B6; #100;
A = 16'h00CA; B = 16'h00B7; #100;
A = 16'h00CA; B = 16'h00B8; #100;
A = 16'h00CA; B = 16'h00B9; #100;
A = 16'h00CA; B = 16'h00BA; #100;
A = 16'h00CA; B = 16'h00BB; #100;
A = 16'h00CA; B = 16'h00BC; #100;
A = 16'h00CA; B = 16'h00BD; #100;
A = 16'h00CA; B = 16'h00BE; #100;
A = 16'h00CA; B = 16'h00BF; #100;
A = 16'h00CA; B = 16'h00C0; #100;
A = 16'h00CA; B = 16'h00C1; #100;
A = 16'h00CA; B = 16'h00C2; #100;
A = 16'h00CA; B = 16'h00C3; #100;
A = 16'h00CA; B = 16'h00C4; #100;
A = 16'h00CA; B = 16'h00C5; #100;
A = 16'h00CA; B = 16'h00C6; #100;
A = 16'h00CA; B = 16'h00C7; #100;
A = 16'h00CA; B = 16'h00C8; #100;
A = 16'h00CA; B = 16'h00C9; #100;
A = 16'h00CA; B = 16'h00CA; #100;
A = 16'h00CA; B = 16'h00CB; #100;
A = 16'h00CA; B = 16'h00CC; #100;
A = 16'h00CA; B = 16'h00CD; #100;
A = 16'h00CA; B = 16'h00CE; #100;
A = 16'h00CA; B = 16'h00CF; #100;
A = 16'h00CA; B = 16'h00D0; #100;
A = 16'h00CA; B = 16'h00D1; #100;
A = 16'h00CA; B = 16'h00D2; #100;
A = 16'h00CA; B = 16'h00D3; #100;
A = 16'h00CA; B = 16'h00D4; #100;
A = 16'h00CA; B = 16'h00D5; #100;
A = 16'h00CA; B = 16'h00D6; #100;
A = 16'h00CA; B = 16'h00D7; #100;
A = 16'h00CA; B = 16'h00D8; #100;
A = 16'h00CA; B = 16'h00D9; #100;
A = 16'h00CA; B = 16'h00DA; #100;
A = 16'h00CA; B = 16'h00DB; #100;
A = 16'h00CA; B = 16'h00DC; #100;
A = 16'h00CA; B = 16'h00DD; #100;
A = 16'h00CA; B = 16'h00DE; #100;
A = 16'h00CA; B = 16'h00DF; #100;
A = 16'h00CA; B = 16'h00E0; #100;
A = 16'h00CA; B = 16'h00E1; #100;
A = 16'h00CA; B = 16'h00E2; #100;
A = 16'h00CA; B = 16'h00E3; #100;
A = 16'h00CA; B = 16'h00E4; #100;
A = 16'h00CA; B = 16'h00E5; #100;
A = 16'h00CA; B = 16'h00E6; #100;
A = 16'h00CA; B = 16'h00E7; #100;
A = 16'h00CA; B = 16'h00E8; #100;
A = 16'h00CA; B = 16'h00E9; #100;
A = 16'h00CA; B = 16'h00EA; #100;
A = 16'h00CA; B = 16'h00EB; #100;
A = 16'h00CA; B = 16'h00EC; #100;
A = 16'h00CA; B = 16'h00ED; #100;
A = 16'h00CA; B = 16'h00EE; #100;
A = 16'h00CA; B = 16'h00EF; #100;
A = 16'h00CA; B = 16'h00F0; #100;
A = 16'h00CA; B = 16'h00F1; #100;
A = 16'h00CA; B = 16'h00F2; #100;
A = 16'h00CA; B = 16'h00F3; #100;
A = 16'h00CA; B = 16'h00F4; #100;
A = 16'h00CA; B = 16'h00F5; #100;
A = 16'h00CA; B = 16'h00F6; #100;
A = 16'h00CA; B = 16'h00F7; #100;
A = 16'h00CA; B = 16'h00F8; #100;
A = 16'h00CA; B = 16'h00F9; #100;
A = 16'h00CA; B = 16'h00FA; #100;
A = 16'h00CA; B = 16'h00FB; #100;
A = 16'h00CA; B = 16'h00FC; #100;
A = 16'h00CA; B = 16'h00FD; #100;
A = 16'h00CA; B = 16'h00FE; #100;
A = 16'h00CA; B = 16'h00FF; #100;
A = 16'h00CB; B = 16'h000; #100;
A = 16'h00CB; B = 16'h001; #100;
A = 16'h00CB; B = 16'h002; #100;
A = 16'h00CB; B = 16'h003; #100;
A = 16'h00CB; B = 16'h004; #100;
A = 16'h00CB; B = 16'h005; #100;
A = 16'h00CB; B = 16'h006; #100;
A = 16'h00CB; B = 16'h007; #100;
A = 16'h00CB; B = 16'h008; #100;
A = 16'h00CB; B = 16'h009; #100;
A = 16'h00CB; B = 16'h00A; #100;
A = 16'h00CB; B = 16'h00B; #100;
A = 16'h00CB; B = 16'h00C; #100;
A = 16'h00CB; B = 16'h00D; #100;
A = 16'h00CB; B = 16'h00E; #100;
A = 16'h00CB; B = 16'h00F; #100;
A = 16'h00CB; B = 16'h0010; #100;
A = 16'h00CB; B = 16'h0011; #100;
A = 16'h00CB; B = 16'h0012; #100;
A = 16'h00CB; B = 16'h0013; #100;
A = 16'h00CB; B = 16'h0014; #100;
A = 16'h00CB; B = 16'h0015; #100;
A = 16'h00CB; B = 16'h0016; #100;
A = 16'h00CB; B = 16'h0017; #100;
A = 16'h00CB; B = 16'h0018; #100;
A = 16'h00CB; B = 16'h0019; #100;
A = 16'h00CB; B = 16'h001A; #100;
A = 16'h00CB; B = 16'h001B; #100;
A = 16'h00CB; B = 16'h001C; #100;
A = 16'h00CB; B = 16'h001D; #100;
A = 16'h00CB; B = 16'h001E; #100;
A = 16'h00CB; B = 16'h001F; #100;
A = 16'h00CB; B = 16'h0020; #100;
A = 16'h00CB; B = 16'h0021; #100;
A = 16'h00CB; B = 16'h0022; #100;
A = 16'h00CB; B = 16'h0023; #100;
A = 16'h00CB; B = 16'h0024; #100;
A = 16'h00CB; B = 16'h0025; #100;
A = 16'h00CB; B = 16'h0026; #100;
A = 16'h00CB; B = 16'h0027; #100;
A = 16'h00CB; B = 16'h0028; #100;
A = 16'h00CB; B = 16'h0029; #100;
A = 16'h00CB; B = 16'h002A; #100;
A = 16'h00CB; B = 16'h002B; #100;
A = 16'h00CB; B = 16'h002C; #100;
A = 16'h00CB; B = 16'h002D; #100;
A = 16'h00CB; B = 16'h002E; #100;
A = 16'h00CB; B = 16'h002F; #100;
A = 16'h00CB; B = 16'h0030; #100;
A = 16'h00CB; B = 16'h0031; #100;
A = 16'h00CB; B = 16'h0032; #100;
A = 16'h00CB; B = 16'h0033; #100;
A = 16'h00CB; B = 16'h0034; #100;
A = 16'h00CB; B = 16'h0035; #100;
A = 16'h00CB; B = 16'h0036; #100;
A = 16'h00CB; B = 16'h0037; #100;
A = 16'h00CB; B = 16'h0038; #100;
A = 16'h00CB; B = 16'h0039; #100;
A = 16'h00CB; B = 16'h003A; #100;
A = 16'h00CB; B = 16'h003B; #100;
A = 16'h00CB; B = 16'h003C; #100;
A = 16'h00CB; B = 16'h003D; #100;
A = 16'h00CB; B = 16'h003E; #100;
A = 16'h00CB; B = 16'h003F; #100;
A = 16'h00CB; B = 16'h0040; #100;
A = 16'h00CB; B = 16'h0041; #100;
A = 16'h00CB; B = 16'h0042; #100;
A = 16'h00CB; B = 16'h0043; #100;
A = 16'h00CB; B = 16'h0044; #100;
A = 16'h00CB; B = 16'h0045; #100;
A = 16'h00CB; B = 16'h0046; #100;
A = 16'h00CB; B = 16'h0047; #100;
A = 16'h00CB; B = 16'h0048; #100;
A = 16'h00CB; B = 16'h0049; #100;
A = 16'h00CB; B = 16'h004A; #100;
A = 16'h00CB; B = 16'h004B; #100;
A = 16'h00CB; B = 16'h004C; #100;
A = 16'h00CB; B = 16'h004D; #100;
A = 16'h00CB; B = 16'h004E; #100;
A = 16'h00CB; B = 16'h004F; #100;
A = 16'h00CB; B = 16'h0050; #100;
A = 16'h00CB; B = 16'h0051; #100;
A = 16'h00CB; B = 16'h0052; #100;
A = 16'h00CB; B = 16'h0053; #100;
A = 16'h00CB; B = 16'h0054; #100;
A = 16'h00CB; B = 16'h0055; #100;
A = 16'h00CB; B = 16'h0056; #100;
A = 16'h00CB; B = 16'h0057; #100;
A = 16'h00CB; B = 16'h0058; #100;
A = 16'h00CB; B = 16'h0059; #100;
A = 16'h00CB; B = 16'h005A; #100;
A = 16'h00CB; B = 16'h005B; #100;
A = 16'h00CB; B = 16'h005C; #100;
A = 16'h00CB; B = 16'h005D; #100;
A = 16'h00CB; B = 16'h005E; #100;
A = 16'h00CB; B = 16'h005F; #100;
A = 16'h00CB; B = 16'h0060; #100;
A = 16'h00CB; B = 16'h0061; #100;
A = 16'h00CB; B = 16'h0062; #100;
A = 16'h00CB; B = 16'h0063; #100;
A = 16'h00CB; B = 16'h0064; #100;
A = 16'h00CB; B = 16'h0065; #100;
A = 16'h00CB; B = 16'h0066; #100;
A = 16'h00CB; B = 16'h0067; #100;
A = 16'h00CB; B = 16'h0068; #100;
A = 16'h00CB; B = 16'h0069; #100;
A = 16'h00CB; B = 16'h006A; #100;
A = 16'h00CB; B = 16'h006B; #100;
A = 16'h00CB; B = 16'h006C; #100;
A = 16'h00CB; B = 16'h006D; #100;
A = 16'h00CB; B = 16'h006E; #100;
A = 16'h00CB; B = 16'h006F; #100;
A = 16'h00CB; B = 16'h0070; #100;
A = 16'h00CB; B = 16'h0071; #100;
A = 16'h00CB; B = 16'h0072; #100;
A = 16'h00CB; B = 16'h0073; #100;
A = 16'h00CB; B = 16'h0074; #100;
A = 16'h00CB; B = 16'h0075; #100;
A = 16'h00CB; B = 16'h0076; #100;
A = 16'h00CB; B = 16'h0077; #100;
A = 16'h00CB; B = 16'h0078; #100;
A = 16'h00CB; B = 16'h0079; #100;
A = 16'h00CB; B = 16'h007A; #100;
A = 16'h00CB; B = 16'h007B; #100;
A = 16'h00CB; B = 16'h007C; #100;
A = 16'h00CB; B = 16'h007D; #100;
A = 16'h00CB; B = 16'h007E; #100;
A = 16'h00CB; B = 16'h007F; #100;
A = 16'h00CB; B = 16'h0080; #100;
A = 16'h00CB; B = 16'h0081; #100;
A = 16'h00CB; B = 16'h0082; #100;
A = 16'h00CB; B = 16'h0083; #100;
A = 16'h00CB; B = 16'h0084; #100;
A = 16'h00CB; B = 16'h0085; #100;
A = 16'h00CB; B = 16'h0086; #100;
A = 16'h00CB; B = 16'h0087; #100;
A = 16'h00CB; B = 16'h0088; #100;
A = 16'h00CB; B = 16'h0089; #100;
A = 16'h00CB; B = 16'h008A; #100;
A = 16'h00CB; B = 16'h008B; #100;
A = 16'h00CB; B = 16'h008C; #100;
A = 16'h00CB; B = 16'h008D; #100;
A = 16'h00CB; B = 16'h008E; #100;
A = 16'h00CB; B = 16'h008F; #100;
A = 16'h00CB; B = 16'h0090; #100;
A = 16'h00CB; B = 16'h0091; #100;
A = 16'h00CB; B = 16'h0092; #100;
A = 16'h00CB; B = 16'h0093; #100;
A = 16'h00CB; B = 16'h0094; #100;
A = 16'h00CB; B = 16'h0095; #100;
A = 16'h00CB; B = 16'h0096; #100;
A = 16'h00CB; B = 16'h0097; #100;
A = 16'h00CB; B = 16'h0098; #100;
A = 16'h00CB; B = 16'h0099; #100;
A = 16'h00CB; B = 16'h009A; #100;
A = 16'h00CB; B = 16'h009B; #100;
A = 16'h00CB; B = 16'h009C; #100;
A = 16'h00CB; B = 16'h009D; #100;
A = 16'h00CB; B = 16'h009E; #100;
A = 16'h00CB; B = 16'h009F; #100;
A = 16'h00CB; B = 16'h00A0; #100;
A = 16'h00CB; B = 16'h00A1; #100;
A = 16'h00CB; B = 16'h00A2; #100;
A = 16'h00CB; B = 16'h00A3; #100;
A = 16'h00CB; B = 16'h00A4; #100;
A = 16'h00CB; B = 16'h00A5; #100;
A = 16'h00CB; B = 16'h00A6; #100;
A = 16'h00CB; B = 16'h00A7; #100;
A = 16'h00CB; B = 16'h00A8; #100;
A = 16'h00CB; B = 16'h00A9; #100;
A = 16'h00CB; B = 16'h00AA; #100;
A = 16'h00CB; B = 16'h00AB; #100;
A = 16'h00CB; B = 16'h00AC; #100;
A = 16'h00CB; B = 16'h00AD; #100;
A = 16'h00CB; B = 16'h00AE; #100;
A = 16'h00CB; B = 16'h00AF; #100;
A = 16'h00CB; B = 16'h00B0; #100;
A = 16'h00CB; B = 16'h00B1; #100;
A = 16'h00CB; B = 16'h00B2; #100;
A = 16'h00CB; B = 16'h00B3; #100;
A = 16'h00CB; B = 16'h00B4; #100;
A = 16'h00CB; B = 16'h00B5; #100;
A = 16'h00CB; B = 16'h00B6; #100;
A = 16'h00CB; B = 16'h00B7; #100;
A = 16'h00CB; B = 16'h00B8; #100;
A = 16'h00CB; B = 16'h00B9; #100;
A = 16'h00CB; B = 16'h00BA; #100;
A = 16'h00CB; B = 16'h00BB; #100;
A = 16'h00CB; B = 16'h00BC; #100;
A = 16'h00CB; B = 16'h00BD; #100;
A = 16'h00CB; B = 16'h00BE; #100;
A = 16'h00CB; B = 16'h00BF; #100;
A = 16'h00CB; B = 16'h00C0; #100;
A = 16'h00CB; B = 16'h00C1; #100;
A = 16'h00CB; B = 16'h00C2; #100;
A = 16'h00CB; B = 16'h00C3; #100;
A = 16'h00CB; B = 16'h00C4; #100;
A = 16'h00CB; B = 16'h00C5; #100;
A = 16'h00CB; B = 16'h00C6; #100;
A = 16'h00CB; B = 16'h00C7; #100;
A = 16'h00CB; B = 16'h00C8; #100;
A = 16'h00CB; B = 16'h00C9; #100;
A = 16'h00CB; B = 16'h00CA; #100;
A = 16'h00CB; B = 16'h00CB; #100;
A = 16'h00CB; B = 16'h00CC; #100;
A = 16'h00CB; B = 16'h00CD; #100;
A = 16'h00CB; B = 16'h00CE; #100;
A = 16'h00CB; B = 16'h00CF; #100;
A = 16'h00CB; B = 16'h00D0; #100;
A = 16'h00CB; B = 16'h00D1; #100;
A = 16'h00CB; B = 16'h00D2; #100;
A = 16'h00CB; B = 16'h00D3; #100;
A = 16'h00CB; B = 16'h00D4; #100;
A = 16'h00CB; B = 16'h00D5; #100;
A = 16'h00CB; B = 16'h00D6; #100;
A = 16'h00CB; B = 16'h00D7; #100;
A = 16'h00CB; B = 16'h00D8; #100;
A = 16'h00CB; B = 16'h00D9; #100;
A = 16'h00CB; B = 16'h00DA; #100;
A = 16'h00CB; B = 16'h00DB; #100;
A = 16'h00CB; B = 16'h00DC; #100;
A = 16'h00CB; B = 16'h00DD; #100;
A = 16'h00CB; B = 16'h00DE; #100;
A = 16'h00CB; B = 16'h00DF; #100;
A = 16'h00CB; B = 16'h00E0; #100;
A = 16'h00CB; B = 16'h00E1; #100;
A = 16'h00CB; B = 16'h00E2; #100;
A = 16'h00CB; B = 16'h00E3; #100;
A = 16'h00CB; B = 16'h00E4; #100;
A = 16'h00CB; B = 16'h00E5; #100;
A = 16'h00CB; B = 16'h00E6; #100;
A = 16'h00CB; B = 16'h00E7; #100;
A = 16'h00CB; B = 16'h00E8; #100;
A = 16'h00CB; B = 16'h00E9; #100;
A = 16'h00CB; B = 16'h00EA; #100;
A = 16'h00CB; B = 16'h00EB; #100;
A = 16'h00CB; B = 16'h00EC; #100;
A = 16'h00CB; B = 16'h00ED; #100;
A = 16'h00CB; B = 16'h00EE; #100;
A = 16'h00CB; B = 16'h00EF; #100;
A = 16'h00CB; B = 16'h00F0; #100;
A = 16'h00CB; B = 16'h00F1; #100;
A = 16'h00CB; B = 16'h00F2; #100;
A = 16'h00CB; B = 16'h00F3; #100;
A = 16'h00CB; B = 16'h00F4; #100;
A = 16'h00CB; B = 16'h00F5; #100;
A = 16'h00CB; B = 16'h00F6; #100;
A = 16'h00CB; B = 16'h00F7; #100;
A = 16'h00CB; B = 16'h00F8; #100;
A = 16'h00CB; B = 16'h00F9; #100;
A = 16'h00CB; B = 16'h00FA; #100;
A = 16'h00CB; B = 16'h00FB; #100;
A = 16'h00CB; B = 16'h00FC; #100;
A = 16'h00CB; B = 16'h00FD; #100;
A = 16'h00CB; B = 16'h00FE; #100;
A = 16'h00CB; B = 16'h00FF; #100;
A = 16'h00CC; B = 16'h000; #100;
A = 16'h00CC; B = 16'h001; #100;
A = 16'h00CC; B = 16'h002; #100;
A = 16'h00CC; B = 16'h003; #100;
A = 16'h00CC; B = 16'h004; #100;
A = 16'h00CC; B = 16'h005; #100;
A = 16'h00CC; B = 16'h006; #100;
A = 16'h00CC; B = 16'h007; #100;
A = 16'h00CC; B = 16'h008; #100;
A = 16'h00CC; B = 16'h009; #100;
A = 16'h00CC; B = 16'h00A; #100;
A = 16'h00CC; B = 16'h00B; #100;
A = 16'h00CC; B = 16'h00C; #100;
A = 16'h00CC; B = 16'h00D; #100;
A = 16'h00CC; B = 16'h00E; #100;
A = 16'h00CC; B = 16'h00F; #100;
A = 16'h00CC; B = 16'h0010; #100;
A = 16'h00CC; B = 16'h0011; #100;
A = 16'h00CC; B = 16'h0012; #100;
A = 16'h00CC; B = 16'h0013; #100;
A = 16'h00CC; B = 16'h0014; #100;
A = 16'h00CC; B = 16'h0015; #100;
A = 16'h00CC; B = 16'h0016; #100;
A = 16'h00CC; B = 16'h0017; #100;
A = 16'h00CC; B = 16'h0018; #100;
A = 16'h00CC; B = 16'h0019; #100;
A = 16'h00CC; B = 16'h001A; #100;
A = 16'h00CC; B = 16'h001B; #100;
A = 16'h00CC; B = 16'h001C; #100;
A = 16'h00CC; B = 16'h001D; #100;
A = 16'h00CC; B = 16'h001E; #100;
A = 16'h00CC; B = 16'h001F; #100;
A = 16'h00CC; B = 16'h0020; #100;
A = 16'h00CC; B = 16'h0021; #100;
A = 16'h00CC; B = 16'h0022; #100;
A = 16'h00CC; B = 16'h0023; #100;
A = 16'h00CC; B = 16'h0024; #100;
A = 16'h00CC; B = 16'h0025; #100;
A = 16'h00CC; B = 16'h0026; #100;
A = 16'h00CC; B = 16'h0027; #100;
A = 16'h00CC; B = 16'h0028; #100;
A = 16'h00CC; B = 16'h0029; #100;
A = 16'h00CC; B = 16'h002A; #100;
A = 16'h00CC; B = 16'h002B; #100;
A = 16'h00CC; B = 16'h002C; #100;
A = 16'h00CC; B = 16'h002D; #100;
A = 16'h00CC; B = 16'h002E; #100;
A = 16'h00CC; B = 16'h002F; #100;
A = 16'h00CC; B = 16'h0030; #100;
A = 16'h00CC; B = 16'h0031; #100;
A = 16'h00CC; B = 16'h0032; #100;
A = 16'h00CC; B = 16'h0033; #100;
A = 16'h00CC; B = 16'h0034; #100;
A = 16'h00CC; B = 16'h0035; #100;
A = 16'h00CC; B = 16'h0036; #100;
A = 16'h00CC; B = 16'h0037; #100;
A = 16'h00CC; B = 16'h0038; #100;
A = 16'h00CC; B = 16'h0039; #100;
A = 16'h00CC; B = 16'h003A; #100;
A = 16'h00CC; B = 16'h003B; #100;
A = 16'h00CC; B = 16'h003C; #100;
A = 16'h00CC; B = 16'h003D; #100;
A = 16'h00CC; B = 16'h003E; #100;
A = 16'h00CC; B = 16'h003F; #100;
A = 16'h00CC; B = 16'h0040; #100;
A = 16'h00CC; B = 16'h0041; #100;
A = 16'h00CC; B = 16'h0042; #100;
A = 16'h00CC; B = 16'h0043; #100;
A = 16'h00CC; B = 16'h0044; #100;
A = 16'h00CC; B = 16'h0045; #100;
A = 16'h00CC; B = 16'h0046; #100;
A = 16'h00CC; B = 16'h0047; #100;
A = 16'h00CC; B = 16'h0048; #100;
A = 16'h00CC; B = 16'h0049; #100;
A = 16'h00CC; B = 16'h004A; #100;
A = 16'h00CC; B = 16'h004B; #100;
A = 16'h00CC; B = 16'h004C; #100;
A = 16'h00CC; B = 16'h004D; #100;
A = 16'h00CC; B = 16'h004E; #100;
A = 16'h00CC; B = 16'h004F; #100;
A = 16'h00CC; B = 16'h0050; #100;
A = 16'h00CC; B = 16'h0051; #100;
A = 16'h00CC; B = 16'h0052; #100;
A = 16'h00CC; B = 16'h0053; #100;
A = 16'h00CC; B = 16'h0054; #100;
A = 16'h00CC; B = 16'h0055; #100;
A = 16'h00CC; B = 16'h0056; #100;
A = 16'h00CC; B = 16'h0057; #100;
A = 16'h00CC; B = 16'h0058; #100;
A = 16'h00CC; B = 16'h0059; #100;
A = 16'h00CC; B = 16'h005A; #100;
A = 16'h00CC; B = 16'h005B; #100;
A = 16'h00CC; B = 16'h005C; #100;
A = 16'h00CC; B = 16'h005D; #100;
A = 16'h00CC; B = 16'h005E; #100;
A = 16'h00CC; B = 16'h005F; #100;
A = 16'h00CC; B = 16'h0060; #100;
A = 16'h00CC; B = 16'h0061; #100;
A = 16'h00CC; B = 16'h0062; #100;
A = 16'h00CC; B = 16'h0063; #100;
A = 16'h00CC; B = 16'h0064; #100;
A = 16'h00CC; B = 16'h0065; #100;
A = 16'h00CC; B = 16'h0066; #100;
A = 16'h00CC; B = 16'h0067; #100;
A = 16'h00CC; B = 16'h0068; #100;
A = 16'h00CC; B = 16'h0069; #100;
A = 16'h00CC; B = 16'h006A; #100;
A = 16'h00CC; B = 16'h006B; #100;
A = 16'h00CC; B = 16'h006C; #100;
A = 16'h00CC; B = 16'h006D; #100;
A = 16'h00CC; B = 16'h006E; #100;
A = 16'h00CC; B = 16'h006F; #100;
A = 16'h00CC; B = 16'h0070; #100;
A = 16'h00CC; B = 16'h0071; #100;
A = 16'h00CC; B = 16'h0072; #100;
A = 16'h00CC; B = 16'h0073; #100;
A = 16'h00CC; B = 16'h0074; #100;
A = 16'h00CC; B = 16'h0075; #100;
A = 16'h00CC; B = 16'h0076; #100;
A = 16'h00CC; B = 16'h0077; #100;
A = 16'h00CC; B = 16'h0078; #100;
A = 16'h00CC; B = 16'h0079; #100;
A = 16'h00CC; B = 16'h007A; #100;
A = 16'h00CC; B = 16'h007B; #100;
A = 16'h00CC; B = 16'h007C; #100;
A = 16'h00CC; B = 16'h007D; #100;
A = 16'h00CC; B = 16'h007E; #100;
A = 16'h00CC; B = 16'h007F; #100;
A = 16'h00CC; B = 16'h0080; #100;
A = 16'h00CC; B = 16'h0081; #100;
A = 16'h00CC; B = 16'h0082; #100;
A = 16'h00CC; B = 16'h0083; #100;
A = 16'h00CC; B = 16'h0084; #100;
A = 16'h00CC; B = 16'h0085; #100;
A = 16'h00CC; B = 16'h0086; #100;
A = 16'h00CC; B = 16'h0087; #100;
A = 16'h00CC; B = 16'h0088; #100;
A = 16'h00CC; B = 16'h0089; #100;
A = 16'h00CC; B = 16'h008A; #100;
A = 16'h00CC; B = 16'h008B; #100;
A = 16'h00CC; B = 16'h008C; #100;
A = 16'h00CC; B = 16'h008D; #100;
A = 16'h00CC; B = 16'h008E; #100;
A = 16'h00CC; B = 16'h008F; #100;
A = 16'h00CC; B = 16'h0090; #100;
A = 16'h00CC; B = 16'h0091; #100;
A = 16'h00CC; B = 16'h0092; #100;
A = 16'h00CC; B = 16'h0093; #100;
A = 16'h00CC; B = 16'h0094; #100;
A = 16'h00CC; B = 16'h0095; #100;
A = 16'h00CC; B = 16'h0096; #100;
A = 16'h00CC; B = 16'h0097; #100;
A = 16'h00CC; B = 16'h0098; #100;
A = 16'h00CC; B = 16'h0099; #100;
A = 16'h00CC; B = 16'h009A; #100;
A = 16'h00CC; B = 16'h009B; #100;
A = 16'h00CC; B = 16'h009C; #100;
A = 16'h00CC; B = 16'h009D; #100;
A = 16'h00CC; B = 16'h009E; #100;
A = 16'h00CC; B = 16'h009F; #100;
A = 16'h00CC; B = 16'h00A0; #100;
A = 16'h00CC; B = 16'h00A1; #100;
A = 16'h00CC; B = 16'h00A2; #100;
A = 16'h00CC; B = 16'h00A3; #100;
A = 16'h00CC; B = 16'h00A4; #100;
A = 16'h00CC; B = 16'h00A5; #100;
A = 16'h00CC; B = 16'h00A6; #100;
A = 16'h00CC; B = 16'h00A7; #100;
A = 16'h00CC; B = 16'h00A8; #100;
A = 16'h00CC; B = 16'h00A9; #100;
A = 16'h00CC; B = 16'h00AA; #100;
A = 16'h00CC; B = 16'h00AB; #100;
A = 16'h00CC; B = 16'h00AC; #100;
A = 16'h00CC; B = 16'h00AD; #100;
A = 16'h00CC; B = 16'h00AE; #100;
A = 16'h00CC; B = 16'h00AF; #100;
A = 16'h00CC; B = 16'h00B0; #100;
A = 16'h00CC; B = 16'h00B1; #100;
A = 16'h00CC; B = 16'h00B2; #100;
A = 16'h00CC; B = 16'h00B3; #100;
A = 16'h00CC; B = 16'h00B4; #100;
A = 16'h00CC; B = 16'h00B5; #100;
A = 16'h00CC; B = 16'h00B6; #100;
A = 16'h00CC; B = 16'h00B7; #100;
A = 16'h00CC; B = 16'h00B8; #100;
A = 16'h00CC; B = 16'h00B9; #100;
A = 16'h00CC; B = 16'h00BA; #100;
A = 16'h00CC; B = 16'h00BB; #100;
A = 16'h00CC; B = 16'h00BC; #100;
A = 16'h00CC; B = 16'h00BD; #100;
A = 16'h00CC; B = 16'h00BE; #100;
A = 16'h00CC; B = 16'h00BF; #100;
A = 16'h00CC; B = 16'h00C0; #100;
A = 16'h00CC; B = 16'h00C1; #100;
A = 16'h00CC; B = 16'h00C2; #100;
A = 16'h00CC; B = 16'h00C3; #100;
A = 16'h00CC; B = 16'h00C4; #100;
A = 16'h00CC; B = 16'h00C5; #100;
A = 16'h00CC; B = 16'h00C6; #100;
A = 16'h00CC; B = 16'h00C7; #100;
A = 16'h00CC; B = 16'h00C8; #100;
A = 16'h00CC; B = 16'h00C9; #100;
A = 16'h00CC; B = 16'h00CA; #100;
A = 16'h00CC; B = 16'h00CB; #100;
A = 16'h00CC; B = 16'h00CC; #100;
A = 16'h00CC; B = 16'h00CD; #100;
A = 16'h00CC; B = 16'h00CE; #100;
A = 16'h00CC; B = 16'h00CF; #100;
A = 16'h00CC; B = 16'h00D0; #100;
A = 16'h00CC; B = 16'h00D1; #100;
A = 16'h00CC; B = 16'h00D2; #100;
A = 16'h00CC; B = 16'h00D3; #100;
A = 16'h00CC; B = 16'h00D4; #100;
A = 16'h00CC; B = 16'h00D5; #100;
A = 16'h00CC; B = 16'h00D6; #100;
A = 16'h00CC; B = 16'h00D7; #100;
A = 16'h00CC; B = 16'h00D8; #100;
A = 16'h00CC; B = 16'h00D9; #100;
A = 16'h00CC; B = 16'h00DA; #100;
A = 16'h00CC; B = 16'h00DB; #100;
A = 16'h00CC; B = 16'h00DC; #100;
A = 16'h00CC; B = 16'h00DD; #100;
A = 16'h00CC; B = 16'h00DE; #100;
A = 16'h00CC; B = 16'h00DF; #100;
A = 16'h00CC; B = 16'h00E0; #100;
A = 16'h00CC; B = 16'h00E1; #100;
A = 16'h00CC; B = 16'h00E2; #100;
A = 16'h00CC; B = 16'h00E3; #100;
A = 16'h00CC; B = 16'h00E4; #100;
A = 16'h00CC; B = 16'h00E5; #100;
A = 16'h00CC; B = 16'h00E6; #100;
A = 16'h00CC; B = 16'h00E7; #100;
A = 16'h00CC; B = 16'h00E8; #100;
A = 16'h00CC; B = 16'h00E9; #100;
A = 16'h00CC; B = 16'h00EA; #100;
A = 16'h00CC; B = 16'h00EB; #100;
A = 16'h00CC; B = 16'h00EC; #100;
A = 16'h00CC; B = 16'h00ED; #100;
A = 16'h00CC; B = 16'h00EE; #100;
A = 16'h00CC; B = 16'h00EF; #100;
A = 16'h00CC; B = 16'h00F0; #100;
A = 16'h00CC; B = 16'h00F1; #100;
A = 16'h00CC; B = 16'h00F2; #100;
A = 16'h00CC; B = 16'h00F3; #100;
A = 16'h00CC; B = 16'h00F4; #100;
A = 16'h00CC; B = 16'h00F5; #100;
A = 16'h00CC; B = 16'h00F6; #100;
A = 16'h00CC; B = 16'h00F7; #100;
A = 16'h00CC; B = 16'h00F8; #100;
A = 16'h00CC; B = 16'h00F9; #100;
A = 16'h00CC; B = 16'h00FA; #100;
A = 16'h00CC; B = 16'h00FB; #100;
A = 16'h00CC; B = 16'h00FC; #100;
A = 16'h00CC; B = 16'h00FD; #100;
A = 16'h00CC; B = 16'h00FE; #100;
A = 16'h00CC; B = 16'h00FF; #100;
A = 16'h00CD; B = 16'h000; #100;
A = 16'h00CD; B = 16'h001; #100;
A = 16'h00CD; B = 16'h002; #100;
A = 16'h00CD; B = 16'h003; #100;
A = 16'h00CD; B = 16'h004; #100;
A = 16'h00CD; B = 16'h005; #100;
A = 16'h00CD; B = 16'h006; #100;
A = 16'h00CD; B = 16'h007; #100;
A = 16'h00CD; B = 16'h008; #100;
A = 16'h00CD; B = 16'h009; #100;
A = 16'h00CD; B = 16'h00A; #100;
A = 16'h00CD; B = 16'h00B; #100;
A = 16'h00CD; B = 16'h00C; #100;
A = 16'h00CD; B = 16'h00D; #100;
A = 16'h00CD; B = 16'h00E; #100;
A = 16'h00CD; B = 16'h00F; #100;
A = 16'h00CD; B = 16'h0010; #100;
A = 16'h00CD; B = 16'h0011; #100;
A = 16'h00CD; B = 16'h0012; #100;
A = 16'h00CD; B = 16'h0013; #100;
A = 16'h00CD; B = 16'h0014; #100;
A = 16'h00CD; B = 16'h0015; #100;
A = 16'h00CD; B = 16'h0016; #100;
A = 16'h00CD; B = 16'h0017; #100;
A = 16'h00CD; B = 16'h0018; #100;
A = 16'h00CD; B = 16'h0019; #100;
A = 16'h00CD; B = 16'h001A; #100;
A = 16'h00CD; B = 16'h001B; #100;
A = 16'h00CD; B = 16'h001C; #100;
A = 16'h00CD; B = 16'h001D; #100;
A = 16'h00CD; B = 16'h001E; #100;
A = 16'h00CD; B = 16'h001F; #100;
A = 16'h00CD; B = 16'h0020; #100;
A = 16'h00CD; B = 16'h0021; #100;
A = 16'h00CD; B = 16'h0022; #100;
A = 16'h00CD; B = 16'h0023; #100;
A = 16'h00CD; B = 16'h0024; #100;
A = 16'h00CD; B = 16'h0025; #100;
A = 16'h00CD; B = 16'h0026; #100;
A = 16'h00CD; B = 16'h0027; #100;
A = 16'h00CD; B = 16'h0028; #100;
A = 16'h00CD; B = 16'h0029; #100;
A = 16'h00CD; B = 16'h002A; #100;
A = 16'h00CD; B = 16'h002B; #100;
A = 16'h00CD; B = 16'h002C; #100;
A = 16'h00CD; B = 16'h002D; #100;
A = 16'h00CD; B = 16'h002E; #100;
A = 16'h00CD; B = 16'h002F; #100;
A = 16'h00CD; B = 16'h0030; #100;
A = 16'h00CD; B = 16'h0031; #100;
A = 16'h00CD; B = 16'h0032; #100;
A = 16'h00CD; B = 16'h0033; #100;
A = 16'h00CD; B = 16'h0034; #100;
A = 16'h00CD; B = 16'h0035; #100;
A = 16'h00CD; B = 16'h0036; #100;
A = 16'h00CD; B = 16'h0037; #100;
A = 16'h00CD; B = 16'h0038; #100;
A = 16'h00CD; B = 16'h0039; #100;
A = 16'h00CD; B = 16'h003A; #100;
A = 16'h00CD; B = 16'h003B; #100;
A = 16'h00CD; B = 16'h003C; #100;
A = 16'h00CD; B = 16'h003D; #100;
A = 16'h00CD; B = 16'h003E; #100;
A = 16'h00CD; B = 16'h003F; #100;
A = 16'h00CD; B = 16'h0040; #100;
A = 16'h00CD; B = 16'h0041; #100;
A = 16'h00CD; B = 16'h0042; #100;
A = 16'h00CD; B = 16'h0043; #100;
A = 16'h00CD; B = 16'h0044; #100;
A = 16'h00CD; B = 16'h0045; #100;
A = 16'h00CD; B = 16'h0046; #100;
A = 16'h00CD; B = 16'h0047; #100;
A = 16'h00CD; B = 16'h0048; #100;
A = 16'h00CD; B = 16'h0049; #100;
A = 16'h00CD; B = 16'h004A; #100;
A = 16'h00CD; B = 16'h004B; #100;
A = 16'h00CD; B = 16'h004C; #100;
A = 16'h00CD; B = 16'h004D; #100;
A = 16'h00CD; B = 16'h004E; #100;
A = 16'h00CD; B = 16'h004F; #100;
A = 16'h00CD; B = 16'h0050; #100;
A = 16'h00CD; B = 16'h0051; #100;
A = 16'h00CD; B = 16'h0052; #100;
A = 16'h00CD; B = 16'h0053; #100;
A = 16'h00CD; B = 16'h0054; #100;
A = 16'h00CD; B = 16'h0055; #100;
A = 16'h00CD; B = 16'h0056; #100;
A = 16'h00CD; B = 16'h0057; #100;
A = 16'h00CD; B = 16'h0058; #100;
A = 16'h00CD; B = 16'h0059; #100;
A = 16'h00CD; B = 16'h005A; #100;
A = 16'h00CD; B = 16'h005B; #100;
A = 16'h00CD; B = 16'h005C; #100;
A = 16'h00CD; B = 16'h005D; #100;
A = 16'h00CD; B = 16'h005E; #100;
A = 16'h00CD; B = 16'h005F; #100;
A = 16'h00CD; B = 16'h0060; #100;
A = 16'h00CD; B = 16'h0061; #100;
A = 16'h00CD; B = 16'h0062; #100;
A = 16'h00CD; B = 16'h0063; #100;
A = 16'h00CD; B = 16'h0064; #100;
A = 16'h00CD; B = 16'h0065; #100;
A = 16'h00CD; B = 16'h0066; #100;
A = 16'h00CD; B = 16'h0067; #100;
A = 16'h00CD; B = 16'h0068; #100;
A = 16'h00CD; B = 16'h0069; #100;
A = 16'h00CD; B = 16'h006A; #100;
A = 16'h00CD; B = 16'h006B; #100;
A = 16'h00CD; B = 16'h006C; #100;
A = 16'h00CD; B = 16'h006D; #100;
A = 16'h00CD; B = 16'h006E; #100;
A = 16'h00CD; B = 16'h006F; #100;
A = 16'h00CD; B = 16'h0070; #100;
A = 16'h00CD; B = 16'h0071; #100;
A = 16'h00CD; B = 16'h0072; #100;
A = 16'h00CD; B = 16'h0073; #100;
A = 16'h00CD; B = 16'h0074; #100;
A = 16'h00CD; B = 16'h0075; #100;
A = 16'h00CD; B = 16'h0076; #100;
A = 16'h00CD; B = 16'h0077; #100;
A = 16'h00CD; B = 16'h0078; #100;
A = 16'h00CD; B = 16'h0079; #100;
A = 16'h00CD; B = 16'h007A; #100;
A = 16'h00CD; B = 16'h007B; #100;
A = 16'h00CD; B = 16'h007C; #100;
A = 16'h00CD; B = 16'h007D; #100;
A = 16'h00CD; B = 16'h007E; #100;
A = 16'h00CD; B = 16'h007F; #100;
A = 16'h00CD; B = 16'h0080; #100;
A = 16'h00CD; B = 16'h0081; #100;
A = 16'h00CD; B = 16'h0082; #100;
A = 16'h00CD; B = 16'h0083; #100;
A = 16'h00CD; B = 16'h0084; #100;
A = 16'h00CD; B = 16'h0085; #100;
A = 16'h00CD; B = 16'h0086; #100;
A = 16'h00CD; B = 16'h0087; #100;
A = 16'h00CD; B = 16'h0088; #100;
A = 16'h00CD; B = 16'h0089; #100;
A = 16'h00CD; B = 16'h008A; #100;
A = 16'h00CD; B = 16'h008B; #100;
A = 16'h00CD; B = 16'h008C; #100;
A = 16'h00CD; B = 16'h008D; #100;
A = 16'h00CD; B = 16'h008E; #100;
A = 16'h00CD; B = 16'h008F; #100;
A = 16'h00CD; B = 16'h0090; #100;
A = 16'h00CD; B = 16'h0091; #100;
A = 16'h00CD; B = 16'h0092; #100;
A = 16'h00CD; B = 16'h0093; #100;
A = 16'h00CD; B = 16'h0094; #100;
A = 16'h00CD; B = 16'h0095; #100;
A = 16'h00CD; B = 16'h0096; #100;
A = 16'h00CD; B = 16'h0097; #100;
A = 16'h00CD; B = 16'h0098; #100;
A = 16'h00CD; B = 16'h0099; #100;
A = 16'h00CD; B = 16'h009A; #100;
A = 16'h00CD; B = 16'h009B; #100;
A = 16'h00CD; B = 16'h009C; #100;
A = 16'h00CD; B = 16'h009D; #100;
A = 16'h00CD; B = 16'h009E; #100;
A = 16'h00CD; B = 16'h009F; #100;
A = 16'h00CD; B = 16'h00A0; #100;
A = 16'h00CD; B = 16'h00A1; #100;
A = 16'h00CD; B = 16'h00A2; #100;
A = 16'h00CD; B = 16'h00A3; #100;
A = 16'h00CD; B = 16'h00A4; #100;
A = 16'h00CD; B = 16'h00A5; #100;
A = 16'h00CD; B = 16'h00A6; #100;
A = 16'h00CD; B = 16'h00A7; #100;
A = 16'h00CD; B = 16'h00A8; #100;
A = 16'h00CD; B = 16'h00A9; #100;
A = 16'h00CD; B = 16'h00AA; #100;
A = 16'h00CD; B = 16'h00AB; #100;
A = 16'h00CD; B = 16'h00AC; #100;
A = 16'h00CD; B = 16'h00AD; #100;
A = 16'h00CD; B = 16'h00AE; #100;
A = 16'h00CD; B = 16'h00AF; #100;
A = 16'h00CD; B = 16'h00B0; #100;
A = 16'h00CD; B = 16'h00B1; #100;
A = 16'h00CD; B = 16'h00B2; #100;
A = 16'h00CD; B = 16'h00B3; #100;
A = 16'h00CD; B = 16'h00B4; #100;
A = 16'h00CD; B = 16'h00B5; #100;
A = 16'h00CD; B = 16'h00B6; #100;
A = 16'h00CD; B = 16'h00B7; #100;
A = 16'h00CD; B = 16'h00B8; #100;
A = 16'h00CD; B = 16'h00B9; #100;
A = 16'h00CD; B = 16'h00BA; #100;
A = 16'h00CD; B = 16'h00BB; #100;
A = 16'h00CD; B = 16'h00BC; #100;
A = 16'h00CD; B = 16'h00BD; #100;
A = 16'h00CD; B = 16'h00BE; #100;
A = 16'h00CD; B = 16'h00BF; #100;
A = 16'h00CD; B = 16'h00C0; #100;
A = 16'h00CD; B = 16'h00C1; #100;
A = 16'h00CD; B = 16'h00C2; #100;
A = 16'h00CD; B = 16'h00C3; #100;
A = 16'h00CD; B = 16'h00C4; #100;
A = 16'h00CD; B = 16'h00C5; #100;
A = 16'h00CD; B = 16'h00C6; #100;
A = 16'h00CD; B = 16'h00C7; #100;
A = 16'h00CD; B = 16'h00C8; #100;
A = 16'h00CD; B = 16'h00C9; #100;
A = 16'h00CD; B = 16'h00CA; #100;
A = 16'h00CD; B = 16'h00CB; #100;
A = 16'h00CD; B = 16'h00CC; #100;
A = 16'h00CD; B = 16'h00CD; #100;
A = 16'h00CD; B = 16'h00CE; #100;
A = 16'h00CD; B = 16'h00CF; #100;
A = 16'h00CD; B = 16'h00D0; #100;
A = 16'h00CD; B = 16'h00D1; #100;
A = 16'h00CD; B = 16'h00D2; #100;
A = 16'h00CD; B = 16'h00D3; #100;
A = 16'h00CD; B = 16'h00D4; #100;
A = 16'h00CD; B = 16'h00D5; #100;
A = 16'h00CD; B = 16'h00D6; #100;
A = 16'h00CD; B = 16'h00D7; #100;
A = 16'h00CD; B = 16'h00D8; #100;
A = 16'h00CD; B = 16'h00D9; #100;
A = 16'h00CD; B = 16'h00DA; #100;
A = 16'h00CD; B = 16'h00DB; #100;
A = 16'h00CD; B = 16'h00DC; #100;
A = 16'h00CD; B = 16'h00DD; #100;
A = 16'h00CD; B = 16'h00DE; #100;
A = 16'h00CD; B = 16'h00DF; #100;
A = 16'h00CD; B = 16'h00E0; #100;
A = 16'h00CD; B = 16'h00E1; #100;
A = 16'h00CD; B = 16'h00E2; #100;
A = 16'h00CD; B = 16'h00E3; #100;
A = 16'h00CD; B = 16'h00E4; #100;
A = 16'h00CD; B = 16'h00E5; #100;
A = 16'h00CD; B = 16'h00E6; #100;
A = 16'h00CD; B = 16'h00E7; #100;
A = 16'h00CD; B = 16'h00E8; #100;
A = 16'h00CD; B = 16'h00E9; #100;
A = 16'h00CD; B = 16'h00EA; #100;
A = 16'h00CD; B = 16'h00EB; #100;
A = 16'h00CD; B = 16'h00EC; #100;
A = 16'h00CD; B = 16'h00ED; #100;
A = 16'h00CD; B = 16'h00EE; #100;
A = 16'h00CD; B = 16'h00EF; #100;
A = 16'h00CD; B = 16'h00F0; #100;
A = 16'h00CD; B = 16'h00F1; #100;
A = 16'h00CD; B = 16'h00F2; #100;
A = 16'h00CD; B = 16'h00F3; #100;
A = 16'h00CD; B = 16'h00F4; #100;
A = 16'h00CD; B = 16'h00F5; #100;
A = 16'h00CD; B = 16'h00F6; #100;
A = 16'h00CD; B = 16'h00F7; #100;
A = 16'h00CD; B = 16'h00F8; #100;
A = 16'h00CD; B = 16'h00F9; #100;
A = 16'h00CD; B = 16'h00FA; #100;
A = 16'h00CD; B = 16'h00FB; #100;
A = 16'h00CD; B = 16'h00FC; #100;
A = 16'h00CD; B = 16'h00FD; #100;
A = 16'h00CD; B = 16'h00FE; #100;
A = 16'h00CD; B = 16'h00FF; #100;
A = 16'h00CE; B = 16'h000; #100;
A = 16'h00CE; B = 16'h001; #100;
A = 16'h00CE; B = 16'h002; #100;
A = 16'h00CE; B = 16'h003; #100;
A = 16'h00CE; B = 16'h004; #100;
A = 16'h00CE; B = 16'h005; #100;
A = 16'h00CE; B = 16'h006; #100;
A = 16'h00CE; B = 16'h007; #100;
A = 16'h00CE; B = 16'h008; #100;
A = 16'h00CE; B = 16'h009; #100;
A = 16'h00CE; B = 16'h00A; #100;
A = 16'h00CE; B = 16'h00B; #100;
A = 16'h00CE; B = 16'h00C; #100;
A = 16'h00CE; B = 16'h00D; #100;
A = 16'h00CE; B = 16'h00E; #100;
A = 16'h00CE; B = 16'h00F; #100;
A = 16'h00CE; B = 16'h0010; #100;
A = 16'h00CE; B = 16'h0011; #100;
A = 16'h00CE; B = 16'h0012; #100;
A = 16'h00CE; B = 16'h0013; #100;
A = 16'h00CE; B = 16'h0014; #100;
A = 16'h00CE; B = 16'h0015; #100;
A = 16'h00CE; B = 16'h0016; #100;
A = 16'h00CE; B = 16'h0017; #100;
A = 16'h00CE; B = 16'h0018; #100;
A = 16'h00CE; B = 16'h0019; #100;
A = 16'h00CE; B = 16'h001A; #100;
A = 16'h00CE; B = 16'h001B; #100;
A = 16'h00CE; B = 16'h001C; #100;
A = 16'h00CE; B = 16'h001D; #100;
A = 16'h00CE; B = 16'h001E; #100;
A = 16'h00CE; B = 16'h001F; #100;
A = 16'h00CE; B = 16'h0020; #100;
A = 16'h00CE; B = 16'h0021; #100;
A = 16'h00CE; B = 16'h0022; #100;
A = 16'h00CE; B = 16'h0023; #100;
A = 16'h00CE; B = 16'h0024; #100;
A = 16'h00CE; B = 16'h0025; #100;
A = 16'h00CE; B = 16'h0026; #100;
A = 16'h00CE; B = 16'h0027; #100;
A = 16'h00CE; B = 16'h0028; #100;
A = 16'h00CE; B = 16'h0029; #100;
A = 16'h00CE; B = 16'h002A; #100;
A = 16'h00CE; B = 16'h002B; #100;
A = 16'h00CE; B = 16'h002C; #100;
A = 16'h00CE; B = 16'h002D; #100;
A = 16'h00CE; B = 16'h002E; #100;
A = 16'h00CE; B = 16'h002F; #100;
A = 16'h00CE; B = 16'h0030; #100;
A = 16'h00CE; B = 16'h0031; #100;
A = 16'h00CE; B = 16'h0032; #100;
A = 16'h00CE; B = 16'h0033; #100;
A = 16'h00CE; B = 16'h0034; #100;
A = 16'h00CE; B = 16'h0035; #100;
A = 16'h00CE; B = 16'h0036; #100;
A = 16'h00CE; B = 16'h0037; #100;
A = 16'h00CE; B = 16'h0038; #100;
A = 16'h00CE; B = 16'h0039; #100;
A = 16'h00CE; B = 16'h003A; #100;
A = 16'h00CE; B = 16'h003B; #100;
A = 16'h00CE; B = 16'h003C; #100;
A = 16'h00CE; B = 16'h003D; #100;
A = 16'h00CE; B = 16'h003E; #100;
A = 16'h00CE; B = 16'h003F; #100;
A = 16'h00CE; B = 16'h0040; #100;
A = 16'h00CE; B = 16'h0041; #100;
A = 16'h00CE; B = 16'h0042; #100;
A = 16'h00CE; B = 16'h0043; #100;
A = 16'h00CE; B = 16'h0044; #100;
A = 16'h00CE; B = 16'h0045; #100;
A = 16'h00CE; B = 16'h0046; #100;
A = 16'h00CE; B = 16'h0047; #100;
A = 16'h00CE; B = 16'h0048; #100;
A = 16'h00CE; B = 16'h0049; #100;
A = 16'h00CE; B = 16'h004A; #100;
A = 16'h00CE; B = 16'h004B; #100;
A = 16'h00CE; B = 16'h004C; #100;
A = 16'h00CE; B = 16'h004D; #100;
A = 16'h00CE; B = 16'h004E; #100;
A = 16'h00CE; B = 16'h004F; #100;
A = 16'h00CE; B = 16'h0050; #100;
A = 16'h00CE; B = 16'h0051; #100;
A = 16'h00CE; B = 16'h0052; #100;
A = 16'h00CE; B = 16'h0053; #100;
A = 16'h00CE; B = 16'h0054; #100;
A = 16'h00CE; B = 16'h0055; #100;
A = 16'h00CE; B = 16'h0056; #100;
A = 16'h00CE; B = 16'h0057; #100;
A = 16'h00CE; B = 16'h0058; #100;
A = 16'h00CE; B = 16'h0059; #100;
A = 16'h00CE; B = 16'h005A; #100;
A = 16'h00CE; B = 16'h005B; #100;
A = 16'h00CE; B = 16'h005C; #100;
A = 16'h00CE; B = 16'h005D; #100;
A = 16'h00CE; B = 16'h005E; #100;
A = 16'h00CE; B = 16'h005F; #100;
A = 16'h00CE; B = 16'h0060; #100;
A = 16'h00CE; B = 16'h0061; #100;
A = 16'h00CE; B = 16'h0062; #100;
A = 16'h00CE; B = 16'h0063; #100;
A = 16'h00CE; B = 16'h0064; #100;
A = 16'h00CE; B = 16'h0065; #100;
A = 16'h00CE; B = 16'h0066; #100;
A = 16'h00CE; B = 16'h0067; #100;
A = 16'h00CE; B = 16'h0068; #100;
A = 16'h00CE; B = 16'h0069; #100;
A = 16'h00CE; B = 16'h006A; #100;
A = 16'h00CE; B = 16'h006B; #100;
A = 16'h00CE; B = 16'h006C; #100;
A = 16'h00CE; B = 16'h006D; #100;
A = 16'h00CE; B = 16'h006E; #100;
A = 16'h00CE; B = 16'h006F; #100;
A = 16'h00CE; B = 16'h0070; #100;
A = 16'h00CE; B = 16'h0071; #100;
A = 16'h00CE; B = 16'h0072; #100;
A = 16'h00CE; B = 16'h0073; #100;
A = 16'h00CE; B = 16'h0074; #100;
A = 16'h00CE; B = 16'h0075; #100;
A = 16'h00CE; B = 16'h0076; #100;
A = 16'h00CE; B = 16'h0077; #100;
A = 16'h00CE; B = 16'h0078; #100;
A = 16'h00CE; B = 16'h0079; #100;
A = 16'h00CE; B = 16'h007A; #100;
A = 16'h00CE; B = 16'h007B; #100;
A = 16'h00CE; B = 16'h007C; #100;
A = 16'h00CE; B = 16'h007D; #100;
A = 16'h00CE; B = 16'h007E; #100;
A = 16'h00CE; B = 16'h007F; #100;
A = 16'h00CE; B = 16'h0080; #100;
A = 16'h00CE; B = 16'h0081; #100;
A = 16'h00CE; B = 16'h0082; #100;
A = 16'h00CE; B = 16'h0083; #100;
A = 16'h00CE; B = 16'h0084; #100;
A = 16'h00CE; B = 16'h0085; #100;
A = 16'h00CE; B = 16'h0086; #100;
A = 16'h00CE; B = 16'h0087; #100;
A = 16'h00CE; B = 16'h0088; #100;
A = 16'h00CE; B = 16'h0089; #100;
A = 16'h00CE; B = 16'h008A; #100;
A = 16'h00CE; B = 16'h008B; #100;
A = 16'h00CE; B = 16'h008C; #100;
A = 16'h00CE; B = 16'h008D; #100;
A = 16'h00CE; B = 16'h008E; #100;
A = 16'h00CE; B = 16'h008F; #100;
A = 16'h00CE; B = 16'h0090; #100;
A = 16'h00CE; B = 16'h0091; #100;
A = 16'h00CE; B = 16'h0092; #100;
A = 16'h00CE; B = 16'h0093; #100;
A = 16'h00CE; B = 16'h0094; #100;
A = 16'h00CE; B = 16'h0095; #100;
A = 16'h00CE; B = 16'h0096; #100;
A = 16'h00CE; B = 16'h0097; #100;
A = 16'h00CE; B = 16'h0098; #100;
A = 16'h00CE; B = 16'h0099; #100;
A = 16'h00CE; B = 16'h009A; #100;
A = 16'h00CE; B = 16'h009B; #100;
A = 16'h00CE; B = 16'h009C; #100;
A = 16'h00CE; B = 16'h009D; #100;
A = 16'h00CE; B = 16'h009E; #100;
A = 16'h00CE; B = 16'h009F; #100;
A = 16'h00CE; B = 16'h00A0; #100;
A = 16'h00CE; B = 16'h00A1; #100;
A = 16'h00CE; B = 16'h00A2; #100;
A = 16'h00CE; B = 16'h00A3; #100;
A = 16'h00CE; B = 16'h00A4; #100;
A = 16'h00CE; B = 16'h00A5; #100;
A = 16'h00CE; B = 16'h00A6; #100;
A = 16'h00CE; B = 16'h00A7; #100;
A = 16'h00CE; B = 16'h00A8; #100;
A = 16'h00CE; B = 16'h00A9; #100;
A = 16'h00CE; B = 16'h00AA; #100;
A = 16'h00CE; B = 16'h00AB; #100;
A = 16'h00CE; B = 16'h00AC; #100;
A = 16'h00CE; B = 16'h00AD; #100;
A = 16'h00CE; B = 16'h00AE; #100;
A = 16'h00CE; B = 16'h00AF; #100;
A = 16'h00CE; B = 16'h00B0; #100;
A = 16'h00CE; B = 16'h00B1; #100;
A = 16'h00CE; B = 16'h00B2; #100;
A = 16'h00CE; B = 16'h00B3; #100;
A = 16'h00CE; B = 16'h00B4; #100;
A = 16'h00CE; B = 16'h00B5; #100;
A = 16'h00CE; B = 16'h00B6; #100;
A = 16'h00CE; B = 16'h00B7; #100;
A = 16'h00CE; B = 16'h00B8; #100;
A = 16'h00CE; B = 16'h00B9; #100;
A = 16'h00CE; B = 16'h00BA; #100;
A = 16'h00CE; B = 16'h00BB; #100;
A = 16'h00CE; B = 16'h00BC; #100;
A = 16'h00CE; B = 16'h00BD; #100;
A = 16'h00CE; B = 16'h00BE; #100;
A = 16'h00CE; B = 16'h00BF; #100;
A = 16'h00CE; B = 16'h00C0; #100;
A = 16'h00CE; B = 16'h00C1; #100;
A = 16'h00CE; B = 16'h00C2; #100;
A = 16'h00CE; B = 16'h00C3; #100;
A = 16'h00CE; B = 16'h00C4; #100;
A = 16'h00CE; B = 16'h00C5; #100;
A = 16'h00CE; B = 16'h00C6; #100;
A = 16'h00CE; B = 16'h00C7; #100;
A = 16'h00CE; B = 16'h00C8; #100;
A = 16'h00CE; B = 16'h00C9; #100;
A = 16'h00CE; B = 16'h00CA; #100;
A = 16'h00CE; B = 16'h00CB; #100;
A = 16'h00CE; B = 16'h00CC; #100;
A = 16'h00CE; B = 16'h00CD; #100;
A = 16'h00CE; B = 16'h00CE; #100;
A = 16'h00CE; B = 16'h00CF; #100;
A = 16'h00CE; B = 16'h00D0; #100;
A = 16'h00CE; B = 16'h00D1; #100;
A = 16'h00CE; B = 16'h00D2; #100;
A = 16'h00CE; B = 16'h00D3; #100;
A = 16'h00CE; B = 16'h00D4; #100;
A = 16'h00CE; B = 16'h00D5; #100;
A = 16'h00CE; B = 16'h00D6; #100;
A = 16'h00CE; B = 16'h00D7; #100;
A = 16'h00CE; B = 16'h00D8; #100;
A = 16'h00CE; B = 16'h00D9; #100;
A = 16'h00CE; B = 16'h00DA; #100;
A = 16'h00CE; B = 16'h00DB; #100;
A = 16'h00CE; B = 16'h00DC; #100;
A = 16'h00CE; B = 16'h00DD; #100;
A = 16'h00CE; B = 16'h00DE; #100;
A = 16'h00CE; B = 16'h00DF; #100;
A = 16'h00CE; B = 16'h00E0; #100;
A = 16'h00CE; B = 16'h00E1; #100;
A = 16'h00CE; B = 16'h00E2; #100;
A = 16'h00CE; B = 16'h00E3; #100;
A = 16'h00CE; B = 16'h00E4; #100;
A = 16'h00CE; B = 16'h00E5; #100;
A = 16'h00CE; B = 16'h00E6; #100;
A = 16'h00CE; B = 16'h00E7; #100;
A = 16'h00CE; B = 16'h00E8; #100;
A = 16'h00CE; B = 16'h00E9; #100;
A = 16'h00CE; B = 16'h00EA; #100;
A = 16'h00CE; B = 16'h00EB; #100;
A = 16'h00CE; B = 16'h00EC; #100;
A = 16'h00CE; B = 16'h00ED; #100;
A = 16'h00CE; B = 16'h00EE; #100;
A = 16'h00CE; B = 16'h00EF; #100;
A = 16'h00CE; B = 16'h00F0; #100;
A = 16'h00CE; B = 16'h00F1; #100;
A = 16'h00CE; B = 16'h00F2; #100;
A = 16'h00CE; B = 16'h00F3; #100;
A = 16'h00CE; B = 16'h00F4; #100;
A = 16'h00CE; B = 16'h00F5; #100;
A = 16'h00CE; B = 16'h00F6; #100;
A = 16'h00CE; B = 16'h00F7; #100;
A = 16'h00CE; B = 16'h00F8; #100;
A = 16'h00CE; B = 16'h00F9; #100;
A = 16'h00CE; B = 16'h00FA; #100;
A = 16'h00CE; B = 16'h00FB; #100;
A = 16'h00CE; B = 16'h00FC; #100;
A = 16'h00CE; B = 16'h00FD; #100;
A = 16'h00CE; B = 16'h00FE; #100;
A = 16'h00CE; B = 16'h00FF; #100;
A = 16'h00CF; B = 16'h000; #100;
A = 16'h00CF; B = 16'h001; #100;
A = 16'h00CF; B = 16'h002; #100;
A = 16'h00CF; B = 16'h003; #100;
A = 16'h00CF; B = 16'h004; #100;
A = 16'h00CF; B = 16'h005; #100;
A = 16'h00CF; B = 16'h006; #100;
A = 16'h00CF; B = 16'h007; #100;
A = 16'h00CF; B = 16'h008; #100;
A = 16'h00CF; B = 16'h009; #100;
A = 16'h00CF; B = 16'h00A; #100;
A = 16'h00CF; B = 16'h00B; #100;
A = 16'h00CF; B = 16'h00C; #100;
A = 16'h00CF; B = 16'h00D; #100;
A = 16'h00CF; B = 16'h00E; #100;
A = 16'h00CF; B = 16'h00F; #100;
A = 16'h00CF; B = 16'h0010; #100;
A = 16'h00CF; B = 16'h0011; #100;
A = 16'h00CF; B = 16'h0012; #100;
A = 16'h00CF; B = 16'h0013; #100;
A = 16'h00CF; B = 16'h0014; #100;
A = 16'h00CF; B = 16'h0015; #100;
A = 16'h00CF; B = 16'h0016; #100;
A = 16'h00CF; B = 16'h0017; #100;
A = 16'h00CF; B = 16'h0018; #100;
A = 16'h00CF; B = 16'h0019; #100;
A = 16'h00CF; B = 16'h001A; #100;
A = 16'h00CF; B = 16'h001B; #100;
A = 16'h00CF; B = 16'h001C; #100;
A = 16'h00CF; B = 16'h001D; #100;
A = 16'h00CF; B = 16'h001E; #100;
A = 16'h00CF; B = 16'h001F; #100;
A = 16'h00CF; B = 16'h0020; #100;
A = 16'h00CF; B = 16'h0021; #100;
A = 16'h00CF; B = 16'h0022; #100;
A = 16'h00CF; B = 16'h0023; #100;
A = 16'h00CF; B = 16'h0024; #100;
A = 16'h00CF; B = 16'h0025; #100;
A = 16'h00CF; B = 16'h0026; #100;
A = 16'h00CF; B = 16'h0027; #100;
A = 16'h00CF; B = 16'h0028; #100;
A = 16'h00CF; B = 16'h0029; #100;
A = 16'h00CF; B = 16'h002A; #100;
A = 16'h00CF; B = 16'h002B; #100;
A = 16'h00CF; B = 16'h002C; #100;
A = 16'h00CF; B = 16'h002D; #100;
A = 16'h00CF; B = 16'h002E; #100;
A = 16'h00CF; B = 16'h002F; #100;
A = 16'h00CF; B = 16'h0030; #100;
A = 16'h00CF; B = 16'h0031; #100;
A = 16'h00CF; B = 16'h0032; #100;
A = 16'h00CF; B = 16'h0033; #100;
A = 16'h00CF; B = 16'h0034; #100;
A = 16'h00CF; B = 16'h0035; #100;
A = 16'h00CF; B = 16'h0036; #100;
A = 16'h00CF; B = 16'h0037; #100;
A = 16'h00CF; B = 16'h0038; #100;
A = 16'h00CF; B = 16'h0039; #100;
A = 16'h00CF; B = 16'h003A; #100;
A = 16'h00CF; B = 16'h003B; #100;
A = 16'h00CF; B = 16'h003C; #100;
A = 16'h00CF; B = 16'h003D; #100;
A = 16'h00CF; B = 16'h003E; #100;
A = 16'h00CF; B = 16'h003F; #100;
A = 16'h00CF; B = 16'h0040; #100;
A = 16'h00CF; B = 16'h0041; #100;
A = 16'h00CF; B = 16'h0042; #100;
A = 16'h00CF; B = 16'h0043; #100;
A = 16'h00CF; B = 16'h0044; #100;
A = 16'h00CF; B = 16'h0045; #100;
A = 16'h00CF; B = 16'h0046; #100;
A = 16'h00CF; B = 16'h0047; #100;
A = 16'h00CF; B = 16'h0048; #100;
A = 16'h00CF; B = 16'h0049; #100;
A = 16'h00CF; B = 16'h004A; #100;
A = 16'h00CF; B = 16'h004B; #100;
A = 16'h00CF; B = 16'h004C; #100;
A = 16'h00CF; B = 16'h004D; #100;
A = 16'h00CF; B = 16'h004E; #100;
A = 16'h00CF; B = 16'h004F; #100;
A = 16'h00CF; B = 16'h0050; #100;
A = 16'h00CF; B = 16'h0051; #100;
A = 16'h00CF; B = 16'h0052; #100;
A = 16'h00CF; B = 16'h0053; #100;
A = 16'h00CF; B = 16'h0054; #100;
A = 16'h00CF; B = 16'h0055; #100;
A = 16'h00CF; B = 16'h0056; #100;
A = 16'h00CF; B = 16'h0057; #100;
A = 16'h00CF; B = 16'h0058; #100;
A = 16'h00CF; B = 16'h0059; #100;
A = 16'h00CF; B = 16'h005A; #100;
A = 16'h00CF; B = 16'h005B; #100;
A = 16'h00CF; B = 16'h005C; #100;
A = 16'h00CF; B = 16'h005D; #100;
A = 16'h00CF; B = 16'h005E; #100;
A = 16'h00CF; B = 16'h005F; #100;
A = 16'h00CF; B = 16'h0060; #100;
A = 16'h00CF; B = 16'h0061; #100;
A = 16'h00CF; B = 16'h0062; #100;
A = 16'h00CF; B = 16'h0063; #100;
A = 16'h00CF; B = 16'h0064; #100;
A = 16'h00CF; B = 16'h0065; #100;
A = 16'h00CF; B = 16'h0066; #100;
A = 16'h00CF; B = 16'h0067; #100;
A = 16'h00CF; B = 16'h0068; #100;
A = 16'h00CF; B = 16'h0069; #100;
A = 16'h00CF; B = 16'h006A; #100;
A = 16'h00CF; B = 16'h006B; #100;
A = 16'h00CF; B = 16'h006C; #100;
A = 16'h00CF; B = 16'h006D; #100;
A = 16'h00CF; B = 16'h006E; #100;
A = 16'h00CF; B = 16'h006F; #100;
A = 16'h00CF; B = 16'h0070; #100;
A = 16'h00CF; B = 16'h0071; #100;
A = 16'h00CF; B = 16'h0072; #100;
A = 16'h00CF; B = 16'h0073; #100;
A = 16'h00CF; B = 16'h0074; #100;
A = 16'h00CF; B = 16'h0075; #100;
A = 16'h00CF; B = 16'h0076; #100;
A = 16'h00CF; B = 16'h0077; #100;
A = 16'h00CF; B = 16'h0078; #100;
A = 16'h00CF; B = 16'h0079; #100;
A = 16'h00CF; B = 16'h007A; #100;
A = 16'h00CF; B = 16'h007B; #100;
A = 16'h00CF; B = 16'h007C; #100;
A = 16'h00CF; B = 16'h007D; #100;
A = 16'h00CF; B = 16'h007E; #100;
A = 16'h00CF; B = 16'h007F; #100;
A = 16'h00CF; B = 16'h0080; #100;
A = 16'h00CF; B = 16'h0081; #100;
A = 16'h00CF; B = 16'h0082; #100;
A = 16'h00CF; B = 16'h0083; #100;
A = 16'h00CF; B = 16'h0084; #100;
A = 16'h00CF; B = 16'h0085; #100;
A = 16'h00CF; B = 16'h0086; #100;
A = 16'h00CF; B = 16'h0087; #100;
A = 16'h00CF; B = 16'h0088; #100;
A = 16'h00CF; B = 16'h0089; #100;
A = 16'h00CF; B = 16'h008A; #100;
A = 16'h00CF; B = 16'h008B; #100;
A = 16'h00CF; B = 16'h008C; #100;
A = 16'h00CF; B = 16'h008D; #100;
A = 16'h00CF; B = 16'h008E; #100;
A = 16'h00CF; B = 16'h008F; #100;
A = 16'h00CF; B = 16'h0090; #100;
A = 16'h00CF; B = 16'h0091; #100;
A = 16'h00CF; B = 16'h0092; #100;
A = 16'h00CF; B = 16'h0093; #100;
A = 16'h00CF; B = 16'h0094; #100;
A = 16'h00CF; B = 16'h0095; #100;
A = 16'h00CF; B = 16'h0096; #100;
A = 16'h00CF; B = 16'h0097; #100;
A = 16'h00CF; B = 16'h0098; #100;
A = 16'h00CF; B = 16'h0099; #100;
A = 16'h00CF; B = 16'h009A; #100;
A = 16'h00CF; B = 16'h009B; #100;
A = 16'h00CF; B = 16'h009C; #100;
A = 16'h00CF; B = 16'h009D; #100;
A = 16'h00CF; B = 16'h009E; #100;
A = 16'h00CF; B = 16'h009F; #100;
A = 16'h00CF; B = 16'h00A0; #100;
A = 16'h00CF; B = 16'h00A1; #100;
A = 16'h00CF; B = 16'h00A2; #100;
A = 16'h00CF; B = 16'h00A3; #100;
A = 16'h00CF; B = 16'h00A4; #100;
A = 16'h00CF; B = 16'h00A5; #100;
A = 16'h00CF; B = 16'h00A6; #100;
A = 16'h00CF; B = 16'h00A7; #100;
A = 16'h00CF; B = 16'h00A8; #100;
A = 16'h00CF; B = 16'h00A9; #100;
A = 16'h00CF; B = 16'h00AA; #100;
A = 16'h00CF; B = 16'h00AB; #100;
A = 16'h00CF; B = 16'h00AC; #100;
A = 16'h00CF; B = 16'h00AD; #100;
A = 16'h00CF; B = 16'h00AE; #100;
A = 16'h00CF; B = 16'h00AF; #100;
A = 16'h00CF; B = 16'h00B0; #100;
A = 16'h00CF; B = 16'h00B1; #100;
A = 16'h00CF; B = 16'h00B2; #100;
A = 16'h00CF; B = 16'h00B3; #100;
A = 16'h00CF; B = 16'h00B4; #100;
A = 16'h00CF; B = 16'h00B5; #100;
A = 16'h00CF; B = 16'h00B6; #100;
A = 16'h00CF; B = 16'h00B7; #100;
A = 16'h00CF; B = 16'h00B8; #100;
A = 16'h00CF; B = 16'h00B9; #100;
A = 16'h00CF; B = 16'h00BA; #100;
A = 16'h00CF; B = 16'h00BB; #100;
A = 16'h00CF; B = 16'h00BC; #100;
A = 16'h00CF; B = 16'h00BD; #100;
A = 16'h00CF; B = 16'h00BE; #100;
A = 16'h00CF; B = 16'h00BF; #100;
A = 16'h00CF; B = 16'h00C0; #100;
A = 16'h00CF; B = 16'h00C1; #100;
A = 16'h00CF; B = 16'h00C2; #100;
A = 16'h00CF; B = 16'h00C3; #100;
A = 16'h00CF; B = 16'h00C4; #100;
A = 16'h00CF; B = 16'h00C5; #100;
A = 16'h00CF; B = 16'h00C6; #100;
A = 16'h00CF; B = 16'h00C7; #100;
A = 16'h00CF; B = 16'h00C8; #100;
A = 16'h00CF; B = 16'h00C9; #100;
A = 16'h00CF; B = 16'h00CA; #100;
A = 16'h00CF; B = 16'h00CB; #100;
A = 16'h00CF; B = 16'h00CC; #100;
A = 16'h00CF; B = 16'h00CD; #100;
A = 16'h00CF; B = 16'h00CE; #100;
A = 16'h00CF; B = 16'h00CF; #100;
A = 16'h00CF; B = 16'h00D0; #100;
A = 16'h00CF; B = 16'h00D1; #100;
A = 16'h00CF; B = 16'h00D2; #100;
A = 16'h00CF; B = 16'h00D3; #100;
A = 16'h00CF; B = 16'h00D4; #100;
A = 16'h00CF; B = 16'h00D5; #100;
A = 16'h00CF; B = 16'h00D6; #100;
A = 16'h00CF; B = 16'h00D7; #100;
A = 16'h00CF; B = 16'h00D8; #100;
A = 16'h00CF; B = 16'h00D9; #100;
A = 16'h00CF; B = 16'h00DA; #100;
A = 16'h00CF; B = 16'h00DB; #100;
A = 16'h00CF; B = 16'h00DC; #100;
A = 16'h00CF; B = 16'h00DD; #100;
A = 16'h00CF; B = 16'h00DE; #100;
A = 16'h00CF; B = 16'h00DF; #100;
A = 16'h00CF; B = 16'h00E0; #100;
A = 16'h00CF; B = 16'h00E1; #100;
A = 16'h00CF; B = 16'h00E2; #100;
A = 16'h00CF; B = 16'h00E3; #100;
A = 16'h00CF; B = 16'h00E4; #100;
A = 16'h00CF; B = 16'h00E5; #100;
A = 16'h00CF; B = 16'h00E6; #100;
A = 16'h00CF; B = 16'h00E7; #100;
A = 16'h00CF; B = 16'h00E8; #100;
A = 16'h00CF; B = 16'h00E9; #100;
A = 16'h00CF; B = 16'h00EA; #100;
A = 16'h00CF; B = 16'h00EB; #100;
A = 16'h00CF; B = 16'h00EC; #100;
A = 16'h00CF; B = 16'h00ED; #100;
A = 16'h00CF; B = 16'h00EE; #100;
A = 16'h00CF; B = 16'h00EF; #100;
A = 16'h00CF; B = 16'h00F0; #100;
A = 16'h00CF; B = 16'h00F1; #100;
A = 16'h00CF; B = 16'h00F2; #100;
A = 16'h00CF; B = 16'h00F3; #100;
A = 16'h00CF; B = 16'h00F4; #100;
A = 16'h00CF; B = 16'h00F5; #100;
A = 16'h00CF; B = 16'h00F6; #100;
A = 16'h00CF; B = 16'h00F7; #100;
A = 16'h00CF; B = 16'h00F8; #100;
A = 16'h00CF; B = 16'h00F9; #100;
A = 16'h00CF; B = 16'h00FA; #100;
A = 16'h00CF; B = 16'h00FB; #100;
A = 16'h00CF; B = 16'h00FC; #100;
A = 16'h00CF; B = 16'h00FD; #100;
A = 16'h00CF; B = 16'h00FE; #100;
A = 16'h00CF; B = 16'h00FF; #100;
A = 16'h00D0; B = 16'h000; #100;
A = 16'h00D0; B = 16'h001; #100;
A = 16'h00D0; B = 16'h002; #100;
A = 16'h00D0; B = 16'h003; #100;
A = 16'h00D0; B = 16'h004; #100;
A = 16'h00D0; B = 16'h005; #100;
A = 16'h00D0; B = 16'h006; #100;
A = 16'h00D0; B = 16'h007; #100;
A = 16'h00D0; B = 16'h008; #100;
A = 16'h00D0; B = 16'h009; #100;
A = 16'h00D0; B = 16'h00A; #100;
A = 16'h00D0; B = 16'h00B; #100;
A = 16'h00D0; B = 16'h00C; #100;
A = 16'h00D0; B = 16'h00D; #100;
A = 16'h00D0; B = 16'h00E; #100;
A = 16'h00D0; B = 16'h00F; #100;
A = 16'h00D0; B = 16'h0010; #100;
A = 16'h00D0; B = 16'h0011; #100;
A = 16'h00D0; B = 16'h0012; #100;
A = 16'h00D0; B = 16'h0013; #100;
A = 16'h00D0; B = 16'h0014; #100;
A = 16'h00D0; B = 16'h0015; #100;
A = 16'h00D0; B = 16'h0016; #100;
A = 16'h00D0; B = 16'h0017; #100;
A = 16'h00D0; B = 16'h0018; #100;
A = 16'h00D0; B = 16'h0019; #100;
A = 16'h00D0; B = 16'h001A; #100;
A = 16'h00D0; B = 16'h001B; #100;
A = 16'h00D0; B = 16'h001C; #100;
A = 16'h00D0; B = 16'h001D; #100;
A = 16'h00D0; B = 16'h001E; #100;
A = 16'h00D0; B = 16'h001F; #100;
A = 16'h00D0; B = 16'h0020; #100;
A = 16'h00D0; B = 16'h0021; #100;
A = 16'h00D0; B = 16'h0022; #100;
A = 16'h00D0; B = 16'h0023; #100;
A = 16'h00D0; B = 16'h0024; #100;
A = 16'h00D0; B = 16'h0025; #100;
A = 16'h00D0; B = 16'h0026; #100;
A = 16'h00D0; B = 16'h0027; #100;
A = 16'h00D0; B = 16'h0028; #100;
A = 16'h00D0; B = 16'h0029; #100;
A = 16'h00D0; B = 16'h002A; #100;
A = 16'h00D0; B = 16'h002B; #100;
A = 16'h00D0; B = 16'h002C; #100;
A = 16'h00D0; B = 16'h002D; #100;
A = 16'h00D0; B = 16'h002E; #100;
A = 16'h00D0; B = 16'h002F; #100;
A = 16'h00D0; B = 16'h0030; #100;
A = 16'h00D0; B = 16'h0031; #100;
A = 16'h00D0; B = 16'h0032; #100;
A = 16'h00D0; B = 16'h0033; #100;
A = 16'h00D0; B = 16'h0034; #100;
A = 16'h00D0; B = 16'h0035; #100;
A = 16'h00D0; B = 16'h0036; #100;
A = 16'h00D0; B = 16'h0037; #100;
A = 16'h00D0; B = 16'h0038; #100;
A = 16'h00D0; B = 16'h0039; #100;
A = 16'h00D0; B = 16'h003A; #100;
A = 16'h00D0; B = 16'h003B; #100;
A = 16'h00D0; B = 16'h003C; #100;
A = 16'h00D0; B = 16'h003D; #100;
A = 16'h00D0; B = 16'h003E; #100;
A = 16'h00D0; B = 16'h003F; #100;
A = 16'h00D0; B = 16'h0040; #100;
A = 16'h00D0; B = 16'h0041; #100;
A = 16'h00D0; B = 16'h0042; #100;
A = 16'h00D0; B = 16'h0043; #100;
A = 16'h00D0; B = 16'h0044; #100;
A = 16'h00D0; B = 16'h0045; #100;
A = 16'h00D0; B = 16'h0046; #100;
A = 16'h00D0; B = 16'h0047; #100;
A = 16'h00D0; B = 16'h0048; #100;
A = 16'h00D0; B = 16'h0049; #100;
A = 16'h00D0; B = 16'h004A; #100;
A = 16'h00D0; B = 16'h004B; #100;
A = 16'h00D0; B = 16'h004C; #100;
A = 16'h00D0; B = 16'h004D; #100;
A = 16'h00D0; B = 16'h004E; #100;
A = 16'h00D0; B = 16'h004F; #100;
A = 16'h00D0; B = 16'h0050; #100;
A = 16'h00D0; B = 16'h0051; #100;
A = 16'h00D0; B = 16'h0052; #100;
A = 16'h00D0; B = 16'h0053; #100;
A = 16'h00D0; B = 16'h0054; #100;
A = 16'h00D0; B = 16'h0055; #100;
A = 16'h00D0; B = 16'h0056; #100;
A = 16'h00D0; B = 16'h0057; #100;
A = 16'h00D0; B = 16'h0058; #100;
A = 16'h00D0; B = 16'h0059; #100;
A = 16'h00D0; B = 16'h005A; #100;
A = 16'h00D0; B = 16'h005B; #100;
A = 16'h00D0; B = 16'h005C; #100;
A = 16'h00D0; B = 16'h005D; #100;
A = 16'h00D0; B = 16'h005E; #100;
A = 16'h00D0; B = 16'h005F; #100;
A = 16'h00D0; B = 16'h0060; #100;
A = 16'h00D0; B = 16'h0061; #100;
A = 16'h00D0; B = 16'h0062; #100;
A = 16'h00D0; B = 16'h0063; #100;
A = 16'h00D0; B = 16'h0064; #100;
A = 16'h00D0; B = 16'h0065; #100;
A = 16'h00D0; B = 16'h0066; #100;
A = 16'h00D0; B = 16'h0067; #100;
A = 16'h00D0; B = 16'h0068; #100;
A = 16'h00D0; B = 16'h0069; #100;
A = 16'h00D0; B = 16'h006A; #100;
A = 16'h00D0; B = 16'h006B; #100;
A = 16'h00D0; B = 16'h006C; #100;
A = 16'h00D0; B = 16'h006D; #100;
A = 16'h00D0; B = 16'h006E; #100;
A = 16'h00D0; B = 16'h006F; #100;
A = 16'h00D0; B = 16'h0070; #100;
A = 16'h00D0; B = 16'h0071; #100;
A = 16'h00D0; B = 16'h0072; #100;
A = 16'h00D0; B = 16'h0073; #100;
A = 16'h00D0; B = 16'h0074; #100;
A = 16'h00D0; B = 16'h0075; #100;
A = 16'h00D0; B = 16'h0076; #100;
A = 16'h00D0; B = 16'h0077; #100;
A = 16'h00D0; B = 16'h0078; #100;
A = 16'h00D0; B = 16'h0079; #100;
A = 16'h00D0; B = 16'h007A; #100;
A = 16'h00D0; B = 16'h007B; #100;
A = 16'h00D0; B = 16'h007C; #100;
A = 16'h00D0; B = 16'h007D; #100;
A = 16'h00D0; B = 16'h007E; #100;
A = 16'h00D0; B = 16'h007F; #100;
A = 16'h00D0; B = 16'h0080; #100;
A = 16'h00D0; B = 16'h0081; #100;
A = 16'h00D0; B = 16'h0082; #100;
A = 16'h00D0; B = 16'h0083; #100;
A = 16'h00D0; B = 16'h0084; #100;
A = 16'h00D0; B = 16'h0085; #100;
A = 16'h00D0; B = 16'h0086; #100;
A = 16'h00D0; B = 16'h0087; #100;
A = 16'h00D0; B = 16'h0088; #100;
A = 16'h00D0; B = 16'h0089; #100;
A = 16'h00D0; B = 16'h008A; #100;
A = 16'h00D0; B = 16'h008B; #100;
A = 16'h00D0; B = 16'h008C; #100;
A = 16'h00D0; B = 16'h008D; #100;
A = 16'h00D0; B = 16'h008E; #100;
A = 16'h00D0; B = 16'h008F; #100;
A = 16'h00D0; B = 16'h0090; #100;
A = 16'h00D0; B = 16'h0091; #100;
A = 16'h00D0; B = 16'h0092; #100;
A = 16'h00D0; B = 16'h0093; #100;
A = 16'h00D0; B = 16'h0094; #100;
A = 16'h00D0; B = 16'h0095; #100;
A = 16'h00D0; B = 16'h0096; #100;
A = 16'h00D0; B = 16'h0097; #100;
A = 16'h00D0; B = 16'h0098; #100;
A = 16'h00D0; B = 16'h0099; #100;
A = 16'h00D0; B = 16'h009A; #100;
A = 16'h00D0; B = 16'h009B; #100;
A = 16'h00D0; B = 16'h009C; #100;
A = 16'h00D0; B = 16'h009D; #100;
A = 16'h00D0; B = 16'h009E; #100;
A = 16'h00D0; B = 16'h009F; #100;
A = 16'h00D0; B = 16'h00A0; #100;
A = 16'h00D0; B = 16'h00A1; #100;
A = 16'h00D0; B = 16'h00A2; #100;
A = 16'h00D0; B = 16'h00A3; #100;
A = 16'h00D0; B = 16'h00A4; #100;
A = 16'h00D0; B = 16'h00A5; #100;
A = 16'h00D0; B = 16'h00A6; #100;
A = 16'h00D0; B = 16'h00A7; #100;
A = 16'h00D0; B = 16'h00A8; #100;
A = 16'h00D0; B = 16'h00A9; #100;
A = 16'h00D0; B = 16'h00AA; #100;
A = 16'h00D0; B = 16'h00AB; #100;
A = 16'h00D0; B = 16'h00AC; #100;
A = 16'h00D0; B = 16'h00AD; #100;
A = 16'h00D0; B = 16'h00AE; #100;
A = 16'h00D0; B = 16'h00AF; #100;
A = 16'h00D0; B = 16'h00B0; #100;
A = 16'h00D0; B = 16'h00B1; #100;
A = 16'h00D0; B = 16'h00B2; #100;
A = 16'h00D0; B = 16'h00B3; #100;
A = 16'h00D0; B = 16'h00B4; #100;
A = 16'h00D0; B = 16'h00B5; #100;
A = 16'h00D0; B = 16'h00B6; #100;
A = 16'h00D0; B = 16'h00B7; #100;
A = 16'h00D0; B = 16'h00B8; #100;
A = 16'h00D0; B = 16'h00B9; #100;
A = 16'h00D0; B = 16'h00BA; #100;
A = 16'h00D0; B = 16'h00BB; #100;
A = 16'h00D0; B = 16'h00BC; #100;
A = 16'h00D0; B = 16'h00BD; #100;
A = 16'h00D0; B = 16'h00BE; #100;
A = 16'h00D0; B = 16'h00BF; #100;
A = 16'h00D0; B = 16'h00C0; #100;
A = 16'h00D0; B = 16'h00C1; #100;
A = 16'h00D0; B = 16'h00C2; #100;
A = 16'h00D0; B = 16'h00C3; #100;
A = 16'h00D0; B = 16'h00C4; #100;
A = 16'h00D0; B = 16'h00C5; #100;
A = 16'h00D0; B = 16'h00C6; #100;
A = 16'h00D0; B = 16'h00C7; #100;
A = 16'h00D0; B = 16'h00C8; #100;
A = 16'h00D0; B = 16'h00C9; #100;
A = 16'h00D0; B = 16'h00CA; #100;
A = 16'h00D0; B = 16'h00CB; #100;
A = 16'h00D0; B = 16'h00CC; #100;
A = 16'h00D0; B = 16'h00CD; #100;
A = 16'h00D0; B = 16'h00CE; #100;
A = 16'h00D0; B = 16'h00CF; #100;
A = 16'h00D0; B = 16'h00D0; #100;
A = 16'h00D0; B = 16'h00D1; #100;
A = 16'h00D0; B = 16'h00D2; #100;
A = 16'h00D0; B = 16'h00D3; #100;
A = 16'h00D0; B = 16'h00D4; #100;
A = 16'h00D0; B = 16'h00D5; #100;
A = 16'h00D0; B = 16'h00D6; #100;
A = 16'h00D0; B = 16'h00D7; #100;
A = 16'h00D0; B = 16'h00D8; #100;
A = 16'h00D0; B = 16'h00D9; #100;
A = 16'h00D0; B = 16'h00DA; #100;
A = 16'h00D0; B = 16'h00DB; #100;
A = 16'h00D0; B = 16'h00DC; #100;
A = 16'h00D0; B = 16'h00DD; #100;
A = 16'h00D0; B = 16'h00DE; #100;
A = 16'h00D0; B = 16'h00DF; #100;
A = 16'h00D0; B = 16'h00E0; #100;
A = 16'h00D0; B = 16'h00E1; #100;
A = 16'h00D0; B = 16'h00E2; #100;
A = 16'h00D0; B = 16'h00E3; #100;
A = 16'h00D0; B = 16'h00E4; #100;
A = 16'h00D0; B = 16'h00E5; #100;
A = 16'h00D0; B = 16'h00E6; #100;
A = 16'h00D0; B = 16'h00E7; #100;
A = 16'h00D0; B = 16'h00E8; #100;
A = 16'h00D0; B = 16'h00E9; #100;
A = 16'h00D0; B = 16'h00EA; #100;
A = 16'h00D0; B = 16'h00EB; #100;
A = 16'h00D0; B = 16'h00EC; #100;
A = 16'h00D0; B = 16'h00ED; #100;
A = 16'h00D0; B = 16'h00EE; #100;
A = 16'h00D0; B = 16'h00EF; #100;
A = 16'h00D0; B = 16'h00F0; #100;
A = 16'h00D0; B = 16'h00F1; #100;
A = 16'h00D0; B = 16'h00F2; #100;
A = 16'h00D0; B = 16'h00F3; #100;
A = 16'h00D0; B = 16'h00F4; #100;
A = 16'h00D0; B = 16'h00F5; #100;
A = 16'h00D0; B = 16'h00F6; #100;
A = 16'h00D0; B = 16'h00F7; #100;
A = 16'h00D0; B = 16'h00F8; #100;
A = 16'h00D0; B = 16'h00F9; #100;
A = 16'h00D0; B = 16'h00FA; #100;
A = 16'h00D0; B = 16'h00FB; #100;
A = 16'h00D0; B = 16'h00FC; #100;
A = 16'h00D0; B = 16'h00FD; #100;
A = 16'h00D0; B = 16'h00FE; #100;
A = 16'h00D0; B = 16'h00FF; #100;
A = 16'h00D1; B = 16'h000; #100;
A = 16'h00D1; B = 16'h001; #100;
A = 16'h00D1; B = 16'h002; #100;
A = 16'h00D1; B = 16'h003; #100;
A = 16'h00D1; B = 16'h004; #100;
A = 16'h00D1; B = 16'h005; #100;
A = 16'h00D1; B = 16'h006; #100;
A = 16'h00D1; B = 16'h007; #100;
A = 16'h00D1; B = 16'h008; #100;
A = 16'h00D1; B = 16'h009; #100;
A = 16'h00D1; B = 16'h00A; #100;
A = 16'h00D1; B = 16'h00B; #100;
A = 16'h00D1; B = 16'h00C; #100;
A = 16'h00D1; B = 16'h00D; #100;
A = 16'h00D1; B = 16'h00E; #100;
A = 16'h00D1; B = 16'h00F; #100;
A = 16'h00D1; B = 16'h0010; #100;
A = 16'h00D1; B = 16'h0011; #100;
A = 16'h00D1; B = 16'h0012; #100;
A = 16'h00D1; B = 16'h0013; #100;
A = 16'h00D1; B = 16'h0014; #100;
A = 16'h00D1; B = 16'h0015; #100;
A = 16'h00D1; B = 16'h0016; #100;
A = 16'h00D1; B = 16'h0017; #100;
A = 16'h00D1; B = 16'h0018; #100;
A = 16'h00D1; B = 16'h0019; #100;
A = 16'h00D1; B = 16'h001A; #100;
A = 16'h00D1; B = 16'h001B; #100;
A = 16'h00D1; B = 16'h001C; #100;
A = 16'h00D1; B = 16'h001D; #100;
A = 16'h00D1; B = 16'h001E; #100;
A = 16'h00D1; B = 16'h001F; #100;
A = 16'h00D1; B = 16'h0020; #100;
A = 16'h00D1; B = 16'h0021; #100;
A = 16'h00D1; B = 16'h0022; #100;
A = 16'h00D1; B = 16'h0023; #100;
A = 16'h00D1; B = 16'h0024; #100;
A = 16'h00D1; B = 16'h0025; #100;
A = 16'h00D1; B = 16'h0026; #100;
A = 16'h00D1; B = 16'h0027; #100;
A = 16'h00D1; B = 16'h0028; #100;
A = 16'h00D1; B = 16'h0029; #100;
A = 16'h00D1; B = 16'h002A; #100;
A = 16'h00D1; B = 16'h002B; #100;
A = 16'h00D1; B = 16'h002C; #100;
A = 16'h00D1; B = 16'h002D; #100;
A = 16'h00D1; B = 16'h002E; #100;
A = 16'h00D1; B = 16'h002F; #100;
A = 16'h00D1; B = 16'h0030; #100;
A = 16'h00D1; B = 16'h0031; #100;
A = 16'h00D1; B = 16'h0032; #100;
A = 16'h00D1; B = 16'h0033; #100;
A = 16'h00D1; B = 16'h0034; #100;
A = 16'h00D1; B = 16'h0035; #100;
A = 16'h00D1; B = 16'h0036; #100;
A = 16'h00D1; B = 16'h0037; #100;
A = 16'h00D1; B = 16'h0038; #100;
A = 16'h00D1; B = 16'h0039; #100;
A = 16'h00D1; B = 16'h003A; #100;
A = 16'h00D1; B = 16'h003B; #100;
A = 16'h00D1; B = 16'h003C; #100;
A = 16'h00D1; B = 16'h003D; #100;
A = 16'h00D1; B = 16'h003E; #100;
A = 16'h00D1; B = 16'h003F; #100;
A = 16'h00D1; B = 16'h0040; #100;
A = 16'h00D1; B = 16'h0041; #100;
A = 16'h00D1; B = 16'h0042; #100;
A = 16'h00D1; B = 16'h0043; #100;
A = 16'h00D1; B = 16'h0044; #100;
A = 16'h00D1; B = 16'h0045; #100;
A = 16'h00D1; B = 16'h0046; #100;
A = 16'h00D1; B = 16'h0047; #100;
A = 16'h00D1; B = 16'h0048; #100;
A = 16'h00D1; B = 16'h0049; #100;
A = 16'h00D1; B = 16'h004A; #100;
A = 16'h00D1; B = 16'h004B; #100;
A = 16'h00D1; B = 16'h004C; #100;
A = 16'h00D1; B = 16'h004D; #100;
A = 16'h00D1; B = 16'h004E; #100;
A = 16'h00D1; B = 16'h004F; #100;
A = 16'h00D1; B = 16'h0050; #100;
A = 16'h00D1; B = 16'h0051; #100;
A = 16'h00D1; B = 16'h0052; #100;
A = 16'h00D1; B = 16'h0053; #100;
A = 16'h00D1; B = 16'h0054; #100;
A = 16'h00D1; B = 16'h0055; #100;
A = 16'h00D1; B = 16'h0056; #100;
A = 16'h00D1; B = 16'h0057; #100;
A = 16'h00D1; B = 16'h0058; #100;
A = 16'h00D1; B = 16'h0059; #100;
A = 16'h00D1; B = 16'h005A; #100;
A = 16'h00D1; B = 16'h005B; #100;
A = 16'h00D1; B = 16'h005C; #100;
A = 16'h00D1; B = 16'h005D; #100;
A = 16'h00D1; B = 16'h005E; #100;
A = 16'h00D1; B = 16'h005F; #100;
A = 16'h00D1; B = 16'h0060; #100;
A = 16'h00D1; B = 16'h0061; #100;
A = 16'h00D1; B = 16'h0062; #100;
A = 16'h00D1; B = 16'h0063; #100;
A = 16'h00D1; B = 16'h0064; #100;
A = 16'h00D1; B = 16'h0065; #100;
A = 16'h00D1; B = 16'h0066; #100;
A = 16'h00D1; B = 16'h0067; #100;
A = 16'h00D1; B = 16'h0068; #100;
A = 16'h00D1; B = 16'h0069; #100;
A = 16'h00D1; B = 16'h006A; #100;
A = 16'h00D1; B = 16'h006B; #100;
A = 16'h00D1; B = 16'h006C; #100;
A = 16'h00D1; B = 16'h006D; #100;
A = 16'h00D1; B = 16'h006E; #100;
A = 16'h00D1; B = 16'h006F; #100;
A = 16'h00D1; B = 16'h0070; #100;
A = 16'h00D1; B = 16'h0071; #100;
A = 16'h00D1; B = 16'h0072; #100;
A = 16'h00D1; B = 16'h0073; #100;
A = 16'h00D1; B = 16'h0074; #100;
A = 16'h00D1; B = 16'h0075; #100;
A = 16'h00D1; B = 16'h0076; #100;
A = 16'h00D1; B = 16'h0077; #100;
A = 16'h00D1; B = 16'h0078; #100;
A = 16'h00D1; B = 16'h0079; #100;
A = 16'h00D1; B = 16'h007A; #100;
A = 16'h00D1; B = 16'h007B; #100;
A = 16'h00D1; B = 16'h007C; #100;
A = 16'h00D1; B = 16'h007D; #100;
A = 16'h00D1; B = 16'h007E; #100;
A = 16'h00D1; B = 16'h007F; #100;
A = 16'h00D1; B = 16'h0080; #100;
A = 16'h00D1; B = 16'h0081; #100;
A = 16'h00D1; B = 16'h0082; #100;
A = 16'h00D1; B = 16'h0083; #100;
A = 16'h00D1; B = 16'h0084; #100;
A = 16'h00D1; B = 16'h0085; #100;
A = 16'h00D1; B = 16'h0086; #100;
A = 16'h00D1; B = 16'h0087; #100;
A = 16'h00D1; B = 16'h0088; #100;
A = 16'h00D1; B = 16'h0089; #100;
A = 16'h00D1; B = 16'h008A; #100;
A = 16'h00D1; B = 16'h008B; #100;
A = 16'h00D1; B = 16'h008C; #100;
A = 16'h00D1; B = 16'h008D; #100;
A = 16'h00D1; B = 16'h008E; #100;
A = 16'h00D1; B = 16'h008F; #100;
A = 16'h00D1; B = 16'h0090; #100;
A = 16'h00D1; B = 16'h0091; #100;
A = 16'h00D1; B = 16'h0092; #100;
A = 16'h00D1; B = 16'h0093; #100;
A = 16'h00D1; B = 16'h0094; #100;
A = 16'h00D1; B = 16'h0095; #100;
A = 16'h00D1; B = 16'h0096; #100;
A = 16'h00D1; B = 16'h0097; #100;
A = 16'h00D1; B = 16'h0098; #100;
A = 16'h00D1; B = 16'h0099; #100;
A = 16'h00D1; B = 16'h009A; #100;
A = 16'h00D1; B = 16'h009B; #100;
A = 16'h00D1; B = 16'h009C; #100;
A = 16'h00D1; B = 16'h009D; #100;
A = 16'h00D1; B = 16'h009E; #100;
A = 16'h00D1; B = 16'h009F; #100;
A = 16'h00D1; B = 16'h00A0; #100;
A = 16'h00D1; B = 16'h00A1; #100;
A = 16'h00D1; B = 16'h00A2; #100;
A = 16'h00D1; B = 16'h00A3; #100;
A = 16'h00D1; B = 16'h00A4; #100;
A = 16'h00D1; B = 16'h00A5; #100;
A = 16'h00D1; B = 16'h00A6; #100;
A = 16'h00D1; B = 16'h00A7; #100;
A = 16'h00D1; B = 16'h00A8; #100;
A = 16'h00D1; B = 16'h00A9; #100;
A = 16'h00D1; B = 16'h00AA; #100;
A = 16'h00D1; B = 16'h00AB; #100;
A = 16'h00D1; B = 16'h00AC; #100;
A = 16'h00D1; B = 16'h00AD; #100;
A = 16'h00D1; B = 16'h00AE; #100;
A = 16'h00D1; B = 16'h00AF; #100;
A = 16'h00D1; B = 16'h00B0; #100;
A = 16'h00D1; B = 16'h00B1; #100;
A = 16'h00D1; B = 16'h00B2; #100;
A = 16'h00D1; B = 16'h00B3; #100;
A = 16'h00D1; B = 16'h00B4; #100;
A = 16'h00D1; B = 16'h00B5; #100;
A = 16'h00D1; B = 16'h00B6; #100;
A = 16'h00D1; B = 16'h00B7; #100;
A = 16'h00D1; B = 16'h00B8; #100;
A = 16'h00D1; B = 16'h00B9; #100;
A = 16'h00D1; B = 16'h00BA; #100;
A = 16'h00D1; B = 16'h00BB; #100;
A = 16'h00D1; B = 16'h00BC; #100;
A = 16'h00D1; B = 16'h00BD; #100;
A = 16'h00D1; B = 16'h00BE; #100;
A = 16'h00D1; B = 16'h00BF; #100;
A = 16'h00D1; B = 16'h00C0; #100;
A = 16'h00D1; B = 16'h00C1; #100;
A = 16'h00D1; B = 16'h00C2; #100;
A = 16'h00D1; B = 16'h00C3; #100;
A = 16'h00D1; B = 16'h00C4; #100;
A = 16'h00D1; B = 16'h00C5; #100;
A = 16'h00D1; B = 16'h00C6; #100;
A = 16'h00D1; B = 16'h00C7; #100;
A = 16'h00D1; B = 16'h00C8; #100;
A = 16'h00D1; B = 16'h00C9; #100;
A = 16'h00D1; B = 16'h00CA; #100;
A = 16'h00D1; B = 16'h00CB; #100;
A = 16'h00D1; B = 16'h00CC; #100;
A = 16'h00D1; B = 16'h00CD; #100;
A = 16'h00D1; B = 16'h00CE; #100;
A = 16'h00D1; B = 16'h00CF; #100;
A = 16'h00D1; B = 16'h00D0; #100;
A = 16'h00D1; B = 16'h00D1; #100;
A = 16'h00D1; B = 16'h00D2; #100;
A = 16'h00D1; B = 16'h00D3; #100;
A = 16'h00D1; B = 16'h00D4; #100;
A = 16'h00D1; B = 16'h00D5; #100;
A = 16'h00D1; B = 16'h00D6; #100;
A = 16'h00D1; B = 16'h00D7; #100;
A = 16'h00D1; B = 16'h00D8; #100;
A = 16'h00D1; B = 16'h00D9; #100;
A = 16'h00D1; B = 16'h00DA; #100;
A = 16'h00D1; B = 16'h00DB; #100;
A = 16'h00D1; B = 16'h00DC; #100;
A = 16'h00D1; B = 16'h00DD; #100;
A = 16'h00D1; B = 16'h00DE; #100;
A = 16'h00D1; B = 16'h00DF; #100;
A = 16'h00D1; B = 16'h00E0; #100;
A = 16'h00D1; B = 16'h00E1; #100;
A = 16'h00D1; B = 16'h00E2; #100;
A = 16'h00D1; B = 16'h00E3; #100;
A = 16'h00D1; B = 16'h00E4; #100;
A = 16'h00D1; B = 16'h00E5; #100;
A = 16'h00D1; B = 16'h00E6; #100;
A = 16'h00D1; B = 16'h00E7; #100;
A = 16'h00D1; B = 16'h00E8; #100;
A = 16'h00D1; B = 16'h00E9; #100;
A = 16'h00D1; B = 16'h00EA; #100;
A = 16'h00D1; B = 16'h00EB; #100;
A = 16'h00D1; B = 16'h00EC; #100;
A = 16'h00D1; B = 16'h00ED; #100;
A = 16'h00D1; B = 16'h00EE; #100;
A = 16'h00D1; B = 16'h00EF; #100;
A = 16'h00D1; B = 16'h00F0; #100;
A = 16'h00D1; B = 16'h00F1; #100;
A = 16'h00D1; B = 16'h00F2; #100;
A = 16'h00D1; B = 16'h00F3; #100;
A = 16'h00D1; B = 16'h00F4; #100;
A = 16'h00D1; B = 16'h00F5; #100;
A = 16'h00D1; B = 16'h00F6; #100;
A = 16'h00D1; B = 16'h00F7; #100;
A = 16'h00D1; B = 16'h00F8; #100;
A = 16'h00D1; B = 16'h00F9; #100;
A = 16'h00D1; B = 16'h00FA; #100;
A = 16'h00D1; B = 16'h00FB; #100;
A = 16'h00D1; B = 16'h00FC; #100;
A = 16'h00D1; B = 16'h00FD; #100;
A = 16'h00D1; B = 16'h00FE; #100;
A = 16'h00D1; B = 16'h00FF; #100;
A = 16'h00D2; B = 16'h000; #100;
A = 16'h00D2; B = 16'h001; #100;
A = 16'h00D2; B = 16'h002; #100;
A = 16'h00D2; B = 16'h003; #100;
A = 16'h00D2; B = 16'h004; #100;
A = 16'h00D2; B = 16'h005; #100;
A = 16'h00D2; B = 16'h006; #100;
A = 16'h00D2; B = 16'h007; #100;
A = 16'h00D2; B = 16'h008; #100;
A = 16'h00D2; B = 16'h009; #100;
A = 16'h00D2; B = 16'h00A; #100;
A = 16'h00D2; B = 16'h00B; #100;
A = 16'h00D2; B = 16'h00C; #100;
A = 16'h00D2; B = 16'h00D; #100;
A = 16'h00D2; B = 16'h00E; #100;
A = 16'h00D2; B = 16'h00F; #100;
A = 16'h00D2; B = 16'h0010; #100;
A = 16'h00D2; B = 16'h0011; #100;
A = 16'h00D2; B = 16'h0012; #100;
A = 16'h00D2; B = 16'h0013; #100;
A = 16'h00D2; B = 16'h0014; #100;
A = 16'h00D2; B = 16'h0015; #100;
A = 16'h00D2; B = 16'h0016; #100;
A = 16'h00D2; B = 16'h0017; #100;
A = 16'h00D2; B = 16'h0018; #100;
A = 16'h00D2; B = 16'h0019; #100;
A = 16'h00D2; B = 16'h001A; #100;
A = 16'h00D2; B = 16'h001B; #100;
A = 16'h00D2; B = 16'h001C; #100;
A = 16'h00D2; B = 16'h001D; #100;
A = 16'h00D2; B = 16'h001E; #100;
A = 16'h00D2; B = 16'h001F; #100;
A = 16'h00D2; B = 16'h0020; #100;
A = 16'h00D2; B = 16'h0021; #100;
A = 16'h00D2; B = 16'h0022; #100;
A = 16'h00D2; B = 16'h0023; #100;
A = 16'h00D2; B = 16'h0024; #100;
A = 16'h00D2; B = 16'h0025; #100;
A = 16'h00D2; B = 16'h0026; #100;
A = 16'h00D2; B = 16'h0027; #100;
A = 16'h00D2; B = 16'h0028; #100;
A = 16'h00D2; B = 16'h0029; #100;
A = 16'h00D2; B = 16'h002A; #100;
A = 16'h00D2; B = 16'h002B; #100;
A = 16'h00D2; B = 16'h002C; #100;
A = 16'h00D2; B = 16'h002D; #100;
A = 16'h00D2; B = 16'h002E; #100;
A = 16'h00D2; B = 16'h002F; #100;
A = 16'h00D2; B = 16'h0030; #100;
A = 16'h00D2; B = 16'h0031; #100;
A = 16'h00D2; B = 16'h0032; #100;
A = 16'h00D2; B = 16'h0033; #100;
A = 16'h00D2; B = 16'h0034; #100;
A = 16'h00D2; B = 16'h0035; #100;
A = 16'h00D2; B = 16'h0036; #100;
A = 16'h00D2; B = 16'h0037; #100;
A = 16'h00D2; B = 16'h0038; #100;
A = 16'h00D2; B = 16'h0039; #100;
A = 16'h00D2; B = 16'h003A; #100;
A = 16'h00D2; B = 16'h003B; #100;
A = 16'h00D2; B = 16'h003C; #100;
A = 16'h00D2; B = 16'h003D; #100;
A = 16'h00D2; B = 16'h003E; #100;
A = 16'h00D2; B = 16'h003F; #100;
A = 16'h00D2; B = 16'h0040; #100;
A = 16'h00D2; B = 16'h0041; #100;
A = 16'h00D2; B = 16'h0042; #100;
A = 16'h00D2; B = 16'h0043; #100;
A = 16'h00D2; B = 16'h0044; #100;
A = 16'h00D2; B = 16'h0045; #100;
A = 16'h00D2; B = 16'h0046; #100;
A = 16'h00D2; B = 16'h0047; #100;
A = 16'h00D2; B = 16'h0048; #100;
A = 16'h00D2; B = 16'h0049; #100;
A = 16'h00D2; B = 16'h004A; #100;
A = 16'h00D2; B = 16'h004B; #100;
A = 16'h00D2; B = 16'h004C; #100;
A = 16'h00D2; B = 16'h004D; #100;
A = 16'h00D2; B = 16'h004E; #100;
A = 16'h00D2; B = 16'h004F; #100;
A = 16'h00D2; B = 16'h0050; #100;
A = 16'h00D2; B = 16'h0051; #100;
A = 16'h00D2; B = 16'h0052; #100;
A = 16'h00D2; B = 16'h0053; #100;
A = 16'h00D2; B = 16'h0054; #100;
A = 16'h00D2; B = 16'h0055; #100;
A = 16'h00D2; B = 16'h0056; #100;
A = 16'h00D2; B = 16'h0057; #100;
A = 16'h00D2; B = 16'h0058; #100;
A = 16'h00D2; B = 16'h0059; #100;
A = 16'h00D2; B = 16'h005A; #100;
A = 16'h00D2; B = 16'h005B; #100;
A = 16'h00D2; B = 16'h005C; #100;
A = 16'h00D2; B = 16'h005D; #100;
A = 16'h00D2; B = 16'h005E; #100;
A = 16'h00D2; B = 16'h005F; #100;
A = 16'h00D2; B = 16'h0060; #100;
A = 16'h00D2; B = 16'h0061; #100;
A = 16'h00D2; B = 16'h0062; #100;
A = 16'h00D2; B = 16'h0063; #100;
A = 16'h00D2; B = 16'h0064; #100;
A = 16'h00D2; B = 16'h0065; #100;
A = 16'h00D2; B = 16'h0066; #100;
A = 16'h00D2; B = 16'h0067; #100;
A = 16'h00D2; B = 16'h0068; #100;
A = 16'h00D2; B = 16'h0069; #100;
A = 16'h00D2; B = 16'h006A; #100;
A = 16'h00D2; B = 16'h006B; #100;
A = 16'h00D2; B = 16'h006C; #100;
A = 16'h00D2; B = 16'h006D; #100;
A = 16'h00D2; B = 16'h006E; #100;
A = 16'h00D2; B = 16'h006F; #100;
A = 16'h00D2; B = 16'h0070; #100;
A = 16'h00D2; B = 16'h0071; #100;
A = 16'h00D2; B = 16'h0072; #100;
A = 16'h00D2; B = 16'h0073; #100;
A = 16'h00D2; B = 16'h0074; #100;
A = 16'h00D2; B = 16'h0075; #100;
A = 16'h00D2; B = 16'h0076; #100;
A = 16'h00D2; B = 16'h0077; #100;
A = 16'h00D2; B = 16'h0078; #100;
A = 16'h00D2; B = 16'h0079; #100;
A = 16'h00D2; B = 16'h007A; #100;
A = 16'h00D2; B = 16'h007B; #100;
A = 16'h00D2; B = 16'h007C; #100;
A = 16'h00D2; B = 16'h007D; #100;
A = 16'h00D2; B = 16'h007E; #100;
A = 16'h00D2; B = 16'h007F; #100;
A = 16'h00D2; B = 16'h0080; #100;
A = 16'h00D2; B = 16'h0081; #100;
A = 16'h00D2; B = 16'h0082; #100;
A = 16'h00D2; B = 16'h0083; #100;
A = 16'h00D2; B = 16'h0084; #100;
A = 16'h00D2; B = 16'h0085; #100;
A = 16'h00D2; B = 16'h0086; #100;
A = 16'h00D2; B = 16'h0087; #100;
A = 16'h00D2; B = 16'h0088; #100;
A = 16'h00D2; B = 16'h0089; #100;
A = 16'h00D2; B = 16'h008A; #100;
A = 16'h00D2; B = 16'h008B; #100;
A = 16'h00D2; B = 16'h008C; #100;
A = 16'h00D2; B = 16'h008D; #100;
A = 16'h00D2; B = 16'h008E; #100;
A = 16'h00D2; B = 16'h008F; #100;
A = 16'h00D2; B = 16'h0090; #100;
A = 16'h00D2; B = 16'h0091; #100;
A = 16'h00D2; B = 16'h0092; #100;
A = 16'h00D2; B = 16'h0093; #100;
A = 16'h00D2; B = 16'h0094; #100;
A = 16'h00D2; B = 16'h0095; #100;
A = 16'h00D2; B = 16'h0096; #100;
A = 16'h00D2; B = 16'h0097; #100;
A = 16'h00D2; B = 16'h0098; #100;
A = 16'h00D2; B = 16'h0099; #100;
A = 16'h00D2; B = 16'h009A; #100;
A = 16'h00D2; B = 16'h009B; #100;
A = 16'h00D2; B = 16'h009C; #100;
A = 16'h00D2; B = 16'h009D; #100;
A = 16'h00D2; B = 16'h009E; #100;
A = 16'h00D2; B = 16'h009F; #100;
A = 16'h00D2; B = 16'h00A0; #100;
A = 16'h00D2; B = 16'h00A1; #100;
A = 16'h00D2; B = 16'h00A2; #100;
A = 16'h00D2; B = 16'h00A3; #100;
A = 16'h00D2; B = 16'h00A4; #100;
A = 16'h00D2; B = 16'h00A5; #100;
A = 16'h00D2; B = 16'h00A6; #100;
A = 16'h00D2; B = 16'h00A7; #100;
A = 16'h00D2; B = 16'h00A8; #100;
A = 16'h00D2; B = 16'h00A9; #100;
A = 16'h00D2; B = 16'h00AA; #100;
A = 16'h00D2; B = 16'h00AB; #100;
A = 16'h00D2; B = 16'h00AC; #100;
A = 16'h00D2; B = 16'h00AD; #100;
A = 16'h00D2; B = 16'h00AE; #100;
A = 16'h00D2; B = 16'h00AF; #100;
A = 16'h00D2; B = 16'h00B0; #100;
A = 16'h00D2; B = 16'h00B1; #100;
A = 16'h00D2; B = 16'h00B2; #100;
A = 16'h00D2; B = 16'h00B3; #100;
A = 16'h00D2; B = 16'h00B4; #100;
A = 16'h00D2; B = 16'h00B5; #100;
A = 16'h00D2; B = 16'h00B6; #100;
A = 16'h00D2; B = 16'h00B7; #100;
A = 16'h00D2; B = 16'h00B8; #100;
A = 16'h00D2; B = 16'h00B9; #100;
A = 16'h00D2; B = 16'h00BA; #100;
A = 16'h00D2; B = 16'h00BB; #100;
A = 16'h00D2; B = 16'h00BC; #100;
A = 16'h00D2; B = 16'h00BD; #100;
A = 16'h00D2; B = 16'h00BE; #100;
A = 16'h00D2; B = 16'h00BF; #100;
A = 16'h00D2; B = 16'h00C0; #100;
A = 16'h00D2; B = 16'h00C1; #100;
A = 16'h00D2; B = 16'h00C2; #100;
A = 16'h00D2; B = 16'h00C3; #100;
A = 16'h00D2; B = 16'h00C4; #100;
A = 16'h00D2; B = 16'h00C5; #100;
A = 16'h00D2; B = 16'h00C6; #100;
A = 16'h00D2; B = 16'h00C7; #100;
A = 16'h00D2; B = 16'h00C8; #100;
A = 16'h00D2; B = 16'h00C9; #100;
A = 16'h00D2; B = 16'h00CA; #100;
A = 16'h00D2; B = 16'h00CB; #100;
A = 16'h00D2; B = 16'h00CC; #100;
A = 16'h00D2; B = 16'h00CD; #100;
A = 16'h00D2; B = 16'h00CE; #100;
A = 16'h00D2; B = 16'h00CF; #100;
A = 16'h00D2; B = 16'h00D0; #100;
A = 16'h00D2; B = 16'h00D1; #100;
A = 16'h00D2; B = 16'h00D2; #100;
A = 16'h00D2; B = 16'h00D3; #100;
A = 16'h00D2; B = 16'h00D4; #100;
A = 16'h00D2; B = 16'h00D5; #100;
A = 16'h00D2; B = 16'h00D6; #100;
A = 16'h00D2; B = 16'h00D7; #100;
A = 16'h00D2; B = 16'h00D8; #100;
A = 16'h00D2; B = 16'h00D9; #100;
A = 16'h00D2; B = 16'h00DA; #100;
A = 16'h00D2; B = 16'h00DB; #100;
A = 16'h00D2; B = 16'h00DC; #100;
A = 16'h00D2; B = 16'h00DD; #100;
A = 16'h00D2; B = 16'h00DE; #100;
A = 16'h00D2; B = 16'h00DF; #100;
A = 16'h00D2; B = 16'h00E0; #100;
A = 16'h00D2; B = 16'h00E1; #100;
A = 16'h00D2; B = 16'h00E2; #100;
A = 16'h00D2; B = 16'h00E3; #100;
A = 16'h00D2; B = 16'h00E4; #100;
A = 16'h00D2; B = 16'h00E5; #100;
A = 16'h00D2; B = 16'h00E6; #100;
A = 16'h00D2; B = 16'h00E7; #100;
A = 16'h00D2; B = 16'h00E8; #100;
A = 16'h00D2; B = 16'h00E9; #100;
A = 16'h00D2; B = 16'h00EA; #100;
A = 16'h00D2; B = 16'h00EB; #100;
A = 16'h00D2; B = 16'h00EC; #100;
A = 16'h00D2; B = 16'h00ED; #100;
A = 16'h00D2; B = 16'h00EE; #100;
A = 16'h00D2; B = 16'h00EF; #100;
A = 16'h00D2; B = 16'h00F0; #100;
A = 16'h00D2; B = 16'h00F1; #100;
A = 16'h00D2; B = 16'h00F2; #100;
A = 16'h00D2; B = 16'h00F3; #100;
A = 16'h00D2; B = 16'h00F4; #100;
A = 16'h00D2; B = 16'h00F5; #100;
A = 16'h00D2; B = 16'h00F6; #100;
A = 16'h00D2; B = 16'h00F7; #100;
A = 16'h00D2; B = 16'h00F8; #100;
A = 16'h00D2; B = 16'h00F9; #100;
A = 16'h00D2; B = 16'h00FA; #100;
A = 16'h00D2; B = 16'h00FB; #100;
A = 16'h00D2; B = 16'h00FC; #100;
A = 16'h00D2; B = 16'h00FD; #100;
A = 16'h00D2; B = 16'h00FE; #100;
A = 16'h00D2; B = 16'h00FF; #100;
A = 16'h00D3; B = 16'h000; #100;
A = 16'h00D3; B = 16'h001; #100;
A = 16'h00D3; B = 16'h002; #100;
A = 16'h00D3; B = 16'h003; #100;
A = 16'h00D3; B = 16'h004; #100;
A = 16'h00D3; B = 16'h005; #100;
A = 16'h00D3; B = 16'h006; #100;
A = 16'h00D3; B = 16'h007; #100;
A = 16'h00D3; B = 16'h008; #100;
A = 16'h00D3; B = 16'h009; #100;
A = 16'h00D3; B = 16'h00A; #100;
A = 16'h00D3; B = 16'h00B; #100;
A = 16'h00D3; B = 16'h00C; #100;
A = 16'h00D3; B = 16'h00D; #100;
A = 16'h00D3; B = 16'h00E; #100;
A = 16'h00D3; B = 16'h00F; #100;
A = 16'h00D3; B = 16'h0010; #100;
A = 16'h00D3; B = 16'h0011; #100;
A = 16'h00D3; B = 16'h0012; #100;
A = 16'h00D3; B = 16'h0013; #100;
A = 16'h00D3; B = 16'h0014; #100;
A = 16'h00D3; B = 16'h0015; #100;
A = 16'h00D3; B = 16'h0016; #100;
A = 16'h00D3; B = 16'h0017; #100;
A = 16'h00D3; B = 16'h0018; #100;
A = 16'h00D3; B = 16'h0019; #100;
A = 16'h00D3; B = 16'h001A; #100;
A = 16'h00D3; B = 16'h001B; #100;
A = 16'h00D3; B = 16'h001C; #100;
A = 16'h00D3; B = 16'h001D; #100;
A = 16'h00D3; B = 16'h001E; #100;
A = 16'h00D3; B = 16'h001F; #100;
A = 16'h00D3; B = 16'h0020; #100;
A = 16'h00D3; B = 16'h0021; #100;
A = 16'h00D3; B = 16'h0022; #100;
A = 16'h00D3; B = 16'h0023; #100;
A = 16'h00D3; B = 16'h0024; #100;
A = 16'h00D3; B = 16'h0025; #100;
A = 16'h00D3; B = 16'h0026; #100;
A = 16'h00D3; B = 16'h0027; #100;
A = 16'h00D3; B = 16'h0028; #100;
A = 16'h00D3; B = 16'h0029; #100;
A = 16'h00D3; B = 16'h002A; #100;
A = 16'h00D3; B = 16'h002B; #100;
A = 16'h00D3; B = 16'h002C; #100;
A = 16'h00D3; B = 16'h002D; #100;
A = 16'h00D3; B = 16'h002E; #100;
A = 16'h00D3; B = 16'h002F; #100;
A = 16'h00D3; B = 16'h0030; #100;
A = 16'h00D3; B = 16'h0031; #100;
A = 16'h00D3; B = 16'h0032; #100;
A = 16'h00D3; B = 16'h0033; #100;
A = 16'h00D3; B = 16'h0034; #100;
A = 16'h00D3; B = 16'h0035; #100;
A = 16'h00D3; B = 16'h0036; #100;
A = 16'h00D3; B = 16'h0037; #100;
A = 16'h00D3; B = 16'h0038; #100;
A = 16'h00D3; B = 16'h0039; #100;
A = 16'h00D3; B = 16'h003A; #100;
A = 16'h00D3; B = 16'h003B; #100;
A = 16'h00D3; B = 16'h003C; #100;
A = 16'h00D3; B = 16'h003D; #100;
A = 16'h00D3; B = 16'h003E; #100;
A = 16'h00D3; B = 16'h003F; #100;
A = 16'h00D3; B = 16'h0040; #100;
A = 16'h00D3; B = 16'h0041; #100;
A = 16'h00D3; B = 16'h0042; #100;
A = 16'h00D3; B = 16'h0043; #100;
A = 16'h00D3; B = 16'h0044; #100;
A = 16'h00D3; B = 16'h0045; #100;
A = 16'h00D3; B = 16'h0046; #100;
A = 16'h00D3; B = 16'h0047; #100;
A = 16'h00D3; B = 16'h0048; #100;
A = 16'h00D3; B = 16'h0049; #100;
A = 16'h00D3; B = 16'h004A; #100;
A = 16'h00D3; B = 16'h004B; #100;
A = 16'h00D3; B = 16'h004C; #100;
A = 16'h00D3; B = 16'h004D; #100;
A = 16'h00D3; B = 16'h004E; #100;
A = 16'h00D3; B = 16'h004F; #100;
A = 16'h00D3; B = 16'h0050; #100;
A = 16'h00D3; B = 16'h0051; #100;
A = 16'h00D3; B = 16'h0052; #100;
A = 16'h00D3; B = 16'h0053; #100;
A = 16'h00D3; B = 16'h0054; #100;
A = 16'h00D3; B = 16'h0055; #100;
A = 16'h00D3; B = 16'h0056; #100;
A = 16'h00D3; B = 16'h0057; #100;
A = 16'h00D3; B = 16'h0058; #100;
A = 16'h00D3; B = 16'h0059; #100;
A = 16'h00D3; B = 16'h005A; #100;
A = 16'h00D3; B = 16'h005B; #100;
A = 16'h00D3; B = 16'h005C; #100;
A = 16'h00D3; B = 16'h005D; #100;
A = 16'h00D3; B = 16'h005E; #100;
A = 16'h00D3; B = 16'h005F; #100;
A = 16'h00D3; B = 16'h0060; #100;
A = 16'h00D3; B = 16'h0061; #100;
A = 16'h00D3; B = 16'h0062; #100;
A = 16'h00D3; B = 16'h0063; #100;
A = 16'h00D3; B = 16'h0064; #100;
A = 16'h00D3; B = 16'h0065; #100;
A = 16'h00D3; B = 16'h0066; #100;
A = 16'h00D3; B = 16'h0067; #100;
A = 16'h00D3; B = 16'h0068; #100;
A = 16'h00D3; B = 16'h0069; #100;
A = 16'h00D3; B = 16'h006A; #100;
A = 16'h00D3; B = 16'h006B; #100;
A = 16'h00D3; B = 16'h006C; #100;
A = 16'h00D3; B = 16'h006D; #100;
A = 16'h00D3; B = 16'h006E; #100;
A = 16'h00D3; B = 16'h006F; #100;
A = 16'h00D3; B = 16'h0070; #100;
A = 16'h00D3; B = 16'h0071; #100;
A = 16'h00D3; B = 16'h0072; #100;
A = 16'h00D3; B = 16'h0073; #100;
A = 16'h00D3; B = 16'h0074; #100;
A = 16'h00D3; B = 16'h0075; #100;
A = 16'h00D3; B = 16'h0076; #100;
A = 16'h00D3; B = 16'h0077; #100;
A = 16'h00D3; B = 16'h0078; #100;
A = 16'h00D3; B = 16'h0079; #100;
A = 16'h00D3; B = 16'h007A; #100;
A = 16'h00D3; B = 16'h007B; #100;
A = 16'h00D3; B = 16'h007C; #100;
A = 16'h00D3; B = 16'h007D; #100;
A = 16'h00D3; B = 16'h007E; #100;
A = 16'h00D3; B = 16'h007F; #100;
A = 16'h00D3; B = 16'h0080; #100;
A = 16'h00D3; B = 16'h0081; #100;
A = 16'h00D3; B = 16'h0082; #100;
A = 16'h00D3; B = 16'h0083; #100;
A = 16'h00D3; B = 16'h0084; #100;
A = 16'h00D3; B = 16'h0085; #100;
A = 16'h00D3; B = 16'h0086; #100;
A = 16'h00D3; B = 16'h0087; #100;
A = 16'h00D3; B = 16'h0088; #100;
A = 16'h00D3; B = 16'h0089; #100;
A = 16'h00D3; B = 16'h008A; #100;
A = 16'h00D3; B = 16'h008B; #100;
A = 16'h00D3; B = 16'h008C; #100;
A = 16'h00D3; B = 16'h008D; #100;
A = 16'h00D3; B = 16'h008E; #100;
A = 16'h00D3; B = 16'h008F; #100;
A = 16'h00D3; B = 16'h0090; #100;
A = 16'h00D3; B = 16'h0091; #100;
A = 16'h00D3; B = 16'h0092; #100;
A = 16'h00D3; B = 16'h0093; #100;
A = 16'h00D3; B = 16'h0094; #100;
A = 16'h00D3; B = 16'h0095; #100;
A = 16'h00D3; B = 16'h0096; #100;
A = 16'h00D3; B = 16'h0097; #100;
A = 16'h00D3; B = 16'h0098; #100;
A = 16'h00D3; B = 16'h0099; #100;
A = 16'h00D3; B = 16'h009A; #100;
A = 16'h00D3; B = 16'h009B; #100;
A = 16'h00D3; B = 16'h009C; #100;
A = 16'h00D3; B = 16'h009D; #100;
A = 16'h00D3; B = 16'h009E; #100;
A = 16'h00D3; B = 16'h009F; #100;
A = 16'h00D3; B = 16'h00A0; #100;
A = 16'h00D3; B = 16'h00A1; #100;
A = 16'h00D3; B = 16'h00A2; #100;
A = 16'h00D3; B = 16'h00A3; #100;
A = 16'h00D3; B = 16'h00A4; #100;
A = 16'h00D3; B = 16'h00A5; #100;
A = 16'h00D3; B = 16'h00A6; #100;
A = 16'h00D3; B = 16'h00A7; #100;
A = 16'h00D3; B = 16'h00A8; #100;
A = 16'h00D3; B = 16'h00A9; #100;
A = 16'h00D3; B = 16'h00AA; #100;
A = 16'h00D3; B = 16'h00AB; #100;
A = 16'h00D3; B = 16'h00AC; #100;
A = 16'h00D3; B = 16'h00AD; #100;
A = 16'h00D3; B = 16'h00AE; #100;
A = 16'h00D3; B = 16'h00AF; #100;
A = 16'h00D3; B = 16'h00B0; #100;
A = 16'h00D3; B = 16'h00B1; #100;
A = 16'h00D3; B = 16'h00B2; #100;
A = 16'h00D3; B = 16'h00B3; #100;
A = 16'h00D3; B = 16'h00B4; #100;
A = 16'h00D3; B = 16'h00B5; #100;
A = 16'h00D3; B = 16'h00B6; #100;
A = 16'h00D3; B = 16'h00B7; #100;
A = 16'h00D3; B = 16'h00B8; #100;
A = 16'h00D3; B = 16'h00B9; #100;
A = 16'h00D3; B = 16'h00BA; #100;
A = 16'h00D3; B = 16'h00BB; #100;
A = 16'h00D3; B = 16'h00BC; #100;
A = 16'h00D3; B = 16'h00BD; #100;
A = 16'h00D3; B = 16'h00BE; #100;
A = 16'h00D3; B = 16'h00BF; #100;
A = 16'h00D3; B = 16'h00C0; #100;
A = 16'h00D3; B = 16'h00C1; #100;
A = 16'h00D3; B = 16'h00C2; #100;
A = 16'h00D3; B = 16'h00C3; #100;
A = 16'h00D3; B = 16'h00C4; #100;
A = 16'h00D3; B = 16'h00C5; #100;
A = 16'h00D3; B = 16'h00C6; #100;
A = 16'h00D3; B = 16'h00C7; #100;
A = 16'h00D3; B = 16'h00C8; #100;
A = 16'h00D3; B = 16'h00C9; #100;
A = 16'h00D3; B = 16'h00CA; #100;
A = 16'h00D3; B = 16'h00CB; #100;
A = 16'h00D3; B = 16'h00CC; #100;
A = 16'h00D3; B = 16'h00CD; #100;
A = 16'h00D3; B = 16'h00CE; #100;
A = 16'h00D3; B = 16'h00CF; #100;
A = 16'h00D3; B = 16'h00D0; #100;
A = 16'h00D3; B = 16'h00D1; #100;
A = 16'h00D3; B = 16'h00D2; #100;
A = 16'h00D3; B = 16'h00D3; #100;
A = 16'h00D3; B = 16'h00D4; #100;
A = 16'h00D3; B = 16'h00D5; #100;
A = 16'h00D3; B = 16'h00D6; #100;
A = 16'h00D3; B = 16'h00D7; #100;
A = 16'h00D3; B = 16'h00D8; #100;
A = 16'h00D3; B = 16'h00D9; #100;
A = 16'h00D3; B = 16'h00DA; #100;
A = 16'h00D3; B = 16'h00DB; #100;
A = 16'h00D3; B = 16'h00DC; #100;
A = 16'h00D3; B = 16'h00DD; #100;
A = 16'h00D3; B = 16'h00DE; #100;
A = 16'h00D3; B = 16'h00DF; #100;
A = 16'h00D3; B = 16'h00E0; #100;
A = 16'h00D3; B = 16'h00E1; #100;
A = 16'h00D3; B = 16'h00E2; #100;
A = 16'h00D3; B = 16'h00E3; #100;
A = 16'h00D3; B = 16'h00E4; #100;
A = 16'h00D3; B = 16'h00E5; #100;
A = 16'h00D3; B = 16'h00E6; #100;
A = 16'h00D3; B = 16'h00E7; #100;
A = 16'h00D3; B = 16'h00E8; #100;
A = 16'h00D3; B = 16'h00E9; #100;
A = 16'h00D3; B = 16'h00EA; #100;
A = 16'h00D3; B = 16'h00EB; #100;
A = 16'h00D3; B = 16'h00EC; #100;
A = 16'h00D3; B = 16'h00ED; #100;
A = 16'h00D3; B = 16'h00EE; #100;
A = 16'h00D3; B = 16'h00EF; #100;
A = 16'h00D3; B = 16'h00F0; #100;
A = 16'h00D3; B = 16'h00F1; #100;
A = 16'h00D3; B = 16'h00F2; #100;
A = 16'h00D3; B = 16'h00F3; #100;
A = 16'h00D3; B = 16'h00F4; #100;
A = 16'h00D3; B = 16'h00F5; #100;
A = 16'h00D3; B = 16'h00F6; #100;
A = 16'h00D3; B = 16'h00F7; #100;
A = 16'h00D3; B = 16'h00F8; #100;
A = 16'h00D3; B = 16'h00F9; #100;
A = 16'h00D3; B = 16'h00FA; #100;
A = 16'h00D3; B = 16'h00FB; #100;
A = 16'h00D3; B = 16'h00FC; #100;
A = 16'h00D3; B = 16'h00FD; #100;
A = 16'h00D3; B = 16'h00FE; #100;
A = 16'h00D3; B = 16'h00FF; #100;
A = 16'h00D4; B = 16'h000; #100;
A = 16'h00D4; B = 16'h001; #100;
A = 16'h00D4; B = 16'h002; #100;
A = 16'h00D4; B = 16'h003; #100;
A = 16'h00D4; B = 16'h004; #100;
A = 16'h00D4; B = 16'h005; #100;
A = 16'h00D4; B = 16'h006; #100;
A = 16'h00D4; B = 16'h007; #100;
A = 16'h00D4; B = 16'h008; #100;
A = 16'h00D4; B = 16'h009; #100;
A = 16'h00D4; B = 16'h00A; #100;
A = 16'h00D4; B = 16'h00B; #100;
A = 16'h00D4; B = 16'h00C; #100;
A = 16'h00D4; B = 16'h00D; #100;
A = 16'h00D4; B = 16'h00E; #100;
A = 16'h00D4; B = 16'h00F; #100;
A = 16'h00D4; B = 16'h0010; #100;
A = 16'h00D4; B = 16'h0011; #100;
A = 16'h00D4; B = 16'h0012; #100;
A = 16'h00D4; B = 16'h0013; #100;
A = 16'h00D4; B = 16'h0014; #100;
A = 16'h00D4; B = 16'h0015; #100;
A = 16'h00D4; B = 16'h0016; #100;
A = 16'h00D4; B = 16'h0017; #100;
A = 16'h00D4; B = 16'h0018; #100;
A = 16'h00D4; B = 16'h0019; #100;
A = 16'h00D4; B = 16'h001A; #100;
A = 16'h00D4; B = 16'h001B; #100;
A = 16'h00D4; B = 16'h001C; #100;
A = 16'h00D4; B = 16'h001D; #100;
A = 16'h00D4; B = 16'h001E; #100;
A = 16'h00D4; B = 16'h001F; #100;
A = 16'h00D4; B = 16'h0020; #100;
A = 16'h00D4; B = 16'h0021; #100;
A = 16'h00D4; B = 16'h0022; #100;
A = 16'h00D4; B = 16'h0023; #100;
A = 16'h00D4; B = 16'h0024; #100;
A = 16'h00D4; B = 16'h0025; #100;
A = 16'h00D4; B = 16'h0026; #100;
A = 16'h00D4; B = 16'h0027; #100;
A = 16'h00D4; B = 16'h0028; #100;
A = 16'h00D4; B = 16'h0029; #100;
A = 16'h00D4; B = 16'h002A; #100;
A = 16'h00D4; B = 16'h002B; #100;
A = 16'h00D4; B = 16'h002C; #100;
A = 16'h00D4; B = 16'h002D; #100;
A = 16'h00D4; B = 16'h002E; #100;
A = 16'h00D4; B = 16'h002F; #100;
A = 16'h00D4; B = 16'h0030; #100;
A = 16'h00D4; B = 16'h0031; #100;
A = 16'h00D4; B = 16'h0032; #100;
A = 16'h00D4; B = 16'h0033; #100;
A = 16'h00D4; B = 16'h0034; #100;
A = 16'h00D4; B = 16'h0035; #100;
A = 16'h00D4; B = 16'h0036; #100;
A = 16'h00D4; B = 16'h0037; #100;
A = 16'h00D4; B = 16'h0038; #100;
A = 16'h00D4; B = 16'h0039; #100;
A = 16'h00D4; B = 16'h003A; #100;
A = 16'h00D4; B = 16'h003B; #100;
A = 16'h00D4; B = 16'h003C; #100;
A = 16'h00D4; B = 16'h003D; #100;
A = 16'h00D4; B = 16'h003E; #100;
A = 16'h00D4; B = 16'h003F; #100;
A = 16'h00D4; B = 16'h0040; #100;
A = 16'h00D4; B = 16'h0041; #100;
A = 16'h00D4; B = 16'h0042; #100;
A = 16'h00D4; B = 16'h0043; #100;
A = 16'h00D4; B = 16'h0044; #100;
A = 16'h00D4; B = 16'h0045; #100;
A = 16'h00D4; B = 16'h0046; #100;
A = 16'h00D4; B = 16'h0047; #100;
A = 16'h00D4; B = 16'h0048; #100;
A = 16'h00D4; B = 16'h0049; #100;
A = 16'h00D4; B = 16'h004A; #100;
A = 16'h00D4; B = 16'h004B; #100;
A = 16'h00D4; B = 16'h004C; #100;
A = 16'h00D4; B = 16'h004D; #100;
A = 16'h00D4; B = 16'h004E; #100;
A = 16'h00D4; B = 16'h004F; #100;
A = 16'h00D4; B = 16'h0050; #100;
A = 16'h00D4; B = 16'h0051; #100;
A = 16'h00D4; B = 16'h0052; #100;
A = 16'h00D4; B = 16'h0053; #100;
A = 16'h00D4; B = 16'h0054; #100;
A = 16'h00D4; B = 16'h0055; #100;
A = 16'h00D4; B = 16'h0056; #100;
A = 16'h00D4; B = 16'h0057; #100;
A = 16'h00D4; B = 16'h0058; #100;
A = 16'h00D4; B = 16'h0059; #100;
A = 16'h00D4; B = 16'h005A; #100;
A = 16'h00D4; B = 16'h005B; #100;
A = 16'h00D4; B = 16'h005C; #100;
A = 16'h00D4; B = 16'h005D; #100;
A = 16'h00D4; B = 16'h005E; #100;
A = 16'h00D4; B = 16'h005F; #100;
A = 16'h00D4; B = 16'h0060; #100;
A = 16'h00D4; B = 16'h0061; #100;
A = 16'h00D4; B = 16'h0062; #100;
A = 16'h00D4; B = 16'h0063; #100;
A = 16'h00D4; B = 16'h0064; #100;
A = 16'h00D4; B = 16'h0065; #100;
A = 16'h00D4; B = 16'h0066; #100;
A = 16'h00D4; B = 16'h0067; #100;
A = 16'h00D4; B = 16'h0068; #100;
A = 16'h00D4; B = 16'h0069; #100;
A = 16'h00D4; B = 16'h006A; #100;
A = 16'h00D4; B = 16'h006B; #100;
A = 16'h00D4; B = 16'h006C; #100;
A = 16'h00D4; B = 16'h006D; #100;
A = 16'h00D4; B = 16'h006E; #100;
A = 16'h00D4; B = 16'h006F; #100;
A = 16'h00D4; B = 16'h0070; #100;
A = 16'h00D4; B = 16'h0071; #100;
A = 16'h00D4; B = 16'h0072; #100;
A = 16'h00D4; B = 16'h0073; #100;
A = 16'h00D4; B = 16'h0074; #100;
A = 16'h00D4; B = 16'h0075; #100;
A = 16'h00D4; B = 16'h0076; #100;
A = 16'h00D4; B = 16'h0077; #100;
A = 16'h00D4; B = 16'h0078; #100;
A = 16'h00D4; B = 16'h0079; #100;
A = 16'h00D4; B = 16'h007A; #100;
A = 16'h00D4; B = 16'h007B; #100;
A = 16'h00D4; B = 16'h007C; #100;
A = 16'h00D4; B = 16'h007D; #100;
A = 16'h00D4; B = 16'h007E; #100;
A = 16'h00D4; B = 16'h007F; #100;
A = 16'h00D4; B = 16'h0080; #100;
A = 16'h00D4; B = 16'h0081; #100;
A = 16'h00D4; B = 16'h0082; #100;
A = 16'h00D4; B = 16'h0083; #100;
A = 16'h00D4; B = 16'h0084; #100;
A = 16'h00D4; B = 16'h0085; #100;
A = 16'h00D4; B = 16'h0086; #100;
A = 16'h00D4; B = 16'h0087; #100;
A = 16'h00D4; B = 16'h0088; #100;
A = 16'h00D4; B = 16'h0089; #100;
A = 16'h00D4; B = 16'h008A; #100;
A = 16'h00D4; B = 16'h008B; #100;
A = 16'h00D4; B = 16'h008C; #100;
A = 16'h00D4; B = 16'h008D; #100;
A = 16'h00D4; B = 16'h008E; #100;
A = 16'h00D4; B = 16'h008F; #100;
A = 16'h00D4; B = 16'h0090; #100;
A = 16'h00D4; B = 16'h0091; #100;
A = 16'h00D4; B = 16'h0092; #100;
A = 16'h00D4; B = 16'h0093; #100;
A = 16'h00D4; B = 16'h0094; #100;
A = 16'h00D4; B = 16'h0095; #100;
A = 16'h00D4; B = 16'h0096; #100;
A = 16'h00D4; B = 16'h0097; #100;
A = 16'h00D4; B = 16'h0098; #100;
A = 16'h00D4; B = 16'h0099; #100;
A = 16'h00D4; B = 16'h009A; #100;
A = 16'h00D4; B = 16'h009B; #100;
A = 16'h00D4; B = 16'h009C; #100;
A = 16'h00D4; B = 16'h009D; #100;
A = 16'h00D4; B = 16'h009E; #100;
A = 16'h00D4; B = 16'h009F; #100;
A = 16'h00D4; B = 16'h00A0; #100;
A = 16'h00D4; B = 16'h00A1; #100;
A = 16'h00D4; B = 16'h00A2; #100;
A = 16'h00D4; B = 16'h00A3; #100;
A = 16'h00D4; B = 16'h00A4; #100;
A = 16'h00D4; B = 16'h00A5; #100;
A = 16'h00D4; B = 16'h00A6; #100;
A = 16'h00D4; B = 16'h00A7; #100;
A = 16'h00D4; B = 16'h00A8; #100;
A = 16'h00D4; B = 16'h00A9; #100;
A = 16'h00D4; B = 16'h00AA; #100;
A = 16'h00D4; B = 16'h00AB; #100;
A = 16'h00D4; B = 16'h00AC; #100;
A = 16'h00D4; B = 16'h00AD; #100;
A = 16'h00D4; B = 16'h00AE; #100;
A = 16'h00D4; B = 16'h00AF; #100;
A = 16'h00D4; B = 16'h00B0; #100;
A = 16'h00D4; B = 16'h00B1; #100;
A = 16'h00D4; B = 16'h00B2; #100;
A = 16'h00D4; B = 16'h00B3; #100;
A = 16'h00D4; B = 16'h00B4; #100;
A = 16'h00D4; B = 16'h00B5; #100;
A = 16'h00D4; B = 16'h00B6; #100;
A = 16'h00D4; B = 16'h00B7; #100;
A = 16'h00D4; B = 16'h00B8; #100;
A = 16'h00D4; B = 16'h00B9; #100;
A = 16'h00D4; B = 16'h00BA; #100;
A = 16'h00D4; B = 16'h00BB; #100;
A = 16'h00D4; B = 16'h00BC; #100;
A = 16'h00D4; B = 16'h00BD; #100;
A = 16'h00D4; B = 16'h00BE; #100;
A = 16'h00D4; B = 16'h00BF; #100;
A = 16'h00D4; B = 16'h00C0; #100;
A = 16'h00D4; B = 16'h00C1; #100;
A = 16'h00D4; B = 16'h00C2; #100;
A = 16'h00D4; B = 16'h00C3; #100;
A = 16'h00D4; B = 16'h00C4; #100;
A = 16'h00D4; B = 16'h00C5; #100;
A = 16'h00D4; B = 16'h00C6; #100;
A = 16'h00D4; B = 16'h00C7; #100;
A = 16'h00D4; B = 16'h00C8; #100;
A = 16'h00D4; B = 16'h00C9; #100;
A = 16'h00D4; B = 16'h00CA; #100;
A = 16'h00D4; B = 16'h00CB; #100;
A = 16'h00D4; B = 16'h00CC; #100;
A = 16'h00D4; B = 16'h00CD; #100;
A = 16'h00D4; B = 16'h00CE; #100;
A = 16'h00D4; B = 16'h00CF; #100;
A = 16'h00D4; B = 16'h00D0; #100;
A = 16'h00D4; B = 16'h00D1; #100;
A = 16'h00D4; B = 16'h00D2; #100;
A = 16'h00D4; B = 16'h00D3; #100;
A = 16'h00D4; B = 16'h00D4; #100;
A = 16'h00D4; B = 16'h00D5; #100;
A = 16'h00D4; B = 16'h00D6; #100;
A = 16'h00D4; B = 16'h00D7; #100;
A = 16'h00D4; B = 16'h00D8; #100;
A = 16'h00D4; B = 16'h00D9; #100;
A = 16'h00D4; B = 16'h00DA; #100;
A = 16'h00D4; B = 16'h00DB; #100;
A = 16'h00D4; B = 16'h00DC; #100;
A = 16'h00D4; B = 16'h00DD; #100;
A = 16'h00D4; B = 16'h00DE; #100;
A = 16'h00D4; B = 16'h00DF; #100;
A = 16'h00D4; B = 16'h00E0; #100;
A = 16'h00D4; B = 16'h00E1; #100;
A = 16'h00D4; B = 16'h00E2; #100;
A = 16'h00D4; B = 16'h00E3; #100;
A = 16'h00D4; B = 16'h00E4; #100;
A = 16'h00D4; B = 16'h00E5; #100;
A = 16'h00D4; B = 16'h00E6; #100;
A = 16'h00D4; B = 16'h00E7; #100;
A = 16'h00D4; B = 16'h00E8; #100;
A = 16'h00D4; B = 16'h00E9; #100;
A = 16'h00D4; B = 16'h00EA; #100;
A = 16'h00D4; B = 16'h00EB; #100;
A = 16'h00D4; B = 16'h00EC; #100;
A = 16'h00D4; B = 16'h00ED; #100;
A = 16'h00D4; B = 16'h00EE; #100;
A = 16'h00D4; B = 16'h00EF; #100;
A = 16'h00D4; B = 16'h00F0; #100;
A = 16'h00D4; B = 16'h00F1; #100;
A = 16'h00D4; B = 16'h00F2; #100;
A = 16'h00D4; B = 16'h00F3; #100;
A = 16'h00D4; B = 16'h00F4; #100;
A = 16'h00D4; B = 16'h00F5; #100;
A = 16'h00D4; B = 16'h00F6; #100;
A = 16'h00D4; B = 16'h00F7; #100;
A = 16'h00D4; B = 16'h00F8; #100;
A = 16'h00D4; B = 16'h00F9; #100;
A = 16'h00D4; B = 16'h00FA; #100;
A = 16'h00D4; B = 16'h00FB; #100;
A = 16'h00D4; B = 16'h00FC; #100;
A = 16'h00D4; B = 16'h00FD; #100;
A = 16'h00D4; B = 16'h00FE; #100;
A = 16'h00D4; B = 16'h00FF; #100;
A = 16'h00D5; B = 16'h000; #100;
A = 16'h00D5; B = 16'h001; #100;
A = 16'h00D5; B = 16'h002; #100;
A = 16'h00D5; B = 16'h003; #100;
A = 16'h00D5; B = 16'h004; #100;
A = 16'h00D5; B = 16'h005; #100;
A = 16'h00D5; B = 16'h006; #100;
A = 16'h00D5; B = 16'h007; #100;
A = 16'h00D5; B = 16'h008; #100;
A = 16'h00D5; B = 16'h009; #100;
A = 16'h00D5; B = 16'h00A; #100;
A = 16'h00D5; B = 16'h00B; #100;
A = 16'h00D5; B = 16'h00C; #100;
A = 16'h00D5; B = 16'h00D; #100;
A = 16'h00D5; B = 16'h00E; #100;
A = 16'h00D5; B = 16'h00F; #100;
A = 16'h00D5; B = 16'h0010; #100;
A = 16'h00D5; B = 16'h0011; #100;
A = 16'h00D5; B = 16'h0012; #100;
A = 16'h00D5; B = 16'h0013; #100;
A = 16'h00D5; B = 16'h0014; #100;
A = 16'h00D5; B = 16'h0015; #100;
A = 16'h00D5; B = 16'h0016; #100;
A = 16'h00D5; B = 16'h0017; #100;
A = 16'h00D5; B = 16'h0018; #100;
A = 16'h00D5; B = 16'h0019; #100;
A = 16'h00D5; B = 16'h001A; #100;
A = 16'h00D5; B = 16'h001B; #100;
A = 16'h00D5; B = 16'h001C; #100;
A = 16'h00D5; B = 16'h001D; #100;
A = 16'h00D5; B = 16'h001E; #100;
A = 16'h00D5; B = 16'h001F; #100;
A = 16'h00D5; B = 16'h0020; #100;
A = 16'h00D5; B = 16'h0021; #100;
A = 16'h00D5; B = 16'h0022; #100;
A = 16'h00D5; B = 16'h0023; #100;
A = 16'h00D5; B = 16'h0024; #100;
A = 16'h00D5; B = 16'h0025; #100;
A = 16'h00D5; B = 16'h0026; #100;
A = 16'h00D5; B = 16'h0027; #100;
A = 16'h00D5; B = 16'h0028; #100;
A = 16'h00D5; B = 16'h0029; #100;
A = 16'h00D5; B = 16'h002A; #100;
A = 16'h00D5; B = 16'h002B; #100;
A = 16'h00D5; B = 16'h002C; #100;
A = 16'h00D5; B = 16'h002D; #100;
A = 16'h00D5; B = 16'h002E; #100;
A = 16'h00D5; B = 16'h002F; #100;
A = 16'h00D5; B = 16'h0030; #100;
A = 16'h00D5; B = 16'h0031; #100;
A = 16'h00D5; B = 16'h0032; #100;
A = 16'h00D5; B = 16'h0033; #100;
A = 16'h00D5; B = 16'h0034; #100;
A = 16'h00D5; B = 16'h0035; #100;
A = 16'h00D5; B = 16'h0036; #100;
A = 16'h00D5; B = 16'h0037; #100;
A = 16'h00D5; B = 16'h0038; #100;
A = 16'h00D5; B = 16'h0039; #100;
A = 16'h00D5; B = 16'h003A; #100;
A = 16'h00D5; B = 16'h003B; #100;
A = 16'h00D5; B = 16'h003C; #100;
A = 16'h00D5; B = 16'h003D; #100;
A = 16'h00D5; B = 16'h003E; #100;
A = 16'h00D5; B = 16'h003F; #100;
A = 16'h00D5; B = 16'h0040; #100;
A = 16'h00D5; B = 16'h0041; #100;
A = 16'h00D5; B = 16'h0042; #100;
A = 16'h00D5; B = 16'h0043; #100;
A = 16'h00D5; B = 16'h0044; #100;
A = 16'h00D5; B = 16'h0045; #100;
A = 16'h00D5; B = 16'h0046; #100;
A = 16'h00D5; B = 16'h0047; #100;
A = 16'h00D5; B = 16'h0048; #100;
A = 16'h00D5; B = 16'h0049; #100;
A = 16'h00D5; B = 16'h004A; #100;
A = 16'h00D5; B = 16'h004B; #100;
A = 16'h00D5; B = 16'h004C; #100;
A = 16'h00D5; B = 16'h004D; #100;
A = 16'h00D5; B = 16'h004E; #100;
A = 16'h00D5; B = 16'h004F; #100;
A = 16'h00D5; B = 16'h0050; #100;
A = 16'h00D5; B = 16'h0051; #100;
A = 16'h00D5; B = 16'h0052; #100;
A = 16'h00D5; B = 16'h0053; #100;
A = 16'h00D5; B = 16'h0054; #100;
A = 16'h00D5; B = 16'h0055; #100;
A = 16'h00D5; B = 16'h0056; #100;
A = 16'h00D5; B = 16'h0057; #100;
A = 16'h00D5; B = 16'h0058; #100;
A = 16'h00D5; B = 16'h0059; #100;
A = 16'h00D5; B = 16'h005A; #100;
A = 16'h00D5; B = 16'h005B; #100;
A = 16'h00D5; B = 16'h005C; #100;
A = 16'h00D5; B = 16'h005D; #100;
A = 16'h00D5; B = 16'h005E; #100;
A = 16'h00D5; B = 16'h005F; #100;
A = 16'h00D5; B = 16'h0060; #100;
A = 16'h00D5; B = 16'h0061; #100;
A = 16'h00D5; B = 16'h0062; #100;
A = 16'h00D5; B = 16'h0063; #100;
A = 16'h00D5; B = 16'h0064; #100;
A = 16'h00D5; B = 16'h0065; #100;
A = 16'h00D5; B = 16'h0066; #100;
A = 16'h00D5; B = 16'h0067; #100;
A = 16'h00D5; B = 16'h0068; #100;
A = 16'h00D5; B = 16'h0069; #100;
A = 16'h00D5; B = 16'h006A; #100;
A = 16'h00D5; B = 16'h006B; #100;
A = 16'h00D5; B = 16'h006C; #100;
A = 16'h00D5; B = 16'h006D; #100;
A = 16'h00D5; B = 16'h006E; #100;
A = 16'h00D5; B = 16'h006F; #100;
A = 16'h00D5; B = 16'h0070; #100;
A = 16'h00D5; B = 16'h0071; #100;
A = 16'h00D5; B = 16'h0072; #100;
A = 16'h00D5; B = 16'h0073; #100;
A = 16'h00D5; B = 16'h0074; #100;
A = 16'h00D5; B = 16'h0075; #100;
A = 16'h00D5; B = 16'h0076; #100;
A = 16'h00D5; B = 16'h0077; #100;
A = 16'h00D5; B = 16'h0078; #100;
A = 16'h00D5; B = 16'h0079; #100;
A = 16'h00D5; B = 16'h007A; #100;
A = 16'h00D5; B = 16'h007B; #100;
A = 16'h00D5; B = 16'h007C; #100;
A = 16'h00D5; B = 16'h007D; #100;
A = 16'h00D5; B = 16'h007E; #100;
A = 16'h00D5; B = 16'h007F; #100;
A = 16'h00D5; B = 16'h0080; #100;
A = 16'h00D5; B = 16'h0081; #100;
A = 16'h00D5; B = 16'h0082; #100;
A = 16'h00D5; B = 16'h0083; #100;
A = 16'h00D5; B = 16'h0084; #100;
A = 16'h00D5; B = 16'h0085; #100;
A = 16'h00D5; B = 16'h0086; #100;
A = 16'h00D5; B = 16'h0087; #100;
A = 16'h00D5; B = 16'h0088; #100;
A = 16'h00D5; B = 16'h0089; #100;
A = 16'h00D5; B = 16'h008A; #100;
A = 16'h00D5; B = 16'h008B; #100;
A = 16'h00D5; B = 16'h008C; #100;
A = 16'h00D5; B = 16'h008D; #100;
A = 16'h00D5; B = 16'h008E; #100;
A = 16'h00D5; B = 16'h008F; #100;
A = 16'h00D5; B = 16'h0090; #100;
A = 16'h00D5; B = 16'h0091; #100;
A = 16'h00D5; B = 16'h0092; #100;
A = 16'h00D5; B = 16'h0093; #100;
A = 16'h00D5; B = 16'h0094; #100;
A = 16'h00D5; B = 16'h0095; #100;
A = 16'h00D5; B = 16'h0096; #100;
A = 16'h00D5; B = 16'h0097; #100;
A = 16'h00D5; B = 16'h0098; #100;
A = 16'h00D5; B = 16'h0099; #100;
A = 16'h00D5; B = 16'h009A; #100;
A = 16'h00D5; B = 16'h009B; #100;
A = 16'h00D5; B = 16'h009C; #100;
A = 16'h00D5; B = 16'h009D; #100;
A = 16'h00D5; B = 16'h009E; #100;
A = 16'h00D5; B = 16'h009F; #100;
A = 16'h00D5; B = 16'h00A0; #100;
A = 16'h00D5; B = 16'h00A1; #100;
A = 16'h00D5; B = 16'h00A2; #100;
A = 16'h00D5; B = 16'h00A3; #100;
A = 16'h00D5; B = 16'h00A4; #100;
A = 16'h00D5; B = 16'h00A5; #100;
A = 16'h00D5; B = 16'h00A6; #100;
A = 16'h00D5; B = 16'h00A7; #100;
A = 16'h00D5; B = 16'h00A8; #100;
A = 16'h00D5; B = 16'h00A9; #100;
A = 16'h00D5; B = 16'h00AA; #100;
A = 16'h00D5; B = 16'h00AB; #100;
A = 16'h00D5; B = 16'h00AC; #100;
A = 16'h00D5; B = 16'h00AD; #100;
A = 16'h00D5; B = 16'h00AE; #100;
A = 16'h00D5; B = 16'h00AF; #100;
A = 16'h00D5; B = 16'h00B0; #100;
A = 16'h00D5; B = 16'h00B1; #100;
A = 16'h00D5; B = 16'h00B2; #100;
A = 16'h00D5; B = 16'h00B3; #100;
A = 16'h00D5; B = 16'h00B4; #100;
A = 16'h00D5; B = 16'h00B5; #100;
A = 16'h00D5; B = 16'h00B6; #100;
A = 16'h00D5; B = 16'h00B7; #100;
A = 16'h00D5; B = 16'h00B8; #100;
A = 16'h00D5; B = 16'h00B9; #100;
A = 16'h00D5; B = 16'h00BA; #100;
A = 16'h00D5; B = 16'h00BB; #100;
A = 16'h00D5; B = 16'h00BC; #100;
A = 16'h00D5; B = 16'h00BD; #100;
A = 16'h00D5; B = 16'h00BE; #100;
A = 16'h00D5; B = 16'h00BF; #100;
A = 16'h00D5; B = 16'h00C0; #100;
A = 16'h00D5; B = 16'h00C1; #100;
A = 16'h00D5; B = 16'h00C2; #100;
A = 16'h00D5; B = 16'h00C3; #100;
A = 16'h00D5; B = 16'h00C4; #100;
A = 16'h00D5; B = 16'h00C5; #100;
A = 16'h00D5; B = 16'h00C6; #100;
A = 16'h00D5; B = 16'h00C7; #100;
A = 16'h00D5; B = 16'h00C8; #100;
A = 16'h00D5; B = 16'h00C9; #100;
A = 16'h00D5; B = 16'h00CA; #100;
A = 16'h00D5; B = 16'h00CB; #100;
A = 16'h00D5; B = 16'h00CC; #100;
A = 16'h00D5; B = 16'h00CD; #100;
A = 16'h00D5; B = 16'h00CE; #100;
A = 16'h00D5; B = 16'h00CF; #100;
A = 16'h00D5; B = 16'h00D0; #100;
A = 16'h00D5; B = 16'h00D1; #100;
A = 16'h00D5; B = 16'h00D2; #100;
A = 16'h00D5; B = 16'h00D3; #100;
A = 16'h00D5; B = 16'h00D4; #100;
A = 16'h00D5; B = 16'h00D5; #100;
A = 16'h00D5; B = 16'h00D6; #100;
A = 16'h00D5; B = 16'h00D7; #100;
A = 16'h00D5; B = 16'h00D8; #100;
A = 16'h00D5; B = 16'h00D9; #100;
A = 16'h00D5; B = 16'h00DA; #100;
A = 16'h00D5; B = 16'h00DB; #100;
A = 16'h00D5; B = 16'h00DC; #100;
A = 16'h00D5; B = 16'h00DD; #100;
A = 16'h00D5; B = 16'h00DE; #100;
A = 16'h00D5; B = 16'h00DF; #100;
A = 16'h00D5; B = 16'h00E0; #100;
A = 16'h00D5; B = 16'h00E1; #100;
A = 16'h00D5; B = 16'h00E2; #100;
A = 16'h00D5; B = 16'h00E3; #100;
A = 16'h00D5; B = 16'h00E4; #100;
A = 16'h00D5; B = 16'h00E5; #100;
A = 16'h00D5; B = 16'h00E6; #100;
A = 16'h00D5; B = 16'h00E7; #100;
A = 16'h00D5; B = 16'h00E8; #100;
A = 16'h00D5; B = 16'h00E9; #100;
A = 16'h00D5; B = 16'h00EA; #100;
A = 16'h00D5; B = 16'h00EB; #100;
A = 16'h00D5; B = 16'h00EC; #100;
A = 16'h00D5; B = 16'h00ED; #100;
A = 16'h00D5; B = 16'h00EE; #100;
A = 16'h00D5; B = 16'h00EF; #100;
A = 16'h00D5; B = 16'h00F0; #100;
A = 16'h00D5; B = 16'h00F1; #100;
A = 16'h00D5; B = 16'h00F2; #100;
A = 16'h00D5; B = 16'h00F3; #100;
A = 16'h00D5; B = 16'h00F4; #100;
A = 16'h00D5; B = 16'h00F5; #100;
A = 16'h00D5; B = 16'h00F6; #100;
A = 16'h00D5; B = 16'h00F7; #100;
A = 16'h00D5; B = 16'h00F8; #100;
A = 16'h00D5; B = 16'h00F9; #100;
A = 16'h00D5; B = 16'h00FA; #100;
A = 16'h00D5; B = 16'h00FB; #100;
A = 16'h00D5; B = 16'h00FC; #100;
A = 16'h00D5; B = 16'h00FD; #100;
A = 16'h00D5; B = 16'h00FE; #100;
A = 16'h00D5; B = 16'h00FF; #100;
A = 16'h00D6; B = 16'h000; #100;
A = 16'h00D6; B = 16'h001; #100;
A = 16'h00D6; B = 16'h002; #100;
A = 16'h00D6; B = 16'h003; #100;
A = 16'h00D6; B = 16'h004; #100;
A = 16'h00D6; B = 16'h005; #100;
A = 16'h00D6; B = 16'h006; #100;
A = 16'h00D6; B = 16'h007; #100;
A = 16'h00D6; B = 16'h008; #100;
A = 16'h00D6; B = 16'h009; #100;
A = 16'h00D6; B = 16'h00A; #100;
A = 16'h00D6; B = 16'h00B; #100;
A = 16'h00D6; B = 16'h00C; #100;
A = 16'h00D6; B = 16'h00D; #100;
A = 16'h00D6; B = 16'h00E; #100;
A = 16'h00D6; B = 16'h00F; #100;
A = 16'h00D6; B = 16'h0010; #100;
A = 16'h00D6; B = 16'h0011; #100;
A = 16'h00D6; B = 16'h0012; #100;
A = 16'h00D6; B = 16'h0013; #100;
A = 16'h00D6; B = 16'h0014; #100;
A = 16'h00D6; B = 16'h0015; #100;
A = 16'h00D6; B = 16'h0016; #100;
A = 16'h00D6; B = 16'h0017; #100;
A = 16'h00D6; B = 16'h0018; #100;
A = 16'h00D6; B = 16'h0019; #100;
A = 16'h00D6; B = 16'h001A; #100;
A = 16'h00D6; B = 16'h001B; #100;
A = 16'h00D6; B = 16'h001C; #100;
A = 16'h00D6; B = 16'h001D; #100;
A = 16'h00D6; B = 16'h001E; #100;
A = 16'h00D6; B = 16'h001F; #100;
A = 16'h00D6; B = 16'h0020; #100;
A = 16'h00D6; B = 16'h0021; #100;
A = 16'h00D6; B = 16'h0022; #100;
A = 16'h00D6; B = 16'h0023; #100;
A = 16'h00D6; B = 16'h0024; #100;
A = 16'h00D6; B = 16'h0025; #100;
A = 16'h00D6; B = 16'h0026; #100;
A = 16'h00D6; B = 16'h0027; #100;
A = 16'h00D6; B = 16'h0028; #100;
A = 16'h00D6; B = 16'h0029; #100;
A = 16'h00D6; B = 16'h002A; #100;
A = 16'h00D6; B = 16'h002B; #100;
A = 16'h00D6; B = 16'h002C; #100;
A = 16'h00D6; B = 16'h002D; #100;
A = 16'h00D6; B = 16'h002E; #100;
A = 16'h00D6; B = 16'h002F; #100;
A = 16'h00D6; B = 16'h0030; #100;
A = 16'h00D6; B = 16'h0031; #100;
A = 16'h00D6; B = 16'h0032; #100;
A = 16'h00D6; B = 16'h0033; #100;
A = 16'h00D6; B = 16'h0034; #100;
A = 16'h00D6; B = 16'h0035; #100;
A = 16'h00D6; B = 16'h0036; #100;
A = 16'h00D6; B = 16'h0037; #100;
A = 16'h00D6; B = 16'h0038; #100;
A = 16'h00D6; B = 16'h0039; #100;
A = 16'h00D6; B = 16'h003A; #100;
A = 16'h00D6; B = 16'h003B; #100;
A = 16'h00D6; B = 16'h003C; #100;
A = 16'h00D6; B = 16'h003D; #100;
A = 16'h00D6; B = 16'h003E; #100;
A = 16'h00D6; B = 16'h003F; #100;
A = 16'h00D6; B = 16'h0040; #100;
A = 16'h00D6; B = 16'h0041; #100;
A = 16'h00D6; B = 16'h0042; #100;
A = 16'h00D6; B = 16'h0043; #100;
A = 16'h00D6; B = 16'h0044; #100;
A = 16'h00D6; B = 16'h0045; #100;
A = 16'h00D6; B = 16'h0046; #100;
A = 16'h00D6; B = 16'h0047; #100;
A = 16'h00D6; B = 16'h0048; #100;
A = 16'h00D6; B = 16'h0049; #100;
A = 16'h00D6; B = 16'h004A; #100;
A = 16'h00D6; B = 16'h004B; #100;
A = 16'h00D6; B = 16'h004C; #100;
A = 16'h00D6; B = 16'h004D; #100;
A = 16'h00D6; B = 16'h004E; #100;
A = 16'h00D6; B = 16'h004F; #100;
A = 16'h00D6; B = 16'h0050; #100;
A = 16'h00D6; B = 16'h0051; #100;
A = 16'h00D6; B = 16'h0052; #100;
A = 16'h00D6; B = 16'h0053; #100;
A = 16'h00D6; B = 16'h0054; #100;
A = 16'h00D6; B = 16'h0055; #100;
A = 16'h00D6; B = 16'h0056; #100;
A = 16'h00D6; B = 16'h0057; #100;
A = 16'h00D6; B = 16'h0058; #100;
A = 16'h00D6; B = 16'h0059; #100;
A = 16'h00D6; B = 16'h005A; #100;
A = 16'h00D6; B = 16'h005B; #100;
A = 16'h00D6; B = 16'h005C; #100;
A = 16'h00D6; B = 16'h005D; #100;
A = 16'h00D6; B = 16'h005E; #100;
A = 16'h00D6; B = 16'h005F; #100;
A = 16'h00D6; B = 16'h0060; #100;
A = 16'h00D6; B = 16'h0061; #100;
A = 16'h00D6; B = 16'h0062; #100;
A = 16'h00D6; B = 16'h0063; #100;
A = 16'h00D6; B = 16'h0064; #100;
A = 16'h00D6; B = 16'h0065; #100;
A = 16'h00D6; B = 16'h0066; #100;
A = 16'h00D6; B = 16'h0067; #100;
A = 16'h00D6; B = 16'h0068; #100;
A = 16'h00D6; B = 16'h0069; #100;
A = 16'h00D6; B = 16'h006A; #100;
A = 16'h00D6; B = 16'h006B; #100;
A = 16'h00D6; B = 16'h006C; #100;
A = 16'h00D6; B = 16'h006D; #100;
A = 16'h00D6; B = 16'h006E; #100;
A = 16'h00D6; B = 16'h006F; #100;
A = 16'h00D6; B = 16'h0070; #100;
A = 16'h00D6; B = 16'h0071; #100;
A = 16'h00D6; B = 16'h0072; #100;
A = 16'h00D6; B = 16'h0073; #100;
A = 16'h00D6; B = 16'h0074; #100;
A = 16'h00D6; B = 16'h0075; #100;
A = 16'h00D6; B = 16'h0076; #100;
A = 16'h00D6; B = 16'h0077; #100;
A = 16'h00D6; B = 16'h0078; #100;
A = 16'h00D6; B = 16'h0079; #100;
A = 16'h00D6; B = 16'h007A; #100;
A = 16'h00D6; B = 16'h007B; #100;
A = 16'h00D6; B = 16'h007C; #100;
A = 16'h00D6; B = 16'h007D; #100;
A = 16'h00D6; B = 16'h007E; #100;
A = 16'h00D6; B = 16'h007F; #100;
A = 16'h00D6; B = 16'h0080; #100;
A = 16'h00D6; B = 16'h0081; #100;
A = 16'h00D6; B = 16'h0082; #100;
A = 16'h00D6; B = 16'h0083; #100;
A = 16'h00D6; B = 16'h0084; #100;
A = 16'h00D6; B = 16'h0085; #100;
A = 16'h00D6; B = 16'h0086; #100;
A = 16'h00D6; B = 16'h0087; #100;
A = 16'h00D6; B = 16'h0088; #100;
A = 16'h00D6; B = 16'h0089; #100;
A = 16'h00D6; B = 16'h008A; #100;
A = 16'h00D6; B = 16'h008B; #100;
A = 16'h00D6; B = 16'h008C; #100;
A = 16'h00D6; B = 16'h008D; #100;
A = 16'h00D6; B = 16'h008E; #100;
A = 16'h00D6; B = 16'h008F; #100;
A = 16'h00D6; B = 16'h0090; #100;
A = 16'h00D6; B = 16'h0091; #100;
A = 16'h00D6; B = 16'h0092; #100;
A = 16'h00D6; B = 16'h0093; #100;
A = 16'h00D6; B = 16'h0094; #100;
A = 16'h00D6; B = 16'h0095; #100;
A = 16'h00D6; B = 16'h0096; #100;
A = 16'h00D6; B = 16'h0097; #100;
A = 16'h00D6; B = 16'h0098; #100;
A = 16'h00D6; B = 16'h0099; #100;
A = 16'h00D6; B = 16'h009A; #100;
A = 16'h00D6; B = 16'h009B; #100;
A = 16'h00D6; B = 16'h009C; #100;
A = 16'h00D6; B = 16'h009D; #100;
A = 16'h00D6; B = 16'h009E; #100;
A = 16'h00D6; B = 16'h009F; #100;
A = 16'h00D6; B = 16'h00A0; #100;
A = 16'h00D6; B = 16'h00A1; #100;
A = 16'h00D6; B = 16'h00A2; #100;
A = 16'h00D6; B = 16'h00A3; #100;
A = 16'h00D6; B = 16'h00A4; #100;
A = 16'h00D6; B = 16'h00A5; #100;
A = 16'h00D6; B = 16'h00A6; #100;
A = 16'h00D6; B = 16'h00A7; #100;
A = 16'h00D6; B = 16'h00A8; #100;
A = 16'h00D6; B = 16'h00A9; #100;
A = 16'h00D6; B = 16'h00AA; #100;
A = 16'h00D6; B = 16'h00AB; #100;
A = 16'h00D6; B = 16'h00AC; #100;
A = 16'h00D6; B = 16'h00AD; #100;
A = 16'h00D6; B = 16'h00AE; #100;
A = 16'h00D6; B = 16'h00AF; #100;
A = 16'h00D6; B = 16'h00B0; #100;
A = 16'h00D6; B = 16'h00B1; #100;
A = 16'h00D6; B = 16'h00B2; #100;
A = 16'h00D6; B = 16'h00B3; #100;
A = 16'h00D6; B = 16'h00B4; #100;
A = 16'h00D6; B = 16'h00B5; #100;
A = 16'h00D6; B = 16'h00B6; #100;
A = 16'h00D6; B = 16'h00B7; #100;
A = 16'h00D6; B = 16'h00B8; #100;
A = 16'h00D6; B = 16'h00B9; #100;
A = 16'h00D6; B = 16'h00BA; #100;
A = 16'h00D6; B = 16'h00BB; #100;
A = 16'h00D6; B = 16'h00BC; #100;
A = 16'h00D6; B = 16'h00BD; #100;
A = 16'h00D6; B = 16'h00BE; #100;
A = 16'h00D6; B = 16'h00BF; #100;
A = 16'h00D6; B = 16'h00C0; #100;
A = 16'h00D6; B = 16'h00C1; #100;
A = 16'h00D6; B = 16'h00C2; #100;
A = 16'h00D6; B = 16'h00C3; #100;
A = 16'h00D6; B = 16'h00C4; #100;
A = 16'h00D6; B = 16'h00C5; #100;
A = 16'h00D6; B = 16'h00C6; #100;
A = 16'h00D6; B = 16'h00C7; #100;
A = 16'h00D6; B = 16'h00C8; #100;
A = 16'h00D6; B = 16'h00C9; #100;
A = 16'h00D6; B = 16'h00CA; #100;
A = 16'h00D6; B = 16'h00CB; #100;
A = 16'h00D6; B = 16'h00CC; #100;
A = 16'h00D6; B = 16'h00CD; #100;
A = 16'h00D6; B = 16'h00CE; #100;
A = 16'h00D6; B = 16'h00CF; #100;
A = 16'h00D6; B = 16'h00D0; #100;
A = 16'h00D6; B = 16'h00D1; #100;
A = 16'h00D6; B = 16'h00D2; #100;
A = 16'h00D6; B = 16'h00D3; #100;
A = 16'h00D6; B = 16'h00D4; #100;
A = 16'h00D6; B = 16'h00D5; #100;
A = 16'h00D6; B = 16'h00D6; #100;
A = 16'h00D6; B = 16'h00D7; #100;
A = 16'h00D6; B = 16'h00D8; #100;
A = 16'h00D6; B = 16'h00D9; #100;
A = 16'h00D6; B = 16'h00DA; #100;
A = 16'h00D6; B = 16'h00DB; #100;
A = 16'h00D6; B = 16'h00DC; #100;
A = 16'h00D6; B = 16'h00DD; #100;
A = 16'h00D6; B = 16'h00DE; #100;
A = 16'h00D6; B = 16'h00DF; #100;
A = 16'h00D6; B = 16'h00E0; #100;
A = 16'h00D6; B = 16'h00E1; #100;
A = 16'h00D6; B = 16'h00E2; #100;
A = 16'h00D6; B = 16'h00E3; #100;
A = 16'h00D6; B = 16'h00E4; #100;
A = 16'h00D6; B = 16'h00E5; #100;
A = 16'h00D6; B = 16'h00E6; #100;
A = 16'h00D6; B = 16'h00E7; #100;
A = 16'h00D6; B = 16'h00E8; #100;
A = 16'h00D6; B = 16'h00E9; #100;
A = 16'h00D6; B = 16'h00EA; #100;
A = 16'h00D6; B = 16'h00EB; #100;
A = 16'h00D6; B = 16'h00EC; #100;
A = 16'h00D6; B = 16'h00ED; #100;
A = 16'h00D6; B = 16'h00EE; #100;
A = 16'h00D6; B = 16'h00EF; #100;
A = 16'h00D6; B = 16'h00F0; #100;
A = 16'h00D6; B = 16'h00F1; #100;
A = 16'h00D6; B = 16'h00F2; #100;
A = 16'h00D6; B = 16'h00F3; #100;
A = 16'h00D6; B = 16'h00F4; #100;
A = 16'h00D6; B = 16'h00F5; #100;
A = 16'h00D6; B = 16'h00F6; #100;
A = 16'h00D6; B = 16'h00F7; #100;
A = 16'h00D6; B = 16'h00F8; #100;
A = 16'h00D6; B = 16'h00F9; #100;
A = 16'h00D6; B = 16'h00FA; #100;
A = 16'h00D6; B = 16'h00FB; #100;
A = 16'h00D6; B = 16'h00FC; #100;
A = 16'h00D6; B = 16'h00FD; #100;
A = 16'h00D6; B = 16'h00FE; #100;
A = 16'h00D6; B = 16'h00FF; #100;
A = 16'h00D7; B = 16'h000; #100;
A = 16'h00D7; B = 16'h001; #100;
A = 16'h00D7; B = 16'h002; #100;
A = 16'h00D7; B = 16'h003; #100;
A = 16'h00D7; B = 16'h004; #100;
A = 16'h00D7; B = 16'h005; #100;
A = 16'h00D7; B = 16'h006; #100;
A = 16'h00D7; B = 16'h007; #100;
A = 16'h00D7; B = 16'h008; #100;
A = 16'h00D7; B = 16'h009; #100;
A = 16'h00D7; B = 16'h00A; #100;
A = 16'h00D7; B = 16'h00B; #100;
A = 16'h00D7; B = 16'h00C; #100;
A = 16'h00D7; B = 16'h00D; #100;
A = 16'h00D7; B = 16'h00E; #100;
A = 16'h00D7; B = 16'h00F; #100;
A = 16'h00D7; B = 16'h0010; #100;
A = 16'h00D7; B = 16'h0011; #100;
A = 16'h00D7; B = 16'h0012; #100;
A = 16'h00D7; B = 16'h0013; #100;
A = 16'h00D7; B = 16'h0014; #100;
A = 16'h00D7; B = 16'h0015; #100;
A = 16'h00D7; B = 16'h0016; #100;
A = 16'h00D7; B = 16'h0017; #100;
A = 16'h00D7; B = 16'h0018; #100;
A = 16'h00D7; B = 16'h0019; #100;
A = 16'h00D7; B = 16'h001A; #100;
A = 16'h00D7; B = 16'h001B; #100;
A = 16'h00D7; B = 16'h001C; #100;
A = 16'h00D7; B = 16'h001D; #100;
A = 16'h00D7; B = 16'h001E; #100;
A = 16'h00D7; B = 16'h001F; #100;
A = 16'h00D7; B = 16'h0020; #100;
A = 16'h00D7; B = 16'h0021; #100;
A = 16'h00D7; B = 16'h0022; #100;
A = 16'h00D7; B = 16'h0023; #100;
A = 16'h00D7; B = 16'h0024; #100;
A = 16'h00D7; B = 16'h0025; #100;
A = 16'h00D7; B = 16'h0026; #100;
A = 16'h00D7; B = 16'h0027; #100;
A = 16'h00D7; B = 16'h0028; #100;
A = 16'h00D7; B = 16'h0029; #100;
A = 16'h00D7; B = 16'h002A; #100;
A = 16'h00D7; B = 16'h002B; #100;
A = 16'h00D7; B = 16'h002C; #100;
A = 16'h00D7; B = 16'h002D; #100;
A = 16'h00D7; B = 16'h002E; #100;
A = 16'h00D7; B = 16'h002F; #100;
A = 16'h00D7; B = 16'h0030; #100;
A = 16'h00D7; B = 16'h0031; #100;
A = 16'h00D7; B = 16'h0032; #100;
A = 16'h00D7; B = 16'h0033; #100;
A = 16'h00D7; B = 16'h0034; #100;
A = 16'h00D7; B = 16'h0035; #100;
A = 16'h00D7; B = 16'h0036; #100;
A = 16'h00D7; B = 16'h0037; #100;
A = 16'h00D7; B = 16'h0038; #100;
A = 16'h00D7; B = 16'h0039; #100;
A = 16'h00D7; B = 16'h003A; #100;
A = 16'h00D7; B = 16'h003B; #100;
A = 16'h00D7; B = 16'h003C; #100;
A = 16'h00D7; B = 16'h003D; #100;
A = 16'h00D7; B = 16'h003E; #100;
A = 16'h00D7; B = 16'h003F; #100;
A = 16'h00D7; B = 16'h0040; #100;
A = 16'h00D7; B = 16'h0041; #100;
A = 16'h00D7; B = 16'h0042; #100;
A = 16'h00D7; B = 16'h0043; #100;
A = 16'h00D7; B = 16'h0044; #100;
A = 16'h00D7; B = 16'h0045; #100;
A = 16'h00D7; B = 16'h0046; #100;
A = 16'h00D7; B = 16'h0047; #100;
A = 16'h00D7; B = 16'h0048; #100;
A = 16'h00D7; B = 16'h0049; #100;
A = 16'h00D7; B = 16'h004A; #100;
A = 16'h00D7; B = 16'h004B; #100;
A = 16'h00D7; B = 16'h004C; #100;
A = 16'h00D7; B = 16'h004D; #100;
A = 16'h00D7; B = 16'h004E; #100;
A = 16'h00D7; B = 16'h004F; #100;
A = 16'h00D7; B = 16'h0050; #100;
A = 16'h00D7; B = 16'h0051; #100;
A = 16'h00D7; B = 16'h0052; #100;
A = 16'h00D7; B = 16'h0053; #100;
A = 16'h00D7; B = 16'h0054; #100;
A = 16'h00D7; B = 16'h0055; #100;
A = 16'h00D7; B = 16'h0056; #100;
A = 16'h00D7; B = 16'h0057; #100;
A = 16'h00D7; B = 16'h0058; #100;
A = 16'h00D7; B = 16'h0059; #100;
A = 16'h00D7; B = 16'h005A; #100;
A = 16'h00D7; B = 16'h005B; #100;
A = 16'h00D7; B = 16'h005C; #100;
A = 16'h00D7; B = 16'h005D; #100;
A = 16'h00D7; B = 16'h005E; #100;
A = 16'h00D7; B = 16'h005F; #100;
A = 16'h00D7; B = 16'h0060; #100;
A = 16'h00D7; B = 16'h0061; #100;
A = 16'h00D7; B = 16'h0062; #100;
A = 16'h00D7; B = 16'h0063; #100;
A = 16'h00D7; B = 16'h0064; #100;
A = 16'h00D7; B = 16'h0065; #100;
A = 16'h00D7; B = 16'h0066; #100;
A = 16'h00D7; B = 16'h0067; #100;
A = 16'h00D7; B = 16'h0068; #100;
A = 16'h00D7; B = 16'h0069; #100;
A = 16'h00D7; B = 16'h006A; #100;
A = 16'h00D7; B = 16'h006B; #100;
A = 16'h00D7; B = 16'h006C; #100;
A = 16'h00D7; B = 16'h006D; #100;
A = 16'h00D7; B = 16'h006E; #100;
A = 16'h00D7; B = 16'h006F; #100;
A = 16'h00D7; B = 16'h0070; #100;
A = 16'h00D7; B = 16'h0071; #100;
A = 16'h00D7; B = 16'h0072; #100;
A = 16'h00D7; B = 16'h0073; #100;
A = 16'h00D7; B = 16'h0074; #100;
A = 16'h00D7; B = 16'h0075; #100;
A = 16'h00D7; B = 16'h0076; #100;
A = 16'h00D7; B = 16'h0077; #100;
A = 16'h00D7; B = 16'h0078; #100;
A = 16'h00D7; B = 16'h0079; #100;
A = 16'h00D7; B = 16'h007A; #100;
A = 16'h00D7; B = 16'h007B; #100;
A = 16'h00D7; B = 16'h007C; #100;
A = 16'h00D7; B = 16'h007D; #100;
A = 16'h00D7; B = 16'h007E; #100;
A = 16'h00D7; B = 16'h007F; #100;
A = 16'h00D7; B = 16'h0080; #100;
A = 16'h00D7; B = 16'h0081; #100;
A = 16'h00D7; B = 16'h0082; #100;
A = 16'h00D7; B = 16'h0083; #100;
A = 16'h00D7; B = 16'h0084; #100;
A = 16'h00D7; B = 16'h0085; #100;
A = 16'h00D7; B = 16'h0086; #100;
A = 16'h00D7; B = 16'h0087; #100;
A = 16'h00D7; B = 16'h0088; #100;
A = 16'h00D7; B = 16'h0089; #100;
A = 16'h00D7; B = 16'h008A; #100;
A = 16'h00D7; B = 16'h008B; #100;
A = 16'h00D7; B = 16'h008C; #100;
A = 16'h00D7; B = 16'h008D; #100;
A = 16'h00D7; B = 16'h008E; #100;
A = 16'h00D7; B = 16'h008F; #100;
A = 16'h00D7; B = 16'h0090; #100;
A = 16'h00D7; B = 16'h0091; #100;
A = 16'h00D7; B = 16'h0092; #100;
A = 16'h00D7; B = 16'h0093; #100;
A = 16'h00D7; B = 16'h0094; #100;
A = 16'h00D7; B = 16'h0095; #100;
A = 16'h00D7; B = 16'h0096; #100;
A = 16'h00D7; B = 16'h0097; #100;
A = 16'h00D7; B = 16'h0098; #100;
A = 16'h00D7; B = 16'h0099; #100;
A = 16'h00D7; B = 16'h009A; #100;
A = 16'h00D7; B = 16'h009B; #100;
A = 16'h00D7; B = 16'h009C; #100;
A = 16'h00D7; B = 16'h009D; #100;
A = 16'h00D7; B = 16'h009E; #100;
A = 16'h00D7; B = 16'h009F; #100;
A = 16'h00D7; B = 16'h00A0; #100;
A = 16'h00D7; B = 16'h00A1; #100;
A = 16'h00D7; B = 16'h00A2; #100;
A = 16'h00D7; B = 16'h00A3; #100;
A = 16'h00D7; B = 16'h00A4; #100;
A = 16'h00D7; B = 16'h00A5; #100;
A = 16'h00D7; B = 16'h00A6; #100;
A = 16'h00D7; B = 16'h00A7; #100;
A = 16'h00D7; B = 16'h00A8; #100;
A = 16'h00D7; B = 16'h00A9; #100;
A = 16'h00D7; B = 16'h00AA; #100;
A = 16'h00D7; B = 16'h00AB; #100;
A = 16'h00D7; B = 16'h00AC; #100;
A = 16'h00D7; B = 16'h00AD; #100;
A = 16'h00D7; B = 16'h00AE; #100;
A = 16'h00D7; B = 16'h00AF; #100;
A = 16'h00D7; B = 16'h00B0; #100;
A = 16'h00D7; B = 16'h00B1; #100;
A = 16'h00D7; B = 16'h00B2; #100;
A = 16'h00D7; B = 16'h00B3; #100;
A = 16'h00D7; B = 16'h00B4; #100;
A = 16'h00D7; B = 16'h00B5; #100;
A = 16'h00D7; B = 16'h00B6; #100;
A = 16'h00D7; B = 16'h00B7; #100;
A = 16'h00D7; B = 16'h00B8; #100;
A = 16'h00D7; B = 16'h00B9; #100;
A = 16'h00D7; B = 16'h00BA; #100;
A = 16'h00D7; B = 16'h00BB; #100;
A = 16'h00D7; B = 16'h00BC; #100;
A = 16'h00D7; B = 16'h00BD; #100;
A = 16'h00D7; B = 16'h00BE; #100;
A = 16'h00D7; B = 16'h00BF; #100;
A = 16'h00D7; B = 16'h00C0; #100;
A = 16'h00D7; B = 16'h00C1; #100;
A = 16'h00D7; B = 16'h00C2; #100;
A = 16'h00D7; B = 16'h00C3; #100;
A = 16'h00D7; B = 16'h00C4; #100;
A = 16'h00D7; B = 16'h00C5; #100;
A = 16'h00D7; B = 16'h00C6; #100;
A = 16'h00D7; B = 16'h00C7; #100;
A = 16'h00D7; B = 16'h00C8; #100;
A = 16'h00D7; B = 16'h00C9; #100;
A = 16'h00D7; B = 16'h00CA; #100;
A = 16'h00D7; B = 16'h00CB; #100;
A = 16'h00D7; B = 16'h00CC; #100;
A = 16'h00D7; B = 16'h00CD; #100;
A = 16'h00D7; B = 16'h00CE; #100;
A = 16'h00D7; B = 16'h00CF; #100;
A = 16'h00D7; B = 16'h00D0; #100;
A = 16'h00D7; B = 16'h00D1; #100;
A = 16'h00D7; B = 16'h00D2; #100;
A = 16'h00D7; B = 16'h00D3; #100;
A = 16'h00D7; B = 16'h00D4; #100;
A = 16'h00D7; B = 16'h00D5; #100;
A = 16'h00D7; B = 16'h00D6; #100;
A = 16'h00D7; B = 16'h00D7; #100;
A = 16'h00D7; B = 16'h00D8; #100;
A = 16'h00D7; B = 16'h00D9; #100;
A = 16'h00D7; B = 16'h00DA; #100;
A = 16'h00D7; B = 16'h00DB; #100;
A = 16'h00D7; B = 16'h00DC; #100;
A = 16'h00D7; B = 16'h00DD; #100;
A = 16'h00D7; B = 16'h00DE; #100;
A = 16'h00D7; B = 16'h00DF; #100;
A = 16'h00D7; B = 16'h00E0; #100;
A = 16'h00D7; B = 16'h00E1; #100;
A = 16'h00D7; B = 16'h00E2; #100;
A = 16'h00D7; B = 16'h00E3; #100;
A = 16'h00D7; B = 16'h00E4; #100;
A = 16'h00D7; B = 16'h00E5; #100;
A = 16'h00D7; B = 16'h00E6; #100;
A = 16'h00D7; B = 16'h00E7; #100;
A = 16'h00D7; B = 16'h00E8; #100;
A = 16'h00D7; B = 16'h00E9; #100;
A = 16'h00D7; B = 16'h00EA; #100;
A = 16'h00D7; B = 16'h00EB; #100;
A = 16'h00D7; B = 16'h00EC; #100;
A = 16'h00D7; B = 16'h00ED; #100;
A = 16'h00D7; B = 16'h00EE; #100;
A = 16'h00D7; B = 16'h00EF; #100;
A = 16'h00D7; B = 16'h00F0; #100;
A = 16'h00D7; B = 16'h00F1; #100;
A = 16'h00D7; B = 16'h00F2; #100;
A = 16'h00D7; B = 16'h00F3; #100;
A = 16'h00D7; B = 16'h00F4; #100;
A = 16'h00D7; B = 16'h00F5; #100;
A = 16'h00D7; B = 16'h00F6; #100;
A = 16'h00D7; B = 16'h00F7; #100;
A = 16'h00D7; B = 16'h00F8; #100;
A = 16'h00D7; B = 16'h00F9; #100;
A = 16'h00D7; B = 16'h00FA; #100;
A = 16'h00D7; B = 16'h00FB; #100;
A = 16'h00D7; B = 16'h00FC; #100;
A = 16'h00D7; B = 16'h00FD; #100;
A = 16'h00D7; B = 16'h00FE; #100;
A = 16'h00D7; B = 16'h00FF; #100;
A = 16'h00D8; B = 16'h000; #100;
A = 16'h00D8; B = 16'h001; #100;
A = 16'h00D8; B = 16'h002; #100;
A = 16'h00D8; B = 16'h003; #100;
A = 16'h00D8; B = 16'h004; #100;
A = 16'h00D8; B = 16'h005; #100;
A = 16'h00D8; B = 16'h006; #100;
A = 16'h00D8; B = 16'h007; #100;
A = 16'h00D8; B = 16'h008; #100;
A = 16'h00D8; B = 16'h009; #100;
A = 16'h00D8; B = 16'h00A; #100;
A = 16'h00D8; B = 16'h00B; #100;
A = 16'h00D8; B = 16'h00C; #100;
A = 16'h00D8; B = 16'h00D; #100;
A = 16'h00D8; B = 16'h00E; #100;
A = 16'h00D8; B = 16'h00F; #100;
A = 16'h00D8; B = 16'h0010; #100;
A = 16'h00D8; B = 16'h0011; #100;
A = 16'h00D8; B = 16'h0012; #100;
A = 16'h00D8; B = 16'h0013; #100;
A = 16'h00D8; B = 16'h0014; #100;
A = 16'h00D8; B = 16'h0015; #100;
A = 16'h00D8; B = 16'h0016; #100;
A = 16'h00D8; B = 16'h0017; #100;
A = 16'h00D8; B = 16'h0018; #100;
A = 16'h00D8; B = 16'h0019; #100;
A = 16'h00D8; B = 16'h001A; #100;
A = 16'h00D8; B = 16'h001B; #100;
A = 16'h00D8; B = 16'h001C; #100;
A = 16'h00D8; B = 16'h001D; #100;
A = 16'h00D8; B = 16'h001E; #100;
A = 16'h00D8; B = 16'h001F; #100;
A = 16'h00D8; B = 16'h0020; #100;
A = 16'h00D8; B = 16'h0021; #100;
A = 16'h00D8; B = 16'h0022; #100;
A = 16'h00D8; B = 16'h0023; #100;
A = 16'h00D8; B = 16'h0024; #100;
A = 16'h00D8; B = 16'h0025; #100;
A = 16'h00D8; B = 16'h0026; #100;
A = 16'h00D8; B = 16'h0027; #100;
A = 16'h00D8; B = 16'h0028; #100;
A = 16'h00D8; B = 16'h0029; #100;
A = 16'h00D8; B = 16'h002A; #100;
A = 16'h00D8; B = 16'h002B; #100;
A = 16'h00D8; B = 16'h002C; #100;
A = 16'h00D8; B = 16'h002D; #100;
A = 16'h00D8; B = 16'h002E; #100;
A = 16'h00D8; B = 16'h002F; #100;
A = 16'h00D8; B = 16'h0030; #100;
A = 16'h00D8; B = 16'h0031; #100;
A = 16'h00D8; B = 16'h0032; #100;
A = 16'h00D8; B = 16'h0033; #100;
A = 16'h00D8; B = 16'h0034; #100;
A = 16'h00D8; B = 16'h0035; #100;
A = 16'h00D8; B = 16'h0036; #100;
A = 16'h00D8; B = 16'h0037; #100;
A = 16'h00D8; B = 16'h0038; #100;
A = 16'h00D8; B = 16'h0039; #100;
A = 16'h00D8; B = 16'h003A; #100;
A = 16'h00D8; B = 16'h003B; #100;
A = 16'h00D8; B = 16'h003C; #100;
A = 16'h00D8; B = 16'h003D; #100;
A = 16'h00D8; B = 16'h003E; #100;
A = 16'h00D8; B = 16'h003F; #100;
A = 16'h00D8; B = 16'h0040; #100;
A = 16'h00D8; B = 16'h0041; #100;
A = 16'h00D8; B = 16'h0042; #100;
A = 16'h00D8; B = 16'h0043; #100;
A = 16'h00D8; B = 16'h0044; #100;
A = 16'h00D8; B = 16'h0045; #100;
A = 16'h00D8; B = 16'h0046; #100;
A = 16'h00D8; B = 16'h0047; #100;
A = 16'h00D8; B = 16'h0048; #100;
A = 16'h00D8; B = 16'h0049; #100;
A = 16'h00D8; B = 16'h004A; #100;
A = 16'h00D8; B = 16'h004B; #100;
A = 16'h00D8; B = 16'h004C; #100;
A = 16'h00D8; B = 16'h004D; #100;
A = 16'h00D8; B = 16'h004E; #100;
A = 16'h00D8; B = 16'h004F; #100;
A = 16'h00D8; B = 16'h0050; #100;
A = 16'h00D8; B = 16'h0051; #100;
A = 16'h00D8; B = 16'h0052; #100;
A = 16'h00D8; B = 16'h0053; #100;
A = 16'h00D8; B = 16'h0054; #100;
A = 16'h00D8; B = 16'h0055; #100;
A = 16'h00D8; B = 16'h0056; #100;
A = 16'h00D8; B = 16'h0057; #100;
A = 16'h00D8; B = 16'h0058; #100;
A = 16'h00D8; B = 16'h0059; #100;
A = 16'h00D8; B = 16'h005A; #100;
A = 16'h00D8; B = 16'h005B; #100;
A = 16'h00D8; B = 16'h005C; #100;
A = 16'h00D8; B = 16'h005D; #100;
A = 16'h00D8; B = 16'h005E; #100;
A = 16'h00D8; B = 16'h005F; #100;
A = 16'h00D8; B = 16'h0060; #100;
A = 16'h00D8; B = 16'h0061; #100;
A = 16'h00D8; B = 16'h0062; #100;
A = 16'h00D8; B = 16'h0063; #100;
A = 16'h00D8; B = 16'h0064; #100;
A = 16'h00D8; B = 16'h0065; #100;
A = 16'h00D8; B = 16'h0066; #100;
A = 16'h00D8; B = 16'h0067; #100;
A = 16'h00D8; B = 16'h0068; #100;
A = 16'h00D8; B = 16'h0069; #100;
A = 16'h00D8; B = 16'h006A; #100;
A = 16'h00D8; B = 16'h006B; #100;
A = 16'h00D8; B = 16'h006C; #100;
A = 16'h00D8; B = 16'h006D; #100;
A = 16'h00D8; B = 16'h006E; #100;
A = 16'h00D8; B = 16'h006F; #100;
A = 16'h00D8; B = 16'h0070; #100;
A = 16'h00D8; B = 16'h0071; #100;
A = 16'h00D8; B = 16'h0072; #100;
A = 16'h00D8; B = 16'h0073; #100;
A = 16'h00D8; B = 16'h0074; #100;
A = 16'h00D8; B = 16'h0075; #100;
A = 16'h00D8; B = 16'h0076; #100;
A = 16'h00D8; B = 16'h0077; #100;
A = 16'h00D8; B = 16'h0078; #100;
A = 16'h00D8; B = 16'h0079; #100;
A = 16'h00D8; B = 16'h007A; #100;
A = 16'h00D8; B = 16'h007B; #100;
A = 16'h00D8; B = 16'h007C; #100;
A = 16'h00D8; B = 16'h007D; #100;
A = 16'h00D8; B = 16'h007E; #100;
A = 16'h00D8; B = 16'h007F; #100;
A = 16'h00D8; B = 16'h0080; #100;
A = 16'h00D8; B = 16'h0081; #100;
A = 16'h00D8; B = 16'h0082; #100;
A = 16'h00D8; B = 16'h0083; #100;
A = 16'h00D8; B = 16'h0084; #100;
A = 16'h00D8; B = 16'h0085; #100;
A = 16'h00D8; B = 16'h0086; #100;
A = 16'h00D8; B = 16'h0087; #100;
A = 16'h00D8; B = 16'h0088; #100;
A = 16'h00D8; B = 16'h0089; #100;
A = 16'h00D8; B = 16'h008A; #100;
A = 16'h00D8; B = 16'h008B; #100;
A = 16'h00D8; B = 16'h008C; #100;
A = 16'h00D8; B = 16'h008D; #100;
A = 16'h00D8; B = 16'h008E; #100;
A = 16'h00D8; B = 16'h008F; #100;
A = 16'h00D8; B = 16'h0090; #100;
A = 16'h00D8; B = 16'h0091; #100;
A = 16'h00D8; B = 16'h0092; #100;
A = 16'h00D8; B = 16'h0093; #100;
A = 16'h00D8; B = 16'h0094; #100;
A = 16'h00D8; B = 16'h0095; #100;
A = 16'h00D8; B = 16'h0096; #100;
A = 16'h00D8; B = 16'h0097; #100;
A = 16'h00D8; B = 16'h0098; #100;
A = 16'h00D8; B = 16'h0099; #100;
A = 16'h00D8; B = 16'h009A; #100;
A = 16'h00D8; B = 16'h009B; #100;
A = 16'h00D8; B = 16'h009C; #100;
A = 16'h00D8; B = 16'h009D; #100;
A = 16'h00D8; B = 16'h009E; #100;
A = 16'h00D8; B = 16'h009F; #100;
A = 16'h00D8; B = 16'h00A0; #100;
A = 16'h00D8; B = 16'h00A1; #100;
A = 16'h00D8; B = 16'h00A2; #100;
A = 16'h00D8; B = 16'h00A3; #100;
A = 16'h00D8; B = 16'h00A4; #100;
A = 16'h00D8; B = 16'h00A5; #100;
A = 16'h00D8; B = 16'h00A6; #100;
A = 16'h00D8; B = 16'h00A7; #100;
A = 16'h00D8; B = 16'h00A8; #100;
A = 16'h00D8; B = 16'h00A9; #100;
A = 16'h00D8; B = 16'h00AA; #100;
A = 16'h00D8; B = 16'h00AB; #100;
A = 16'h00D8; B = 16'h00AC; #100;
A = 16'h00D8; B = 16'h00AD; #100;
A = 16'h00D8; B = 16'h00AE; #100;
A = 16'h00D8; B = 16'h00AF; #100;
A = 16'h00D8; B = 16'h00B0; #100;
A = 16'h00D8; B = 16'h00B1; #100;
A = 16'h00D8; B = 16'h00B2; #100;
A = 16'h00D8; B = 16'h00B3; #100;
A = 16'h00D8; B = 16'h00B4; #100;
A = 16'h00D8; B = 16'h00B5; #100;
A = 16'h00D8; B = 16'h00B6; #100;
A = 16'h00D8; B = 16'h00B7; #100;
A = 16'h00D8; B = 16'h00B8; #100;
A = 16'h00D8; B = 16'h00B9; #100;
A = 16'h00D8; B = 16'h00BA; #100;
A = 16'h00D8; B = 16'h00BB; #100;
A = 16'h00D8; B = 16'h00BC; #100;
A = 16'h00D8; B = 16'h00BD; #100;
A = 16'h00D8; B = 16'h00BE; #100;
A = 16'h00D8; B = 16'h00BF; #100;
A = 16'h00D8; B = 16'h00C0; #100;
A = 16'h00D8; B = 16'h00C1; #100;
A = 16'h00D8; B = 16'h00C2; #100;
A = 16'h00D8; B = 16'h00C3; #100;
A = 16'h00D8; B = 16'h00C4; #100;
A = 16'h00D8; B = 16'h00C5; #100;
A = 16'h00D8; B = 16'h00C6; #100;
A = 16'h00D8; B = 16'h00C7; #100;
A = 16'h00D8; B = 16'h00C8; #100;
A = 16'h00D8; B = 16'h00C9; #100;
A = 16'h00D8; B = 16'h00CA; #100;
A = 16'h00D8; B = 16'h00CB; #100;
A = 16'h00D8; B = 16'h00CC; #100;
A = 16'h00D8; B = 16'h00CD; #100;
A = 16'h00D8; B = 16'h00CE; #100;
A = 16'h00D8; B = 16'h00CF; #100;
A = 16'h00D8; B = 16'h00D0; #100;
A = 16'h00D8; B = 16'h00D1; #100;
A = 16'h00D8; B = 16'h00D2; #100;
A = 16'h00D8; B = 16'h00D3; #100;
A = 16'h00D8; B = 16'h00D4; #100;
A = 16'h00D8; B = 16'h00D5; #100;
A = 16'h00D8; B = 16'h00D6; #100;
A = 16'h00D8; B = 16'h00D7; #100;
A = 16'h00D8; B = 16'h00D8; #100;
A = 16'h00D8; B = 16'h00D9; #100;
A = 16'h00D8; B = 16'h00DA; #100;
A = 16'h00D8; B = 16'h00DB; #100;
A = 16'h00D8; B = 16'h00DC; #100;
A = 16'h00D8; B = 16'h00DD; #100;
A = 16'h00D8; B = 16'h00DE; #100;
A = 16'h00D8; B = 16'h00DF; #100;
A = 16'h00D8; B = 16'h00E0; #100;
A = 16'h00D8; B = 16'h00E1; #100;
A = 16'h00D8; B = 16'h00E2; #100;
A = 16'h00D8; B = 16'h00E3; #100;
A = 16'h00D8; B = 16'h00E4; #100;
A = 16'h00D8; B = 16'h00E5; #100;
A = 16'h00D8; B = 16'h00E6; #100;
A = 16'h00D8; B = 16'h00E7; #100;
A = 16'h00D8; B = 16'h00E8; #100;
A = 16'h00D8; B = 16'h00E9; #100;
A = 16'h00D8; B = 16'h00EA; #100;
A = 16'h00D8; B = 16'h00EB; #100;
A = 16'h00D8; B = 16'h00EC; #100;
A = 16'h00D8; B = 16'h00ED; #100;
A = 16'h00D8; B = 16'h00EE; #100;
A = 16'h00D8; B = 16'h00EF; #100;
A = 16'h00D8; B = 16'h00F0; #100;
A = 16'h00D8; B = 16'h00F1; #100;
A = 16'h00D8; B = 16'h00F2; #100;
A = 16'h00D8; B = 16'h00F3; #100;
A = 16'h00D8; B = 16'h00F4; #100;
A = 16'h00D8; B = 16'h00F5; #100;
A = 16'h00D8; B = 16'h00F6; #100;
A = 16'h00D8; B = 16'h00F7; #100;
A = 16'h00D8; B = 16'h00F8; #100;
A = 16'h00D8; B = 16'h00F9; #100;
A = 16'h00D8; B = 16'h00FA; #100;
A = 16'h00D8; B = 16'h00FB; #100;
A = 16'h00D8; B = 16'h00FC; #100;
A = 16'h00D8; B = 16'h00FD; #100;
A = 16'h00D8; B = 16'h00FE; #100;
A = 16'h00D8; B = 16'h00FF; #100;
A = 16'h00D9; B = 16'h000; #100;
A = 16'h00D9; B = 16'h001; #100;
A = 16'h00D9; B = 16'h002; #100;
A = 16'h00D9; B = 16'h003; #100;
A = 16'h00D9; B = 16'h004; #100;
A = 16'h00D9; B = 16'h005; #100;
A = 16'h00D9; B = 16'h006; #100;
A = 16'h00D9; B = 16'h007; #100;
A = 16'h00D9; B = 16'h008; #100;
A = 16'h00D9; B = 16'h009; #100;
A = 16'h00D9; B = 16'h00A; #100;
A = 16'h00D9; B = 16'h00B; #100;
A = 16'h00D9; B = 16'h00C; #100;
A = 16'h00D9; B = 16'h00D; #100;
A = 16'h00D9; B = 16'h00E; #100;
A = 16'h00D9; B = 16'h00F; #100;
A = 16'h00D9; B = 16'h0010; #100;
A = 16'h00D9; B = 16'h0011; #100;
A = 16'h00D9; B = 16'h0012; #100;
A = 16'h00D9; B = 16'h0013; #100;
A = 16'h00D9; B = 16'h0014; #100;
A = 16'h00D9; B = 16'h0015; #100;
A = 16'h00D9; B = 16'h0016; #100;
A = 16'h00D9; B = 16'h0017; #100;
A = 16'h00D9; B = 16'h0018; #100;
A = 16'h00D9; B = 16'h0019; #100;
A = 16'h00D9; B = 16'h001A; #100;
A = 16'h00D9; B = 16'h001B; #100;
A = 16'h00D9; B = 16'h001C; #100;
A = 16'h00D9; B = 16'h001D; #100;
A = 16'h00D9; B = 16'h001E; #100;
A = 16'h00D9; B = 16'h001F; #100;
A = 16'h00D9; B = 16'h0020; #100;
A = 16'h00D9; B = 16'h0021; #100;
A = 16'h00D9; B = 16'h0022; #100;
A = 16'h00D9; B = 16'h0023; #100;
A = 16'h00D9; B = 16'h0024; #100;
A = 16'h00D9; B = 16'h0025; #100;
A = 16'h00D9; B = 16'h0026; #100;
A = 16'h00D9; B = 16'h0027; #100;
A = 16'h00D9; B = 16'h0028; #100;
A = 16'h00D9; B = 16'h0029; #100;
A = 16'h00D9; B = 16'h002A; #100;
A = 16'h00D9; B = 16'h002B; #100;
A = 16'h00D9; B = 16'h002C; #100;
A = 16'h00D9; B = 16'h002D; #100;
A = 16'h00D9; B = 16'h002E; #100;
A = 16'h00D9; B = 16'h002F; #100;
A = 16'h00D9; B = 16'h0030; #100;
A = 16'h00D9; B = 16'h0031; #100;
A = 16'h00D9; B = 16'h0032; #100;
A = 16'h00D9; B = 16'h0033; #100;
A = 16'h00D9; B = 16'h0034; #100;
A = 16'h00D9; B = 16'h0035; #100;
A = 16'h00D9; B = 16'h0036; #100;
A = 16'h00D9; B = 16'h0037; #100;
A = 16'h00D9; B = 16'h0038; #100;
A = 16'h00D9; B = 16'h0039; #100;
A = 16'h00D9; B = 16'h003A; #100;
A = 16'h00D9; B = 16'h003B; #100;
A = 16'h00D9; B = 16'h003C; #100;
A = 16'h00D9; B = 16'h003D; #100;
A = 16'h00D9; B = 16'h003E; #100;
A = 16'h00D9; B = 16'h003F; #100;
A = 16'h00D9; B = 16'h0040; #100;
A = 16'h00D9; B = 16'h0041; #100;
A = 16'h00D9; B = 16'h0042; #100;
A = 16'h00D9; B = 16'h0043; #100;
A = 16'h00D9; B = 16'h0044; #100;
A = 16'h00D9; B = 16'h0045; #100;
A = 16'h00D9; B = 16'h0046; #100;
A = 16'h00D9; B = 16'h0047; #100;
A = 16'h00D9; B = 16'h0048; #100;
A = 16'h00D9; B = 16'h0049; #100;
A = 16'h00D9; B = 16'h004A; #100;
A = 16'h00D9; B = 16'h004B; #100;
A = 16'h00D9; B = 16'h004C; #100;
A = 16'h00D9; B = 16'h004D; #100;
A = 16'h00D9; B = 16'h004E; #100;
A = 16'h00D9; B = 16'h004F; #100;
A = 16'h00D9; B = 16'h0050; #100;
A = 16'h00D9; B = 16'h0051; #100;
A = 16'h00D9; B = 16'h0052; #100;
A = 16'h00D9; B = 16'h0053; #100;
A = 16'h00D9; B = 16'h0054; #100;
A = 16'h00D9; B = 16'h0055; #100;
A = 16'h00D9; B = 16'h0056; #100;
A = 16'h00D9; B = 16'h0057; #100;
A = 16'h00D9; B = 16'h0058; #100;
A = 16'h00D9; B = 16'h0059; #100;
A = 16'h00D9; B = 16'h005A; #100;
A = 16'h00D9; B = 16'h005B; #100;
A = 16'h00D9; B = 16'h005C; #100;
A = 16'h00D9; B = 16'h005D; #100;
A = 16'h00D9; B = 16'h005E; #100;
A = 16'h00D9; B = 16'h005F; #100;
A = 16'h00D9; B = 16'h0060; #100;
A = 16'h00D9; B = 16'h0061; #100;
A = 16'h00D9; B = 16'h0062; #100;
A = 16'h00D9; B = 16'h0063; #100;
A = 16'h00D9; B = 16'h0064; #100;
A = 16'h00D9; B = 16'h0065; #100;
A = 16'h00D9; B = 16'h0066; #100;
A = 16'h00D9; B = 16'h0067; #100;
A = 16'h00D9; B = 16'h0068; #100;
A = 16'h00D9; B = 16'h0069; #100;
A = 16'h00D9; B = 16'h006A; #100;
A = 16'h00D9; B = 16'h006B; #100;
A = 16'h00D9; B = 16'h006C; #100;
A = 16'h00D9; B = 16'h006D; #100;
A = 16'h00D9; B = 16'h006E; #100;
A = 16'h00D9; B = 16'h006F; #100;
A = 16'h00D9; B = 16'h0070; #100;
A = 16'h00D9; B = 16'h0071; #100;
A = 16'h00D9; B = 16'h0072; #100;
A = 16'h00D9; B = 16'h0073; #100;
A = 16'h00D9; B = 16'h0074; #100;
A = 16'h00D9; B = 16'h0075; #100;
A = 16'h00D9; B = 16'h0076; #100;
A = 16'h00D9; B = 16'h0077; #100;
A = 16'h00D9; B = 16'h0078; #100;
A = 16'h00D9; B = 16'h0079; #100;
A = 16'h00D9; B = 16'h007A; #100;
A = 16'h00D9; B = 16'h007B; #100;
A = 16'h00D9; B = 16'h007C; #100;
A = 16'h00D9; B = 16'h007D; #100;
A = 16'h00D9; B = 16'h007E; #100;
A = 16'h00D9; B = 16'h007F; #100;
A = 16'h00D9; B = 16'h0080; #100;
A = 16'h00D9; B = 16'h0081; #100;
A = 16'h00D9; B = 16'h0082; #100;
A = 16'h00D9; B = 16'h0083; #100;
A = 16'h00D9; B = 16'h0084; #100;
A = 16'h00D9; B = 16'h0085; #100;
A = 16'h00D9; B = 16'h0086; #100;
A = 16'h00D9; B = 16'h0087; #100;
A = 16'h00D9; B = 16'h0088; #100;
A = 16'h00D9; B = 16'h0089; #100;
A = 16'h00D9; B = 16'h008A; #100;
A = 16'h00D9; B = 16'h008B; #100;
A = 16'h00D9; B = 16'h008C; #100;
A = 16'h00D9; B = 16'h008D; #100;
A = 16'h00D9; B = 16'h008E; #100;
A = 16'h00D9; B = 16'h008F; #100;
A = 16'h00D9; B = 16'h0090; #100;
A = 16'h00D9; B = 16'h0091; #100;
A = 16'h00D9; B = 16'h0092; #100;
A = 16'h00D9; B = 16'h0093; #100;
A = 16'h00D9; B = 16'h0094; #100;
A = 16'h00D9; B = 16'h0095; #100;
A = 16'h00D9; B = 16'h0096; #100;
A = 16'h00D9; B = 16'h0097; #100;
A = 16'h00D9; B = 16'h0098; #100;
A = 16'h00D9; B = 16'h0099; #100;
A = 16'h00D9; B = 16'h009A; #100;
A = 16'h00D9; B = 16'h009B; #100;
A = 16'h00D9; B = 16'h009C; #100;
A = 16'h00D9; B = 16'h009D; #100;
A = 16'h00D9; B = 16'h009E; #100;
A = 16'h00D9; B = 16'h009F; #100;
A = 16'h00D9; B = 16'h00A0; #100;
A = 16'h00D9; B = 16'h00A1; #100;
A = 16'h00D9; B = 16'h00A2; #100;
A = 16'h00D9; B = 16'h00A3; #100;
A = 16'h00D9; B = 16'h00A4; #100;
A = 16'h00D9; B = 16'h00A5; #100;
A = 16'h00D9; B = 16'h00A6; #100;
A = 16'h00D9; B = 16'h00A7; #100;
A = 16'h00D9; B = 16'h00A8; #100;
A = 16'h00D9; B = 16'h00A9; #100;
A = 16'h00D9; B = 16'h00AA; #100;
A = 16'h00D9; B = 16'h00AB; #100;
A = 16'h00D9; B = 16'h00AC; #100;
A = 16'h00D9; B = 16'h00AD; #100;
A = 16'h00D9; B = 16'h00AE; #100;
A = 16'h00D9; B = 16'h00AF; #100;
A = 16'h00D9; B = 16'h00B0; #100;
A = 16'h00D9; B = 16'h00B1; #100;
A = 16'h00D9; B = 16'h00B2; #100;
A = 16'h00D9; B = 16'h00B3; #100;
A = 16'h00D9; B = 16'h00B4; #100;
A = 16'h00D9; B = 16'h00B5; #100;
A = 16'h00D9; B = 16'h00B6; #100;
A = 16'h00D9; B = 16'h00B7; #100;
A = 16'h00D9; B = 16'h00B8; #100;
A = 16'h00D9; B = 16'h00B9; #100;
A = 16'h00D9; B = 16'h00BA; #100;
A = 16'h00D9; B = 16'h00BB; #100;
A = 16'h00D9; B = 16'h00BC; #100;
A = 16'h00D9; B = 16'h00BD; #100;
A = 16'h00D9; B = 16'h00BE; #100;
A = 16'h00D9; B = 16'h00BF; #100;
A = 16'h00D9; B = 16'h00C0; #100;
A = 16'h00D9; B = 16'h00C1; #100;
A = 16'h00D9; B = 16'h00C2; #100;
A = 16'h00D9; B = 16'h00C3; #100;
A = 16'h00D9; B = 16'h00C4; #100;
A = 16'h00D9; B = 16'h00C5; #100;
A = 16'h00D9; B = 16'h00C6; #100;
A = 16'h00D9; B = 16'h00C7; #100;
A = 16'h00D9; B = 16'h00C8; #100;
A = 16'h00D9; B = 16'h00C9; #100;
A = 16'h00D9; B = 16'h00CA; #100;
A = 16'h00D9; B = 16'h00CB; #100;
A = 16'h00D9; B = 16'h00CC; #100;
A = 16'h00D9; B = 16'h00CD; #100;
A = 16'h00D9; B = 16'h00CE; #100;
A = 16'h00D9; B = 16'h00CF; #100;
A = 16'h00D9; B = 16'h00D0; #100;
A = 16'h00D9; B = 16'h00D1; #100;
A = 16'h00D9; B = 16'h00D2; #100;
A = 16'h00D9; B = 16'h00D3; #100;
A = 16'h00D9; B = 16'h00D4; #100;
A = 16'h00D9; B = 16'h00D5; #100;
A = 16'h00D9; B = 16'h00D6; #100;
A = 16'h00D9; B = 16'h00D7; #100;
A = 16'h00D9; B = 16'h00D8; #100;
A = 16'h00D9; B = 16'h00D9; #100;
A = 16'h00D9; B = 16'h00DA; #100;
A = 16'h00D9; B = 16'h00DB; #100;
A = 16'h00D9; B = 16'h00DC; #100;
A = 16'h00D9; B = 16'h00DD; #100;
A = 16'h00D9; B = 16'h00DE; #100;
A = 16'h00D9; B = 16'h00DF; #100;
A = 16'h00D9; B = 16'h00E0; #100;
A = 16'h00D9; B = 16'h00E1; #100;
A = 16'h00D9; B = 16'h00E2; #100;
A = 16'h00D9; B = 16'h00E3; #100;
A = 16'h00D9; B = 16'h00E4; #100;
A = 16'h00D9; B = 16'h00E5; #100;
A = 16'h00D9; B = 16'h00E6; #100;
A = 16'h00D9; B = 16'h00E7; #100;
A = 16'h00D9; B = 16'h00E8; #100;
A = 16'h00D9; B = 16'h00E9; #100;
A = 16'h00D9; B = 16'h00EA; #100;
A = 16'h00D9; B = 16'h00EB; #100;
A = 16'h00D9; B = 16'h00EC; #100;
A = 16'h00D9; B = 16'h00ED; #100;
A = 16'h00D9; B = 16'h00EE; #100;
A = 16'h00D9; B = 16'h00EF; #100;
A = 16'h00D9; B = 16'h00F0; #100;
A = 16'h00D9; B = 16'h00F1; #100;
A = 16'h00D9; B = 16'h00F2; #100;
A = 16'h00D9; B = 16'h00F3; #100;
A = 16'h00D9; B = 16'h00F4; #100;
A = 16'h00D9; B = 16'h00F5; #100;
A = 16'h00D9; B = 16'h00F6; #100;
A = 16'h00D9; B = 16'h00F7; #100;
A = 16'h00D9; B = 16'h00F8; #100;
A = 16'h00D9; B = 16'h00F9; #100;
A = 16'h00D9; B = 16'h00FA; #100;
A = 16'h00D9; B = 16'h00FB; #100;
A = 16'h00D9; B = 16'h00FC; #100;
A = 16'h00D9; B = 16'h00FD; #100;
A = 16'h00D9; B = 16'h00FE; #100;
A = 16'h00D9; B = 16'h00FF; #100;
A = 16'h00DA; B = 16'h000; #100;
A = 16'h00DA; B = 16'h001; #100;
A = 16'h00DA; B = 16'h002; #100;
A = 16'h00DA; B = 16'h003; #100;
A = 16'h00DA; B = 16'h004; #100;
A = 16'h00DA; B = 16'h005; #100;
A = 16'h00DA; B = 16'h006; #100;
A = 16'h00DA; B = 16'h007; #100;
A = 16'h00DA; B = 16'h008; #100;
A = 16'h00DA; B = 16'h009; #100;
A = 16'h00DA; B = 16'h00A; #100;
A = 16'h00DA; B = 16'h00B; #100;
A = 16'h00DA; B = 16'h00C; #100;
A = 16'h00DA; B = 16'h00D; #100;
A = 16'h00DA; B = 16'h00E; #100;
A = 16'h00DA; B = 16'h00F; #100;
A = 16'h00DA; B = 16'h0010; #100;
A = 16'h00DA; B = 16'h0011; #100;
A = 16'h00DA; B = 16'h0012; #100;
A = 16'h00DA; B = 16'h0013; #100;
A = 16'h00DA; B = 16'h0014; #100;
A = 16'h00DA; B = 16'h0015; #100;
A = 16'h00DA; B = 16'h0016; #100;
A = 16'h00DA; B = 16'h0017; #100;
A = 16'h00DA; B = 16'h0018; #100;
A = 16'h00DA; B = 16'h0019; #100;
A = 16'h00DA; B = 16'h001A; #100;
A = 16'h00DA; B = 16'h001B; #100;
A = 16'h00DA; B = 16'h001C; #100;
A = 16'h00DA; B = 16'h001D; #100;
A = 16'h00DA; B = 16'h001E; #100;
A = 16'h00DA; B = 16'h001F; #100;
A = 16'h00DA; B = 16'h0020; #100;
A = 16'h00DA; B = 16'h0021; #100;
A = 16'h00DA; B = 16'h0022; #100;
A = 16'h00DA; B = 16'h0023; #100;
A = 16'h00DA; B = 16'h0024; #100;
A = 16'h00DA; B = 16'h0025; #100;
A = 16'h00DA; B = 16'h0026; #100;
A = 16'h00DA; B = 16'h0027; #100;
A = 16'h00DA; B = 16'h0028; #100;
A = 16'h00DA; B = 16'h0029; #100;
A = 16'h00DA; B = 16'h002A; #100;
A = 16'h00DA; B = 16'h002B; #100;
A = 16'h00DA; B = 16'h002C; #100;
A = 16'h00DA; B = 16'h002D; #100;
A = 16'h00DA; B = 16'h002E; #100;
A = 16'h00DA; B = 16'h002F; #100;
A = 16'h00DA; B = 16'h0030; #100;
A = 16'h00DA; B = 16'h0031; #100;
A = 16'h00DA; B = 16'h0032; #100;
A = 16'h00DA; B = 16'h0033; #100;
A = 16'h00DA; B = 16'h0034; #100;
A = 16'h00DA; B = 16'h0035; #100;
A = 16'h00DA; B = 16'h0036; #100;
A = 16'h00DA; B = 16'h0037; #100;
A = 16'h00DA; B = 16'h0038; #100;
A = 16'h00DA; B = 16'h0039; #100;
A = 16'h00DA; B = 16'h003A; #100;
A = 16'h00DA; B = 16'h003B; #100;
A = 16'h00DA; B = 16'h003C; #100;
A = 16'h00DA; B = 16'h003D; #100;
A = 16'h00DA; B = 16'h003E; #100;
A = 16'h00DA; B = 16'h003F; #100;
A = 16'h00DA; B = 16'h0040; #100;
A = 16'h00DA; B = 16'h0041; #100;
A = 16'h00DA; B = 16'h0042; #100;
A = 16'h00DA; B = 16'h0043; #100;
A = 16'h00DA; B = 16'h0044; #100;
A = 16'h00DA; B = 16'h0045; #100;
A = 16'h00DA; B = 16'h0046; #100;
A = 16'h00DA; B = 16'h0047; #100;
A = 16'h00DA; B = 16'h0048; #100;
A = 16'h00DA; B = 16'h0049; #100;
A = 16'h00DA; B = 16'h004A; #100;
A = 16'h00DA; B = 16'h004B; #100;
A = 16'h00DA; B = 16'h004C; #100;
A = 16'h00DA; B = 16'h004D; #100;
A = 16'h00DA; B = 16'h004E; #100;
A = 16'h00DA; B = 16'h004F; #100;
A = 16'h00DA; B = 16'h0050; #100;
A = 16'h00DA; B = 16'h0051; #100;
A = 16'h00DA; B = 16'h0052; #100;
A = 16'h00DA; B = 16'h0053; #100;
A = 16'h00DA; B = 16'h0054; #100;
A = 16'h00DA; B = 16'h0055; #100;
A = 16'h00DA; B = 16'h0056; #100;
A = 16'h00DA; B = 16'h0057; #100;
A = 16'h00DA; B = 16'h0058; #100;
A = 16'h00DA; B = 16'h0059; #100;
A = 16'h00DA; B = 16'h005A; #100;
A = 16'h00DA; B = 16'h005B; #100;
A = 16'h00DA; B = 16'h005C; #100;
A = 16'h00DA; B = 16'h005D; #100;
A = 16'h00DA; B = 16'h005E; #100;
A = 16'h00DA; B = 16'h005F; #100;
A = 16'h00DA; B = 16'h0060; #100;
A = 16'h00DA; B = 16'h0061; #100;
A = 16'h00DA; B = 16'h0062; #100;
A = 16'h00DA; B = 16'h0063; #100;
A = 16'h00DA; B = 16'h0064; #100;
A = 16'h00DA; B = 16'h0065; #100;
A = 16'h00DA; B = 16'h0066; #100;
A = 16'h00DA; B = 16'h0067; #100;
A = 16'h00DA; B = 16'h0068; #100;
A = 16'h00DA; B = 16'h0069; #100;
A = 16'h00DA; B = 16'h006A; #100;
A = 16'h00DA; B = 16'h006B; #100;
A = 16'h00DA; B = 16'h006C; #100;
A = 16'h00DA; B = 16'h006D; #100;
A = 16'h00DA; B = 16'h006E; #100;
A = 16'h00DA; B = 16'h006F; #100;
A = 16'h00DA; B = 16'h0070; #100;
A = 16'h00DA; B = 16'h0071; #100;
A = 16'h00DA; B = 16'h0072; #100;
A = 16'h00DA; B = 16'h0073; #100;
A = 16'h00DA; B = 16'h0074; #100;
A = 16'h00DA; B = 16'h0075; #100;
A = 16'h00DA; B = 16'h0076; #100;
A = 16'h00DA; B = 16'h0077; #100;
A = 16'h00DA; B = 16'h0078; #100;
A = 16'h00DA; B = 16'h0079; #100;
A = 16'h00DA; B = 16'h007A; #100;
A = 16'h00DA; B = 16'h007B; #100;
A = 16'h00DA; B = 16'h007C; #100;
A = 16'h00DA; B = 16'h007D; #100;
A = 16'h00DA; B = 16'h007E; #100;
A = 16'h00DA; B = 16'h007F; #100;
A = 16'h00DA; B = 16'h0080; #100;
A = 16'h00DA; B = 16'h0081; #100;
A = 16'h00DA; B = 16'h0082; #100;
A = 16'h00DA; B = 16'h0083; #100;
A = 16'h00DA; B = 16'h0084; #100;
A = 16'h00DA; B = 16'h0085; #100;
A = 16'h00DA; B = 16'h0086; #100;
A = 16'h00DA; B = 16'h0087; #100;
A = 16'h00DA; B = 16'h0088; #100;
A = 16'h00DA; B = 16'h0089; #100;
A = 16'h00DA; B = 16'h008A; #100;
A = 16'h00DA; B = 16'h008B; #100;
A = 16'h00DA; B = 16'h008C; #100;
A = 16'h00DA; B = 16'h008D; #100;
A = 16'h00DA; B = 16'h008E; #100;
A = 16'h00DA; B = 16'h008F; #100;
A = 16'h00DA; B = 16'h0090; #100;
A = 16'h00DA; B = 16'h0091; #100;
A = 16'h00DA; B = 16'h0092; #100;
A = 16'h00DA; B = 16'h0093; #100;
A = 16'h00DA; B = 16'h0094; #100;
A = 16'h00DA; B = 16'h0095; #100;
A = 16'h00DA; B = 16'h0096; #100;
A = 16'h00DA; B = 16'h0097; #100;
A = 16'h00DA; B = 16'h0098; #100;
A = 16'h00DA; B = 16'h0099; #100;
A = 16'h00DA; B = 16'h009A; #100;
A = 16'h00DA; B = 16'h009B; #100;
A = 16'h00DA; B = 16'h009C; #100;
A = 16'h00DA; B = 16'h009D; #100;
A = 16'h00DA; B = 16'h009E; #100;
A = 16'h00DA; B = 16'h009F; #100;
A = 16'h00DA; B = 16'h00A0; #100;
A = 16'h00DA; B = 16'h00A1; #100;
A = 16'h00DA; B = 16'h00A2; #100;
A = 16'h00DA; B = 16'h00A3; #100;
A = 16'h00DA; B = 16'h00A4; #100;
A = 16'h00DA; B = 16'h00A5; #100;
A = 16'h00DA; B = 16'h00A6; #100;
A = 16'h00DA; B = 16'h00A7; #100;
A = 16'h00DA; B = 16'h00A8; #100;
A = 16'h00DA; B = 16'h00A9; #100;
A = 16'h00DA; B = 16'h00AA; #100;
A = 16'h00DA; B = 16'h00AB; #100;
A = 16'h00DA; B = 16'h00AC; #100;
A = 16'h00DA; B = 16'h00AD; #100;
A = 16'h00DA; B = 16'h00AE; #100;
A = 16'h00DA; B = 16'h00AF; #100;
A = 16'h00DA; B = 16'h00B0; #100;
A = 16'h00DA; B = 16'h00B1; #100;
A = 16'h00DA; B = 16'h00B2; #100;
A = 16'h00DA; B = 16'h00B3; #100;
A = 16'h00DA; B = 16'h00B4; #100;
A = 16'h00DA; B = 16'h00B5; #100;
A = 16'h00DA; B = 16'h00B6; #100;
A = 16'h00DA; B = 16'h00B7; #100;
A = 16'h00DA; B = 16'h00B8; #100;
A = 16'h00DA; B = 16'h00B9; #100;
A = 16'h00DA; B = 16'h00BA; #100;
A = 16'h00DA; B = 16'h00BB; #100;
A = 16'h00DA; B = 16'h00BC; #100;
A = 16'h00DA; B = 16'h00BD; #100;
A = 16'h00DA; B = 16'h00BE; #100;
A = 16'h00DA; B = 16'h00BF; #100;
A = 16'h00DA; B = 16'h00C0; #100;
A = 16'h00DA; B = 16'h00C1; #100;
A = 16'h00DA; B = 16'h00C2; #100;
A = 16'h00DA; B = 16'h00C3; #100;
A = 16'h00DA; B = 16'h00C4; #100;
A = 16'h00DA; B = 16'h00C5; #100;
A = 16'h00DA; B = 16'h00C6; #100;
A = 16'h00DA; B = 16'h00C7; #100;
A = 16'h00DA; B = 16'h00C8; #100;
A = 16'h00DA; B = 16'h00C9; #100;
A = 16'h00DA; B = 16'h00CA; #100;
A = 16'h00DA; B = 16'h00CB; #100;
A = 16'h00DA; B = 16'h00CC; #100;
A = 16'h00DA; B = 16'h00CD; #100;
A = 16'h00DA; B = 16'h00CE; #100;
A = 16'h00DA; B = 16'h00CF; #100;
A = 16'h00DA; B = 16'h00D0; #100;
A = 16'h00DA; B = 16'h00D1; #100;
A = 16'h00DA; B = 16'h00D2; #100;
A = 16'h00DA; B = 16'h00D3; #100;
A = 16'h00DA; B = 16'h00D4; #100;
A = 16'h00DA; B = 16'h00D5; #100;
A = 16'h00DA; B = 16'h00D6; #100;
A = 16'h00DA; B = 16'h00D7; #100;
A = 16'h00DA; B = 16'h00D8; #100;
A = 16'h00DA; B = 16'h00D9; #100;
A = 16'h00DA; B = 16'h00DA; #100;
A = 16'h00DA; B = 16'h00DB; #100;
A = 16'h00DA; B = 16'h00DC; #100;
A = 16'h00DA; B = 16'h00DD; #100;
A = 16'h00DA; B = 16'h00DE; #100;
A = 16'h00DA; B = 16'h00DF; #100;
A = 16'h00DA; B = 16'h00E0; #100;
A = 16'h00DA; B = 16'h00E1; #100;
A = 16'h00DA; B = 16'h00E2; #100;
A = 16'h00DA; B = 16'h00E3; #100;
A = 16'h00DA; B = 16'h00E4; #100;
A = 16'h00DA; B = 16'h00E5; #100;
A = 16'h00DA; B = 16'h00E6; #100;
A = 16'h00DA; B = 16'h00E7; #100;
A = 16'h00DA; B = 16'h00E8; #100;
A = 16'h00DA; B = 16'h00E9; #100;
A = 16'h00DA; B = 16'h00EA; #100;
A = 16'h00DA; B = 16'h00EB; #100;
A = 16'h00DA; B = 16'h00EC; #100;
A = 16'h00DA; B = 16'h00ED; #100;
A = 16'h00DA; B = 16'h00EE; #100;
A = 16'h00DA; B = 16'h00EF; #100;
A = 16'h00DA; B = 16'h00F0; #100;
A = 16'h00DA; B = 16'h00F1; #100;
A = 16'h00DA; B = 16'h00F2; #100;
A = 16'h00DA; B = 16'h00F3; #100;
A = 16'h00DA; B = 16'h00F4; #100;
A = 16'h00DA; B = 16'h00F5; #100;
A = 16'h00DA; B = 16'h00F6; #100;
A = 16'h00DA; B = 16'h00F7; #100;
A = 16'h00DA; B = 16'h00F8; #100;
A = 16'h00DA; B = 16'h00F9; #100;
A = 16'h00DA; B = 16'h00FA; #100;
A = 16'h00DA; B = 16'h00FB; #100;
A = 16'h00DA; B = 16'h00FC; #100;
A = 16'h00DA; B = 16'h00FD; #100;
A = 16'h00DA; B = 16'h00FE; #100;
A = 16'h00DA; B = 16'h00FF; #100;
A = 16'h00DB; B = 16'h000; #100;
A = 16'h00DB; B = 16'h001; #100;
A = 16'h00DB; B = 16'h002; #100;
A = 16'h00DB; B = 16'h003; #100;
A = 16'h00DB; B = 16'h004; #100;
A = 16'h00DB; B = 16'h005; #100;
A = 16'h00DB; B = 16'h006; #100;
A = 16'h00DB; B = 16'h007; #100;
A = 16'h00DB; B = 16'h008; #100;
A = 16'h00DB; B = 16'h009; #100;
A = 16'h00DB; B = 16'h00A; #100;
A = 16'h00DB; B = 16'h00B; #100;
A = 16'h00DB; B = 16'h00C; #100;
A = 16'h00DB; B = 16'h00D; #100;
A = 16'h00DB; B = 16'h00E; #100;
A = 16'h00DB; B = 16'h00F; #100;
A = 16'h00DB; B = 16'h0010; #100;
A = 16'h00DB; B = 16'h0011; #100;
A = 16'h00DB; B = 16'h0012; #100;
A = 16'h00DB; B = 16'h0013; #100;
A = 16'h00DB; B = 16'h0014; #100;
A = 16'h00DB; B = 16'h0015; #100;
A = 16'h00DB; B = 16'h0016; #100;
A = 16'h00DB; B = 16'h0017; #100;
A = 16'h00DB; B = 16'h0018; #100;
A = 16'h00DB; B = 16'h0019; #100;
A = 16'h00DB; B = 16'h001A; #100;
A = 16'h00DB; B = 16'h001B; #100;
A = 16'h00DB; B = 16'h001C; #100;
A = 16'h00DB; B = 16'h001D; #100;
A = 16'h00DB; B = 16'h001E; #100;
A = 16'h00DB; B = 16'h001F; #100;
A = 16'h00DB; B = 16'h0020; #100;
A = 16'h00DB; B = 16'h0021; #100;
A = 16'h00DB; B = 16'h0022; #100;
A = 16'h00DB; B = 16'h0023; #100;
A = 16'h00DB; B = 16'h0024; #100;
A = 16'h00DB; B = 16'h0025; #100;
A = 16'h00DB; B = 16'h0026; #100;
A = 16'h00DB; B = 16'h0027; #100;
A = 16'h00DB; B = 16'h0028; #100;
A = 16'h00DB; B = 16'h0029; #100;
A = 16'h00DB; B = 16'h002A; #100;
A = 16'h00DB; B = 16'h002B; #100;
A = 16'h00DB; B = 16'h002C; #100;
A = 16'h00DB; B = 16'h002D; #100;
A = 16'h00DB; B = 16'h002E; #100;
A = 16'h00DB; B = 16'h002F; #100;
A = 16'h00DB; B = 16'h0030; #100;
A = 16'h00DB; B = 16'h0031; #100;
A = 16'h00DB; B = 16'h0032; #100;
A = 16'h00DB; B = 16'h0033; #100;
A = 16'h00DB; B = 16'h0034; #100;
A = 16'h00DB; B = 16'h0035; #100;
A = 16'h00DB; B = 16'h0036; #100;
A = 16'h00DB; B = 16'h0037; #100;
A = 16'h00DB; B = 16'h0038; #100;
A = 16'h00DB; B = 16'h0039; #100;
A = 16'h00DB; B = 16'h003A; #100;
A = 16'h00DB; B = 16'h003B; #100;
A = 16'h00DB; B = 16'h003C; #100;
A = 16'h00DB; B = 16'h003D; #100;
A = 16'h00DB; B = 16'h003E; #100;
A = 16'h00DB; B = 16'h003F; #100;
A = 16'h00DB; B = 16'h0040; #100;
A = 16'h00DB; B = 16'h0041; #100;
A = 16'h00DB; B = 16'h0042; #100;
A = 16'h00DB; B = 16'h0043; #100;
A = 16'h00DB; B = 16'h0044; #100;
A = 16'h00DB; B = 16'h0045; #100;
A = 16'h00DB; B = 16'h0046; #100;
A = 16'h00DB; B = 16'h0047; #100;
A = 16'h00DB; B = 16'h0048; #100;
A = 16'h00DB; B = 16'h0049; #100;
A = 16'h00DB; B = 16'h004A; #100;
A = 16'h00DB; B = 16'h004B; #100;
A = 16'h00DB; B = 16'h004C; #100;
A = 16'h00DB; B = 16'h004D; #100;
A = 16'h00DB; B = 16'h004E; #100;
A = 16'h00DB; B = 16'h004F; #100;
A = 16'h00DB; B = 16'h0050; #100;
A = 16'h00DB; B = 16'h0051; #100;
A = 16'h00DB; B = 16'h0052; #100;
A = 16'h00DB; B = 16'h0053; #100;
A = 16'h00DB; B = 16'h0054; #100;
A = 16'h00DB; B = 16'h0055; #100;
A = 16'h00DB; B = 16'h0056; #100;
A = 16'h00DB; B = 16'h0057; #100;
A = 16'h00DB; B = 16'h0058; #100;
A = 16'h00DB; B = 16'h0059; #100;
A = 16'h00DB; B = 16'h005A; #100;
A = 16'h00DB; B = 16'h005B; #100;
A = 16'h00DB; B = 16'h005C; #100;
A = 16'h00DB; B = 16'h005D; #100;
A = 16'h00DB; B = 16'h005E; #100;
A = 16'h00DB; B = 16'h005F; #100;
A = 16'h00DB; B = 16'h0060; #100;
A = 16'h00DB; B = 16'h0061; #100;
A = 16'h00DB; B = 16'h0062; #100;
A = 16'h00DB; B = 16'h0063; #100;
A = 16'h00DB; B = 16'h0064; #100;
A = 16'h00DB; B = 16'h0065; #100;
A = 16'h00DB; B = 16'h0066; #100;
A = 16'h00DB; B = 16'h0067; #100;
A = 16'h00DB; B = 16'h0068; #100;
A = 16'h00DB; B = 16'h0069; #100;
A = 16'h00DB; B = 16'h006A; #100;
A = 16'h00DB; B = 16'h006B; #100;
A = 16'h00DB; B = 16'h006C; #100;
A = 16'h00DB; B = 16'h006D; #100;
A = 16'h00DB; B = 16'h006E; #100;
A = 16'h00DB; B = 16'h006F; #100;
A = 16'h00DB; B = 16'h0070; #100;
A = 16'h00DB; B = 16'h0071; #100;
A = 16'h00DB; B = 16'h0072; #100;
A = 16'h00DB; B = 16'h0073; #100;
A = 16'h00DB; B = 16'h0074; #100;
A = 16'h00DB; B = 16'h0075; #100;
A = 16'h00DB; B = 16'h0076; #100;
A = 16'h00DB; B = 16'h0077; #100;
A = 16'h00DB; B = 16'h0078; #100;
A = 16'h00DB; B = 16'h0079; #100;
A = 16'h00DB; B = 16'h007A; #100;
A = 16'h00DB; B = 16'h007B; #100;
A = 16'h00DB; B = 16'h007C; #100;
A = 16'h00DB; B = 16'h007D; #100;
A = 16'h00DB; B = 16'h007E; #100;
A = 16'h00DB; B = 16'h007F; #100;
A = 16'h00DB; B = 16'h0080; #100;
A = 16'h00DB; B = 16'h0081; #100;
A = 16'h00DB; B = 16'h0082; #100;
A = 16'h00DB; B = 16'h0083; #100;
A = 16'h00DB; B = 16'h0084; #100;
A = 16'h00DB; B = 16'h0085; #100;
A = 16'h00DB; B = 16'h0086; #100;
A = 16'h00DB; B = 16'h0087; #100;
A = 16'h00DB; B = 16'h0088; #100;
A = 16'h00DB; B = 16'h0089; #100;
A = 16'h00DB; B = 16'h008A; #100;
A = 16'h00DB; B = 16'h008B; #100;
A = 16'h00DB; B = 16'h008C; #100;
A = 16'h00DB; B = 16'h008D; #100;
A = 16'h00DB; B = 16'h008E; #100;
A = 16'h00DB; B = 16'h008F; #100;
A = 16'h00DB; B = 16'h0090; #100;
A = 16'h00DB; B = 16'h0091; #100;
A = 16'h00DB; B = 16'h0092; #100;
A = 16'h00DB; B = 16'h0093; #100;
A = 16'h00DB; B = 16'h0094; #100;
A = 16'h00DB; B = 16'h0095; #100;
A = 16'h00DB; B = 16'h0096; #100;
A = 16'h00DB; B = 16'h0097; #100;
A = 16'h00DB; B = 16'h0098; #100;
A = 16'h00DB; B = 16'h0099; #100;
A = 16'h00DB; B = 16'h009A; #100;
A = 16'h00DB; B = 16'h009B; #100;
A = 16'h00DB; B = 16'h009C; #100;
A = 16'h00DB; B = 16'h009D; #100;
A = 16'h00DB; B = 16'h009E; #100;
A = 16'h00DB; B = 16'h009F; #100;
A = 16'h00DB; B = 16'h00A0; #100;
A = 16'h00DB; B = 16'h00A1; #100;
A = 16'h00DB; B = 16'h00A2; #100;
A = 16'h00DB; B = 16'h00A3; #100;
A = 16'h00DB; B = 16'h00A4; #100;
A = 16'h00DB; B = 16'h00A5; #100;
A = 16'h00DB; B = 16'h00A6; #100;
A = 16'h00DB; B = 16'h00A7; #100;
A = 16'h00DB; B = 16'h00A8; #100;
A = 16'h00DB; B = 16'h00A9; #100;
A = 16'h00DB; B = 16'h00AA; #100;
A = 16'h00DB; B = 16'h00AB; #100;
A = 16'h00DB; B = 16'h00AC; #100;
A = 16'h00DB; B = 16'h00AD; #100;
A = 16'h00DB; B = 16'h00AE; #100;
A = 16'h00DB; B = 16'h00AF; #100;
A = 16'h00DB; B = 16'h00B0; #100;
A = 16'h00DB; B = 16'h00B1; #100;
A = 16'h00DB; B = 16'h00B2; #100;
A = 16'h00DB; B = 16'h00B3; #100;
A = 16'h00DB; B = 16'h00B4; #100;
A = 16'h00DB; B = 16'h00B5; #100;
A = 16'h00DB; B = 16'h00B6; #100;
A = 16'h00DB; B = 16'h00B7; #100;
A = 16'h00DB; B = 16'h00B8; #100;
A = 16'h00DB; B = 16'h00B9; #100;
A = 16'h00DB; B = 16'h00BA; #100;
A = 16'h00DB; B = 16'h00BB; #100;
A = 16'h00DB; B = 16'h00BC; #100;
A = 16'h00DB; B = 16'h00BD; #100;
A = 16'h00DB; B = 16'h00BE; #100;
A = 16'h00DB; B = 16'h00BF; #100;
A = 16'h00DB; B = 16'h00C0; #100;
A = 16'h00DB; B = 16'h00C1; #100;
A = 16'h00DB; B = 16'h00C2; #100;
A = 16'h00DB; B = 16'h00C3; #100;
A = 16'h00DB; B = 16'h00C4; #100;
A = 16'h00DB; B = 16'h00C5; #100;
A = 16'h00DB; B = 16'h00C6; #100;
A = 16'h00DB; B = 16'h00C7; #100;
A = 16'h00DB; B = 16'h00C8; #100;
A = 16'h00DB; B = 16'h00C9; #100;
A = 16'h00DB; B = 16'h00CA; #100;
A = 16'h00DB; B = 16'h00CB; #100;
A = 16'h00DB; B = 16'h00CC; #100;
A = 16'h00DB; B = 16'h00CD; #100;
A = 16'h00DB; B = 16'h00CE; #100;
A = 16'h00DB; B = 16'h00CF; #100;
A = 16'h00DB; B = 16'h00D0; #100;
A = 16'h00DB; B = 16'h00D1; #100;
A = 16'h00DB; B = 16'h00D2; #100;
A = 16'h00DB; B = 16'h00D3; #100;
A = 16'h00DB; B = 16'h00D4; #100;
A = 16'h00DB; B = 16'h00D5; #100;
A = 16'h00DB; B = 16'h00D6; #100;
A = 16'h00DB; B = 16'h00D7; #100;
A = 16'h00DB; B = 16'h00D8; #100;
A = 16'h00DB; B = 16'h00D9; #100;
A = 16'h00DB; B = 16'h00DA; #100;
A = 16'h00DB; B = 16'h00DB; #100;
A = 16'h00DB; B = 16'h00DC; #100;
A = 16'h00DB; B = 16'h00DD; #100;
A = 16'h00DB; B = 16'h00DE; #100;
A = 16'h00DB; B = 16'h00DF; #100;
A = 16'h00DB; B = 16'h00E0; #100;
A = 16'h00DB; B = 16'h00E1; #100;
A = 16'h00DB; B = 16'h00E2; #100;
A = 16'h00DB; B = 16'h00E3; #100;
A = 16'h00DB; B = 16'h00E4; #100;
A = 16'h00DB; B = 16'h00E5; #100;
A = 16'h00DB; B = 16'h00E6; #100;
A = 16'h00DB; B = 16'h00E7; #100;
A = 16'h00DB; B = 16'h00E8; #100;
A = 16'h00DB; B = 16'h00E9; #100;
A = 16'h00DB; B = 16'h00EA; #100;
A = 16'h00DB; B = 16'h00EB; #100;
A = 16'h00DB; B = 16'h00EC; #100;
A = 16'h00DB; B = 16'h00ED; #100;
A = 16'h00DB; B = 16'h00EE; #100;
A = 16'h00DB; B = 16'h00EF; #100;
A = 16'h00DB; B = 16'h00F0; #100;
A = 16'h00DB; B = 16'h00F1; #100;
A = 16'h00DB; B = 16'h00F2; #100;
A = 16'h00DB; B = 16'h00F3; #100;
A = 16'h00DB; B = 16'h00F4; #100;
A = 16'h00DB; B = 16'h00F5; #100;
A = 16'h00DB; B = 16'h00F6; #100;
A = 16'h00DB; B = 16'h00F7; #100;
A = 16'h00DB; B = 16'h00F8; #100;
A = 16'h00DB; B = 16'h00F9; #100;
A = 16'h00DB; B = 16'h00FA; #100;
A = 16'h00DB; B = 16'h00FB; #100;
A = 16'h00DB; B = 16'h00FC; #100;
A = 16'h00DB; B = 16'h00FD; #100;
A = 16'h00DB; B = 16'h00FE; #100;
A = 16'h00DB; B = 16'h00FF; #100;
A = 16'h00DC; B = 16'h000; #100;
A = 16'h00DC; B = 16'h001; #100;
A = 16'h00DC; B = 16'h002; #100;
A = 16'h00DC; B = 16'h003; #100;
A = 16'h00DC; B = 16'h004; #100;
A = 16'h00DC; B = 16'h005; #100;
A = 16'h00DC; B = 16'h006; #100;
A = 16'h00DC; B = 16'h007; #100;
A = 16'h00DC; B = 16'h008; #100;
A = 16'h00DC; B = 16'h009; #100;
A = 16'h00DC; B = 16'h00A; #100;
A = 16'h00DC; B = 16'h00B; #100;
A = 16'h00DC; B = 16'h00C; #100;
A = 16'h00DC; B = 16'h00D; #100;
A = 16'h00DC; B = 16'h00E; #100;
A = 16'h00DC; B = 16'h00F; #100;
A = 16'h00DC; B = 16'h0010; #100;
A = 16'h00DC; B = 16'h0011; #100;
A = 16'h00DC; B = 16'h0012; #100;
A = 16'h00DC; B = 16'h0013; #100;
A = 16'h00DC; B = 16'h0014; #100;
A = 16'h00DC; B = 16'h0015; #100;
A = 16'h00DC; B = 16'h0016; #100;
A = 16'h00DC; B = 16'h0017; #100;
A = 16'h00DC; B = 16'h0018; #100;
A = 16'h00DC; B = 16'h0019; #100;
A = 16'h00DC; B = 16'h001A; #100;
A = 16'h00DC; B = 16'h001B; #100;
A = 16'h00DC; B = 16'h001C; #100;
A = 16'h00DC; B = 16'h001D; #100;
A = 16'h00DC; B = 16'h001E; #100;
A = 16'h00DC; B = 16'h001F; #100;
A = 16'h00DC; B = 16'h0020; #100;
A = 16'h00DC; B = 16'h0021; #100;
A = 16'h00DC; B = 16'h0022; #100;
A = 16'h00DC; B = 16'h0023; #100;
A = 16'h00DC; B = 16'h0024; #100;
A = 16'h00DC; B = 16'h0025; #100;
A = 16'h00DC; B = 16'h0026; #100;
A = 16'h00DC; B = 16'h0027; #100;
A = 16'h00DC; B = 16'h0028; #100;
A = 16'h00DC; B = 16'h0029; #100;
A = 16'h00DC; B = 16'h002A; #100;
A = 16'h00DC; B = 16'h002B; #100;
A = 16'h00DC; B = 16'h002C; #100;
A = 16'h00DC; B = 16'h002D; #100;
A = 16'h00DC; B = 16'h002E; #100;
A = 16'h00DC; B = 16'h002F; #100;
A = 16'h00DC; B = 16'h0030; #100;
A = 16'h00DC; B = 16'h0031; #100;
A = 16'h00DC; B = 16'h0032; #100;
A = 16'h00DC; B = 16'h0033; #100;
A = 16'h00DC; B = 16'h0034; #100;
A = 16'h00DC; B = 16'h0035; #100;
A = 16'h00DC; B = 16'h0036; #100;
A = 16'h00DC; B = 16'h0037; #100;
A = 16'h00DC; B = 16'h0038; #100;
A = 16'h00DC; B = 16'h0039; #100;
A = 16'h00DC; B = 16'h003A; #100;
A = 16'h00DC; B = 16'h003B; #100;
A = 16'h00DC; B = 16'h003C; #100;
A = 16'h00DC; B = 16'h003D; #100;
A = 16'h00DC; B = 16'h003E; #100;
A = 16'h00DC; B = 16'h003F; #100;
A = 16'h00DC; B = 16'h0040; #100;
A = 16'h00DC; B = 16'h0041; #100;
A = 16'h00DC; B = 16'h0042; #100;
A = 16'h00DC; B = 16'h0043; #100;
A = 16'h00DC; B = 16'h0044; #100;
A = 16'h00DC; B = 16'h0045; #100;
A = 16'h00DC; B = 16'h0046; #100;
A = 16'h00DC; B = 16'h0047; #100;
A = 16'h00DC; B = 16'h0048; #100;
A = 16'h00DC; B = 16'h0049; #100;
A = 16'h00DC; B = 16'h004A; #100;
A = 16'h00DC; B = 16'h004B; #100;
A = 16'h00DC; B = 16'h004C; #100;
A = 16'h00DC; B = 16'h004D; #100;
A = 16'h00DC; B = 16'h004E; #100;
A = 16'h00DC; B = 16'h004F; #100;
A = 16'h00DC; B = 16'h0050; #100;
A = 16'h00DC; B = 16'h0051; #100;
A = 16'h00DC; B = 16'h0052; #100;
A = 16'h00DC; B = 16'h0053; #100;
A = 16'h00DC; B = 16'h0054; #100;
A = 16'h00DC; B = 16'h0055; #100;
A = 16'h00DC; B = 16'h0056; #100;
A = 16'h00DC; B = 16'h0057; #100;
A = 16'h00DC; B = 16'h0058; #100;
A = 16'h00DC; B = 16'h0059; #100;
A = 16'h00DC; B = 16'h005A; #100;
A = 16'h00DC; B = 16'h005B; #100;
A = 16'h00DC; B = 16'h005C; #100;
A = 16'h00DC; B = 16'h005D; #100;
A = 16'h00DC; B = 16'h005E; #100;
A = 16'h00DC; B = 16'h005F; #100;
A = 16'h00DC; B = 16'h0060; #100;
A = 16'h00DC; B = 16'h0061; #100;
A = 16'h00DC; B = 16'h0062; #100;
A = 16'h00DC; B = 16'h0063; #100;
A = 16'h00DC; B = 16'h0064; #100;
A = 16'h00DC; B = 16'h0065; #100;
A = 16'h00DC; B = 16'h0066; #100;
A = 16'h00DC; B = 16'h0067; #100;
A = 16'h00DC; B = 16'h0068; #100;
A = 16'h00DC; B = 16'h0069; #100;
A = 16'h00DC; B = 16'h006A; #100;
A = 16'h00DC; B = 16'h006B; #100;
A = 16'h00DC; B = 16'h006C; #100;
A = 16'h00DC; B = 16'h006D; #100;
A = 16'h00DC; B = 16'h006E; #100;
A = 16'h00DC; B = 16'h006F; #100;
A = 16'h00DC; B = 16'h0070; #100;
A = 16'h00DC; B = 16'h0071; #100;
A = 16'h00DC; B = 16'h0072; #100;
A = 16'h00DC; B = 16'h0073; #100;
A = 16'h00DC; B = 16'h0074; #100;
A = 16'h00DC; B = 16'h0075; #100;
A = 16'h00DC; B = 16'h0076; #100;
A = 16'h00DC; B = 16'h0077; #100;
A = 16'h00DC; B = 16'h0078; #100;
A = 16'h00DC; B = 16'h0079; #100;
A = 16'h00DC; B = 16'h007A; #100;
A = 16'h00DC; B = 16'h007B; #100;
A = 16'h00DC; B = 16'h007C; #100;
A = 16'h00DC; B = 16'h007D; #100;
A = 16'h00DC; B = 16'h007E; #100;
A = 16'h00DC; B = 16'h007F; #100;
A = 16'h00DC; B = 16'h0080; #100;
A = 16'h00DC; B = 16'h0081; #100;
A = 16'h00DC; B = 16'h0082; #100;
A = 16'h00DC; B = 16'h0083; #100;
A = 16'h00DC; B = 16'h0084; #100;
A = 16'h00DC; B = 16'h0085; #100;
A = 16'h00DC; B = 16'h0086; #100;
A = 16'h00DC; B = 16'h0087; #100;
A = 16'h00DC; B = 16'h0088; #100;
A = 16'h00DC; B = 16'h0089; #100;
A = 16'h00DC; B = 16'h008A; #100;
A = 16'h00DC; B = 16'h008B; #100;
A = 16'h00DC; B = 16'h008C; #100;
A = 16'h00DC; B = 16'h008D; #100;
A = 16'h00DC; B = 16'h008E; #100;
A = 16'h00DC; B = 16'h008F; #100;
A = 16'h00DC; B = 16'h0090; #100;
A = 16'h00DC; B = 16'h0091; #100;
A = 16'h00DC; B = 16'h0092; #100;
A = 16'h00DC; B = 16'h0093; #100;
A = 16'h00DC; B = 16'h0094; #100;
A = 16'h00DC; B = 16'h0095; #100;
A = 16'h00DC; B = 16'h0096; #100;
A = 16'h00DC; B = 16'h0097; #100;
A = 16'h00DC; B = 16'h0098; #100;
A = 16'h00DC; B = 16'h0099; #100;
A = 16'h00DC; B = 16'h009A; #100;
A = 16'h00DC; B = 16'h009B; #100;
A = 16'h00DC; B = 16'h009C; #100;
A = 16'h00DC; B = 16'h009D; #100;
A = 16'h00DC; B = 16'h009E; #100;
A = 16'h00DC; B = 16'h009F; #100;
A = 16'h00DC; B = 16'h00A0; #100;
A = 16'h00DC; B = 16'h00A1; #100;
A = 16'h00DC; B = 16'h00A2; #100;
A = 16'h00DC; B = 16'h00A3; #100;
A = 16'h00DC; B = 16'h00A4; #100;
A = 16'h00DC; B = 16'h00A5; #100;
A = 16'h00DC; B = 16'h00A6; #100;
A = 16'h00DC; B = 16'h00A7; #100;
A = 16'h00DC; B = 16'h00A8; #100;
A = 16'h00DC; B = 16'h00A9; #100;
A = 16'h00DC; B = 16'h00AA; #100;
A = 16'h00DC; B = 16'h00AB; #100;
A = 16'h00DC; B = 16'h00AC; #100;
A = 16'h00DC; B = 16'h00AD; #100;
A = 16'h00DC; B = 16'h00AE; #100;
A = 16'h00DC; B = 16'h00AF; #100;
A = 16'h00DC; B = 16'h00B0; #100;
A = 16'h00DC; B = 16'h00B1; #100;
A = 16'h00DC; B = 16'h00B2; #100;
A = 16'h00DC; B = 16'h00B3; #100;
A = 16'h00DC; B = 16'h00B4; #100;
A = 16'h00DC; B = 16'h00B5; #100;
A = 16'h00DC; B = 16'h00B6; #100;
A = 16'h00DC; B = 16'h00B7; #100;
A = 16'h00DC; B = 16'h00B8; #100;
A = 16'h00DC; B = 16'h00B9; #100;
A = 16'h00DC; B = 16'h00BA; #100;
A = 16'h00DC; B = 16'h00BB; #100;
A = 16'h00DC; B = 16'h00BC; #100;
A = 16'h00DC; B = 16'h00BD; #100;
A = 16'h00DC; B = 16'h00BE; #100;
A = 16'h00DC; B = 16'h00BF; #100;
A = 16'h00DC; B = 16'h00C0; #100;
A = 16'h00DC; B = 16'h00C1; #100;
A = 16'h00DC; B = 16'h00C2; #100;
A = 16'h00DC; B = 16'h00C3; #100;
A = 16'h00DC; B = 16'h00C4; #100;
A = 16'h00DC; B = 16'h00C5; #100;
A = 16'h00DC; B = 16'h00C6; #100;
A = 16'h00DC; B = 16'h00C7; #100;
A = 16'h00DC; B = 16'h00C8; #100;
A = 16'h00DC; B = 16'h00C9; #100;
A = 16'h00DC; B = 16'h00CA; #100;
A = 16'h00DC; B = 16'h00CB; #100;
A = 16'h00DC; B = 16'h00CC; #100;
A = 16'h00DC; B = 16'h00CD; #100;
A = 16'h00DC; B = 16'h00CE; #100;
A = 16'h00DC; B = 16'h00CF; #100;
A = 16'h00DC; B = 16'h00D0; #100;
A = 16'h00DC; B = 16'h00D1; #100;
A = 16'h00DC; B = 16'h00D2; #100;
A = 16'h00DC; B = 16'h00D3; #100;
A = 16'h00DC; B = 16'h00D4; #100;
A = 16'h00DC; B = 16'h00D5; #100;
A = 16'h00DC; B = 16'h00D6; #100;
A = 16'h00DC; B = 16'h00D7; #100;
A = 16'h00DC; B = 16'h00D8; #100;
A = 16'h00DC; B = 16'h00D9; #100;
A = 16'h00DC; B = 16'h00DA; #100;
A = 16'h00DC; B = 16'h00DB; #100;
A = 16'h00DC; B = 16'h00DC; #100;
A = 16'h00DC; B = 16'h00DD; #100;
A = 16'h00DC; B = 16'h00DE; #100;
A = 16'h00DC; B = 16'h00DF; #100;
A = 16'h00DC; B = 16'h00E0; #100;
A = 16'h00DC; B = 16'h00E1; #100;
A = 16'h00DC; B = 16'h00E2; #100;
A = 16'h00DC; B = 16'h00E3; #100;
A = 16'h00DC; B = 16'h00E4; #100;
A = 16'h00DC; B = 16'h00E5; #100;
A = 16'h00DC; B = 16'h00E6; #100;
A = 16'h00DC; B = 16'h00E7; #100;
A = 16'h00DC; B = 16'h00E8; #100;
A = 16'h00DC; B = 16'h00E9; #100;
A = 16'h00DC; B = 16'h00EA; #100;
A = 16'h00DC; B = 16'h00EB; #100;
A = 16'h00DC; B = 16'h00EC; #100;
A = 16'h00DC; B = 16'h00ED; #100;
A = 16'h00DC; B = 16'h00EE; #100;
A = 16'h00DC; B = 16'h00EF; #100;
A = 16'h00DC; B = 16'h00F0; #100;
A = 16'h00DC; B = 16'h00F1; #100;
A = 16'h00DC; B = 16'h00F2; #100;
A = 16'h00DC; B = 16'h00F3; #100;
A = 16'h00DC; B = 16'h00F4; #100;
A = 16'h00DC; B = 16'h00F5; #100;
A = 16'h00DC; B = 16'h00F6; #100;
A = 16'h00DC; B = 16'h00F7; #100;
A = 16'h00DC; B = 16'h00F8; #100;
A = 16'h00DC; B = 16'h00F9; #100;
A = 16'h00DC; B = 16'h00FA; #100;
A = 16'h00DC; B = 16'h00FB; #100;
A = 16'h00DC; B = 16'h00FC; #100;
A = 16'h00DC; B = 16'h00FD; #100;
A = 16'h00DC; B = 16'h00FE; #100;
A = 16'h00DC; B = 16'h00FF; #100;
A = 16'h00DD; B = 16'h000; #100;
A = 16'h00DD; B = 16'h001; #100;
A = 16'h00DD; B = 16'h002; #100;
A = 16'h00DD; B = 16'h003; #100;
A = 16'h00DD; B = 16'h004; #100;
A = 16'h00DD; B = 16'h005; #100;
A = 16'h00DD; B = 16'h006; #100;
A = 16'h00DD; B = 16'h007; #100;
A = 16'h00DD; B = 16'h008; #100;
A = 16'h00DD; B = 16'h009; #100;
A = 16'h00DD; B = 16'h00A; #100;
A = 16'h00DD; B = 16'h00B; #100;
A = 16'h00DD; B = 16'h00C; #100;
A = 16'h00DD; B = 16'h00D; #100;
A = 16'h00DD; B = 16'h00E; #100;
A = 16'h00DD; B = 16'h00F; #100;
A = 16'h00DD; B = 16'h0010; #100;
A = 16'h00DD; B = 16'h0011; #100;
A = 16'h00DD; B = 16'h0012; #100;
A = 16'h00DD; B = 16'h0013; #100;
A = 16'h00DD; B = 16'h0014; #100;
A = 16'h00DD; B = 16'h0015; #100;
A = 16'h00DD; B = 16'h0016; #100;
A = 16'h00DD; B = 16'h0017; #100;
A = 16'h00DD; B = 16'h0018; #100;
A = 16'h00DD; B = 16'h0019; #100;
A = 16'h00DD; B = 16'h001A; #100;
A = 16'h00DD; B = 16'h001B; #100;
A = 16'h00DD; B = 16'h001C; #100;
A = 16'h00DD; B = 16'h001D; #100;
A = 16'h00DD; B = 16'h001E; #100;
A = 16'h00DD; B = 16'h001F; #100;
A = 16'h00DD; B = 16'h0020; #100;
A = 16'h00DD; B = 16'h0021; #100;
A = 16'h00DD; B = 16'h0022; #100;
A = 16'h00DD; B = 16'h0023; #100;
A = 16'h00DD; B = 16'h0024; #100;
A = 16'h00DD; B = 16'h0025; #100;
A = 16'h00DD; B = 16'h0026; #100;
A = 16'h00DD; B = 16'h0027; #100;
A = 16'h00DD; B = 16'h0028; #100;
A = 16'h00DD; B = 16'h0029; #100;
A = 16'h00DD; B = 16'h002A; #100;
A = 16'h00DD; B = 16'h002B; #100;
A = 16'h00DD; B = 16'h002C; #100;
A = 16'h00DD; B = 16'h002D; #100;
A = 16'h00DD; B = 16'h002E; #100;
A = 16'h00DD; B = 16'h002F; #100;
A = 16'h00DD; B = 16'h0030; #100;
A = 16'h00DD; B = 16'h0031; #100;
A = 16'h00DD; B = 16'h0032; #100;
A = 16'h00DD; B = 16'h0033; #100;
A = 16'h00DD; B = 16'h0034; #100;
A = 16'h00DD; B = 16'h0035; #100;
A = 16'h00DD; B = 16'h0036; #100;
A = 16'h00DD; B = 16'h0037; #100;
A = 16'h00DD; B = 16'h0038; #100;
A = 16'h00DD; B = 16'h0039; #100;
A = 16'h00DD; B = 16'h003A; #100;
A = 16'h00DD; B = 16'h003B; #100;
A = 16'h00DD; B = 16'h003C; #100;
A = 16'h00DD; B = 16'h003D; #100;
A = 16'h00DD; B = 16'h003E; #100;
A = 16'h00DD; B = 16'h003F; #100;
A = 16'h00DD; B = 16'h0040; #100;
A = 16'h00DD; B = 16'h0041; #100;
A = 16'h00DD; B = 16'h0042; #100;
A = 16'h00DD; B = 16'h0043; #100;
A = 16'h00DD; B = 16'h0044; #100;
A = 16'h00DD; B = 16'h0045; #100;
A = 16'h00DD; B = 16'h0046; #100;
A = 16'h00DD; B = 16'h0047; #100;
A = 16'h00DD; B = 16'h0048; #100;
A = 16'h00DD; B = 16'h0049; #100;
A = 16'h00DD; B = 16'h004A; #100;
A = 16'h00DD; B = 16'h004B; #100;
A = 16'h00DD; B = 16'h004C; #100;
A = 16'h00DD; B = 16'h004D; #100;
A = 16'h00DD; B = 16'h004E; #100;
A = 16'h00DD; B = 16'h004F; #100;
A = 16'h00DD; B = 16'h0050; #100;
A = 16'h00DD; B = 16'h0051; #100;
A = 16'h00DD; B = 16'h0052; #100;
A = 16'h00DD; B = 16'h0053; #100;
A = 16'h00DD; B = 16'h0054; #100;
A = 16'h00DD; B = 16'h0055; #100;
A = 16'h00DD; B = 16'h0056; #100;
A = 16'h00DD; B = 16'h0057; #100;
A = 16'h00DD; B = 16'h0058; #100;
A = 16'h00DD; B = 16'h0059; #100;
A = 16'h00DD; B = 16'h005A; #100;
A = 16'h00DD; B = 16'h005B; #100;
A = 16'h00DD; B = 16'h005C; #100;
A = 16'h00DD; B = 16'h005D; #100;
A = 16'h00DD; B = 16'h005E; #100;
A = 16'h00DD; B = 16'h005F; #100;
A = 16'h00DD; B = 16'h0060; #100;
A = 16'h00DD; B = 16'h0061; #100;
A = 16'h00DD; B = 16'h0062; #100;
A = 16'h00DD; B = 16'h0063; #100;
A = 16'h00DD; B = 16'h0064; #100;
A = 16'h00DD; B = 16'h0065; #100;
A = 16'h00DD; B = 16'h0066; #100;
A = 16'h00DD; B = 16'h0067; #100;
A = 16'h00DD; B = 16'h0068; #100;
A = 16'h00DD; B = 16'h0069; #100;
A = 16'h00DD; B = 16'h006A; #100;
A = 16'h00DD; B = 16'h006B; #100;
A = 16'h00DD; B = 16'h006C; #100;
A = 16'h00DD; B = 16'h006D; #100;
A = 16'h00DD; B = 16'h006E; #100;
A = 16'h00DD; B = 16'h006F; #100;
A = 16'h00DD; B = 16'h0070; #100;
A = 16'h00DD; B = 16'h0071; #100;
A = 16'h00DD; B = 16'h0072; #100;
A = 16'h00DD; B = 16'h0073; #100;
A = 16'h00DD; B = 16'h0074; #100;
A = 16'h00DD; B = 16'h0075; #100;
A = 16'h00DD; B = 16'h0076; #100;
A = 16'h00DD; B = 16'h0077; #100;
A = 16'h00DD; B = 16'h0078; #100;
A = 16'h00DD; B = 16'h0079; #100;
A = 16'h00DD; B = 16'h007A; #100;
A = 16'h00DD; B = 16'h007B; #100;
A = 16'h00DD; B = 16'h007C; #100;
A = 16'h00DD; B = 16'h007D; #100;
A = 16'h00DD; B = 16'h007E; #100;
A = 16'h00DD; B = 16'h007F; #100;
A = 16'h00DD; B = 16'h0080; #100;
A = 16'h00DD; B = 16'h0081; #100;
A = 16'h00DD; B = 16'h0082; #100;
A = 16'h00DD; B = 16'h0083; #100;
A = 16'h00DD; B = 16'h0084; #100;
A = 16'h00DD; B = 16'h0085; #100;
A = 16'h00DD; B = 16'h0086; #100;
A = 16'h00DD; B = 16'h0087; #100;
A = 16'h00DD; B = 16'h0088; #100;
A = 16'h00DD; B = 16'h0089; #100;
A = 16'h00DD; B = 16'h008A; #100;
A = 16'h00DD; B = 16'h008B; #100;
A = 16'h00DD; B = 16'h008C; #100;
A = 16'h00DD; B = 16'h008D; #100;
A = 16'h00DD; B = 16'h008E; #100;
A = 16'h00DD; B = 16'h008F; #100;
A = 16'h00DD; B = 16'h0090; #100;
A = 16'h00DD; B = 16'h0091; #100;
A = 16'h00DD; B = 16'h0092; #100;
A = 16'h00DD; B = 16'h0093; #100;
A = 16'h00DD; B = 16'h0094; #100;
A = 16'h00DD; B = 16'h0095; #100;
A = 16'h00DD; B = 16'h0096; #100;
A = 16'h00DD; B = 16'h0097; #100;
A = 16'h00DD; B = 16'h0098; #100;
A = 16'h00DD; B = 16'h0099; #100;
A = 16'h00DD; B = 16'h009A; #100;
A = 16'h00DD; B = 16'h009B; #100;
A = 16'h00DD; B = 16'h009C; #100;
A = 16'h00DD; B = 16'h009D; #100;
A = 16'h00DD; B = 16'h009E; #100;
A = 16'h00DD; B = 16'h009F; #100;
A = 16'h00DD; B = 16'h00A0; #100;
A = 16'h00DD; B = 16'h00A1; #100;
A = 16'h00DD; B = 16'h00A2; #100;
A = 16'h00DD; B = 16'h00A3; #100;
A = 16'h00DD; B = 16'h00A4; #100;
A = 16'h00DD; B = 16'h00A5; #100;
A = 16'h00DD; B = 16'h00A6; #100;
A = 16'h00DD; B = 16'h00A7; #100;
A = 16'h00DD; B = 16'h00A8; #100;
A = 16'h00DD; B = 16'h00A9; #100;
A = 16'h00DD; B = 16'h00AA; #100;
A = 16'h00DD; B = 16'h00AB; #100;
A = 16'h00DD; B = 16'h00AC; #100;
A = 16'h00DD; B = 16'h00AD; #100;
A = 16'h00DD; B = 16'h00AE; #100;
A = 16'h00DD; B = 16'h00AF; #100;
A = 16'h00DD; B = 16'h00B0; #100;
A = 16'h00DD; B = 16'h00B1; #100;
A = 16'h00DD; B = 16'h00B2; #100;
A = 16'h00DD; B = 16'h00B3; #100;
A = 16'h00DD; B = 16'h00B4; #100;
A = 16'h00DD; B = 16'h00B5; #100;
A = 16'h00DD; B = 16'h00B6; #100;
A = 16'h00DD; B = 16'h00B7; #100;
A = 16'h00DD; B = 16'h00B8; #100;
A = 16'h00DD; B = 16'h00B9; #100;
A = 16'h00DD; B = 16'h00BA; #100;
A = 16'h00DD; B = 16'h00BB; #100;
A = 16'h00DD; B = 16'h00BC; #100;
A = 16'h00DD; B = 16'h00BD; #100;
A = 16'h00DD; B = 16'h00BE; #100;
A = 16'h00DD; B = 16'h00BF; #100;
A = 16'h00DD; B = 16'h00C0; #100;
A = 16'h00DD; B = 16'h00C1; #100;
A = 16'h00DD; B = 16'h00C2; #100;
A = 16'h00DD; B = 16'h00C3; #100;
A = 16'h00DD; B = 16'h00C4; #100;
A = 16'h00DD; B = 16'h00C5; #100;
A = 16'h00DD; B = 16'h00C6; #100;
A = 16'h00DD; B = 16'h00C7; #100;
A = 16'h00DD; B = 16'h00C8; #100;
A = 16'h00DD; B = 16'h00C9; #100;
A = 16'h00DD; B = 16'h00CA; #100;
A = 16'h00DD; B = 16'h00CB; #100;
A = 16'h00DD; B = 16'h00CC; #100;
A = 16'h00DD; B = 16'h00CD; #100;
A = 16'h00DD; B = 16'h00CE; #100;
A = 16'h00DD; B = 16'h00CF; #100;
A = 16'h00DD; B = 16'h00D0; #100;
A = 16'h00DD; B = 16'h00D1; #100;
A = 16'h00DD; B = 16'h00D2; #100;
A = 16'h00DD; B = 16'h00D3; #100;
A = 16'h00DD; B = 16'h00D4; #100;
A = 16'h00DD; B = 16'h00D5; #100;
A = 16'h00DD; B = 16'h00D6; #100;
A = 16'h00DD; B = 16'h00D7; #100;
A = 16'h00DD; B = 16'h00D8; #100;
A = 16'h00DD; B = 16'h00D9; #100;
A = 16'h00DD; B = 16'h00DA; #100;
A = 16'h00DD; B = 16'h00DB; #100;
A = 16'h00DD; B = 16'h00DC; #100;
A = 16'h00DD; B = 16'h00DD; #100;
A = 16'h00DD; B = 16'h00DE; #100;
A = 16'h00DD; B = 16'h00DF; #100;
A = 16'h00DD; B = 16'h00E0; #100;
A = 16'h00DD; B = 16'h00E1; #100;
A = 16'h00DD; B = 16'h00E2; #100;
A = 16'h00DD; B = 16'h00E3; #100;
A = 16'h00DD; B = 16'h00E4; #100;
A = 16'h00DD; B = 16'h00E5; #100;
A = 16'h00DD; B = 16'h00E6; #100;
A = 16'h00DD; B = 16'h00E7; #100;
A = 16'h00DD; B = 16'h00E8; #100;
A = 16'h00DD; B = 16'h00E9; #100;
A = 16'h00DD; B = 16'h00EA; #100;
A = 16'h00DD; B = 16'h00EB; #100;
A = 16'h00DD; B = 16'h00EC; #100;
A = 16'h00DD; B = 16'h00ED; #100;
A = 16'h00DD; B = 16'h00EE; #100;
A = 16'h00DD; B = 16'h00EF; #100;
A = 16'h00DD; B = 16'h00F0; #100;
A = 16'h00DD; B = 16'h00F1; #100;
A = 16'h00DD; B = 16'h00F2; #100;
A = 16'h00DD; B = 16'h00F3; #100;
A = 16'h00DD; B = 16'h00F4; #100;
A = 16'h00DD; B = 16'h00F5; #100;
A = 16'h00DD; B = 16'h00F6; #100;
A = 16'h00DD; B = 16'h00F7; #100;
A = 16'h00DD; B = 16'h00F8; #100;
A = 16'h00DD; B = 16'h00F9; #100;
A = 16'h00DD; B = 16'h00FA; #100;
A = 16'h00DD; B = 16'h00FB; #100;
A = 16'h00DD; B = 16'h00FC; #100;
A = 16'h00DD; B = 16'h00FD; #100;
A = 16'h00DD; B = 16'h00FE; #100;
A = 16'h00DD; B = 16'h00FF; #100;
A = 16'h00DE; B = 16'h000; #100;
A = 16'h00DE; B = 16'h001; #100;
A = 16'h00DE; B = 16'h002; #100;
A = 16'h00DE; B = 16'h003; #100;
A = 16'h00DE; B = 16'h004; #100;
A = 16'h00DE; B = 16'h005; #100;
A = 16'h00DE; B = 16'h006; #100;
A = 16'h00DE; B = 16'h007; #100;
A = 16'h00DE; B = 16'h008; #100;
A = 16'h00DE; B = 16'h009; #100;
A = 16'h00DE; B = 16'h00A; #100;
A = 16'h00DE; B = 16'h00B; #100;
A = 16'h00DE; B = 16'h00C; #100;
A = 16'h00DE; B = 16'h00D; #100;
A = 16'h00DE; B = 16'h00E; #100;
A = 16'h00DE; B = 16'h00F; #100;
A = 16'h00DE; B = 16'h0010; #100;
A = 16'h00DE; B = 16'h0011; #100;
A = 16'h00DE; B = 16'h0012; #100;
A = 16'h00DE; B = 16'h0013; #100;
A = 16'h00DE; B = 16'h0014; #100;
A = 16'h00DE; B = 16'h0015; #100;
A = 16'h00DE; B = 16'h0016; #100;
A = 16'h00DE; B = 16'h0017; #100;
A = 16'h00DE; B = 16'h0018; #100;
A = 16'h00DE; B = 16'h0019; #100;
A = 16'h00DE; B = 16'h001A; #100;
A = 16'h00DE; B = 16'h001B; #100;
A = 16'h00DE; B = 16'h001C; #100;
A = 16'h00DE; B = 16'h001D; #100;
A = 16'h00DE; B = 16'h001E; #100;
A = 16'h00DE; B = 16'h001F; #100;
A = 16'h00DE; B = 16'h0020; #100;
A = 16'h00DE; B = 16'h0021; #100;
A = 16'h00DE; B = 16'h0022; #100;
A = 16'h00DE; B = 16'h0023; #100;
A = 16'h00DE; B = 16'h0024; #100;
A = 16'h00DE; B = 16'h0025; #100;
A = 16'h00DE; B = 16'h0026; #100;
A = 16'h00DE; B = 16'h0027; #100;
A = 16'h00DE; B = 16'h0028; #100;
A = 16'h00DE; B = 16'h0029; #100;
A = 16'h00DE; B = 16'h002A; #100;
A = 16'h00DE; B = 16'h002B; #100;
A = 16'h00DE; B = 16'h002C; #100;
A = 16'h00DE; B = 16'h002D; #100;
A = 16'h00DE; B = 16'h002E; #100;
A = 16'h00DE; B = 16'h002F; #100;
A = 16'h00DE; B = 16'h0030; #100;
A = 16'h00DE; B = 16'h0031; #100;
A = 16'h00DE; B = 16'h0032; #100;
A = 16'h00DE; B = 16'h0033; #100;
A = 16'h00DE; B = 16'h0034; #100;
A = 16'h00DE; B = 16'h0035; #100;
A = 16'h00DE; B = 16'h0036; #100;
A = 16'h00DE; B = 16'h0037; #100;
A = 16'h00DE; B = 16'h0038; #100;
A = 16'h00DE; B = 16'h0039; #100;
A = 16'h00DE; B = 16'h003A; #100;
A = 16'h00DE; B = 16'h003B; #100;
A = 16'h00DE; B = 16'h003C; #100;
A = 16'h00DE; B = 16'h003D; #100;
A = 16'h00DE; B = 16'h003E; #100;
A = 16'h00DE; B = 16'h003F; #100;
A = 16'h00DE; B = 16'h0040; #100;
A = 16'h00DE; B = 16'h0041; #100;
A = 16'h00DE; B = 16'h0042; #100;
A = 16'h00DE; B = 16'h0043; #100;
A = 16'h00DE; B = 16'h0044; #100;
A = 16'h00DE; B = 16'h0045; #100;
A = 16'h00DE; B = 16'h0046; #100;
A = 16'h00DE; B = 16'h0047; #100;
A = 16'h00DE; B = 16'h0048; #100;
A = 16'h00DE; B = 16'h0049; #100;
A = 16'h00DE; B = 16'h004A; #100;
A = 16'h00DE; B = 16'h004B; #100;
A = 16'h00DE; B = 16'h004C; #100;
A = 16'h00DE; B = 16'h004D; #100;
A = 16'h00DE; B = 16'h004E; #100;
A = 16'h00DE; B = 16'h004F; #100;
A = 16'h00DE; B = 16'h0050; #100;
A = 16'h00DE; B = 16'h0051; #100;
A = 16'h00DE; B = 16'h0052; #100;
A = 16'h00DE; B = 16'h0053; #100;
A = 16'h00DE; B = 16'h0054; #100;
A = 16'h00DE; B = 16'h0055; #100;
A = 16'h00DE; B = 16'h0056; #100;
A = 16'h00DE; B = 16'h0057; #100;
A = 16'h00DE; B = 16'h0058; #100;
A = 16'h00DE; B = 16'h0059; #100;
A = 16'h00DE; B = 16'h005A; #100;
A = 16'h00DE; B = 16'h005B; #100;
A = 16'h00DE; B = 16'h005C; #100;
A = 16'h00DE; B = 16'h005D; #100;
A = 16'h00DE; B = 16'h005E; #100;
A = 16'h00DE; B = 16'h005F; #100;
A = 16'h00DE; B = 16'h0060; #100;
A = 16'h00DE; B = 16'h0061; #100;
A = 16'h00DE; B = 16'h0062; #100;
A = 16'h00DE; B = 16'h0063; #100;
A = 16'h00DE; B = 16'h0064; #100;
A = 16'h00DE; B = 16'h0065; #100;
A = 16'h00DE; B = 16'h0066; #100;
A = 16'h00DE; B = 16'h0067; #100;
A = 16'h00DE; B = 16'h0068; #100;
A = 16'h00DE; B = 16'h0069; #100;
A = 16'h00DE; B = 16'h006A; #100;
A = 16'h00DE; B = 16'h006B; #100;
A = 16'h00DE; B = 16'h006C; #100;
A = 16'h00DE; B = 16'h006D; #100;
A = 16'h00DE; B = 16'h006E; #100;
A = 16'h00DE; B = 16'h006F; #100;
A = 16'h00DE; B = 16'h0070; #100;
A = 16'h00DE; B = 16'h0071; #100;
A = 16'h00DE; B = 16'h0072; #100;
A = 16'h00DE; B = 16'h0073; #100;
A = 16'h00DE; B = 16'h0074; #100;
A = 16'h00DE; B = 16'h0075; #100;
A = 16'h00DE; B = 16'h0076; #100;
A = 16'h00DE; B = 16'h0077; #100;
A = 16'h00DE; B = 16'h0078; #100;
A = 16'h00DE; B = 16'h0079; #100;
A = 16'h00DE; B = 16'h007A; #100;
A = 16'h00DE; B = 16'h007B; #100;
A = 16'h00DE; B = 16'h007C; #100;
A = 16'h00DE; B = 16'h007D; #100;
A = 16'h00DE; B = 16'h007E; #100;
A = 16'h00DE; B = 16'h007F; #100;
A = 16'h00DE; B = 16'h0080; #100;
A = 16'h00DE; B = 16'h0081; #100;
A = 16'h00DE; B = 16'h0082; #100;
A = 16'h00DE; B = 16'h0083; #100;
A = 16'h00DE; B = 16'h0084; #100;
A = 16'h00DE; B = 16'h0085; #100;
A = 16'h00DE; B = 16'h0086; #100;
A = 16'h00DE; B = 16'h0087; #100;
A = 16'h00DE; B = 16'h0088; #100;
A = 16'h00DE; B = 16'h0089; #100;
A = 16'h00DE; B = 16'h008A; #100;
A = 16'h00DE; B = 16'h008B; #100;
A = 16'h00DE; B = 16'h008C; #100;
A = 16'h00DE; B = 16'h008D; #100;
A = 16'h00DE; B = 16'h008E; #100;
A = 16'h00DE; B = 16'h008F; #100;
A = 16'h00DE; B = 16'h0090; #100;
A = 16'h00DE; B = 16'h0091; #100;
A = 16'h00DE; B = 16'h0092; #100;
A = 16'h00DE; B = 16'h0093; #100;
A = 16'h00DE; B = 16'h0094; #100;
A = 16'h00DE; B = 16'h0095; #100;
A = 16'h00DE; B = 16'h0096; #100;
A = 16'h00DE; B = 16'h0097; #100;
A = 16'h00DE; B = 16'h0098; #100;
A = 16'h00DE; B = 16'h0099; #100;
A = 16'h00DE; B = 16'h009A; #100;
A = 16'h00DE; B = 16'h009B; #100;
A = 16'h00DE; B = 16'h009C; #100;
A = 16'h00DE; B = 16'h009D; #100;
A = 16'h00DE; B = 16'h009E; #100;
A = 16'h00DE; B = 16'h009F; #100;
A = 16'h00DE; B = 16'h00A0; #100;
A = 16'h00DE; B = 16'h00A1; #100;
A = 16'h00DE; B = 16'h00A2; #100;
A = 16'h00DE; B = 16'h00A3; #100;
A = 16'h00DE; B = 16'h00A4; #100;
A = 16'h00DE; B = 16'h00A5; #100;
A = 16'h00DE; B = 16'h00A6; #100;
A = 16'h00DE; B = 16'h00A7; #100;
A = 16'h00DE; B = 16'h00A8; #100;
A = 16'h00DE; B = 16'h00A9; #100;
A = 16'h00DE; B = 16'h00AA; #100;
A = 16'h00DE; B = 16'h00AB; #100;
A = 16'h00DE; B = 16'h00AC; #100;
A = 16'h00DE; B = 16'h00AD; #100;
A = 16'h00DE; B = 16'h00AE; #100;
A = 16'h00DE; B = 16'h00AF; #100;
A = 16'h00DE; B = 16'h00B0; #100;
A = 16'h00DE; B = 16'h00B1; #100;
A = 16'h00DE; B = 16'h00B2; #100;
A = 16'h00DE; B = 16'h00B3; #100;
A = 16'h00DE; B = 16'h00B4; #100;
A = 16'h00DE; B = 16'h00B5; #100;
A = 16'h00DE; B = 16'h00B6; #100;
A = 16'h00DE; B = 16'h00B7; #100;
A = 16'h00DE; B = 16'h00B8; #100;
A = 16'h00DE; B = 16'h00B9; #100;
A = 16'h00DE; B = 16'h00BA; #100;
A = 16'h00DE; B = 16'h00BB; #100;
A = 16'h00DE; B = 16'h00BC; #100;
A = 16'h00DE; B = 16'h00BD; #100;
A = 16'h00DE; B = 16'h00BE; #100;
A = 16'h00DE; B = 16'h00BF; #100;
A = 16'h00DE; B = 16'h00C0; #100;
A = 16'h00DE; B = 16'h00C1; #100;
A = 16'h00DE; B = 16'h00C2; #100;
A = 16'h00DE; B = 16'h00C3; #100;
A = 16'h00DE; B = 16'h00C4; #100;
A = 16'h00DE; B = 16'h00C5; #100;
A = 16'h00DE; B = 16'h00C6; #100;
A = 16'h00DE; B = 16'h00C7; #100;
A = 16'h00DE; B = 16'h00C8; #100;
A = 16'h00DE; B = 16'h00C9; #100;
A = 16'h00DE; B = 16'h00CA; #100;
A = 16'h00DE; B = 16'h00CB; #100;
A = 16'h00DE; B = 16'h00CC; #100;
A = 16'h00DE; B = 16'h00CD; #100;
A = 16'h00DE; B = 16'h00CE; #100;
A = 16'h00DE; B = 16'h00CF; #100;
A = 16'h00DE; B = 16'h00D0; #100;
A = 16'h00DE; B = 16'h00D1; #100;
A = 16'h00DE; B = 16'h00D2; #100;
A = 16'h00DE; B = 16'h00D3; #100;
A = 16'h00DE; B = 16'h00D4; #100;
A = 16'h00DE; B = 16'h00D5; #100;
A = 16'h00DE; B = 16'h00D6; #100;
A = 16'h00DE; B = 16'h00D7; #100;
A = 16'h00DE; B = 16'h00D8; #100;
A = 16'h00DE; B = 16'h00D9; #100;
A = 16'h00DE; B = 16'h00DA; #100;
A = 16'h00DE; B = 16'h00DB; #100;
A = 16'h00DE; B = 16'h00DC; #100;
A = 16'h00DE; B = 16'h00DD; #100;
A = 16'h00DE; B = 16'h00DE; #100;
A = 16'h00DE; B = 16'h00DF; #100;
A = 16'h00DE; B = 16'h00E0; #100;
A = 16'h00DE; B = 16'h00E1; #100;
A = 16'h00DE; B = 16'h00E2; #100;
A = 16'h00DE; B = 16'h00E3; #100;
A = 16'h00DE; B = 16'h00E4; #100;
A = 16'h00DE; B = 16'h00E5; #100;
A = 16'h00DE; B = 16'h00E6; #100;
A = 16'h00DE; B = 16'h00E7; #100;
A = 16'h00DE; B = 16'h00E8; #100;
A = 16'h00DE; B = 16'h00E9; #100;
A = 16'h00DE; B = 16'h00EA; #100;
A = 16'h00DE; B = 16'h00EB; #100;
A = 16'h00DE; B = 16'h00EC; #100;
A = 16'h00DE; B = 16'h00ED; #100;
A = 16'h00DE; B = 16'h00EE; #100;
A = 16'h00DE; B = 16'h00EF; #100;
A = 16'h00DE; B = 16'h00F0; #100;
A = 16'h00DE; B = 16'h00F1; #100;
A = 16'h00DE; B = 16'h00F2; #100;
A = 16'h00DE; B = 16'h00F3; #100;
A = 16'h00DE; B = 16'h00F4; #100;
A = 16'h00DE; B = 16'h00F5; #100;
A = 16'h00DE; B = 16'h00F6; #100;
A = 16'h00DE; B = 16'h00F7; #100;
A = 16'h00DE; B = 16'h00F8; #100;
A = 16'h00DE; B = 16'h00F9; #100;
A = 16'h00DE; B = 16'h00FA; #100;
A = 16'h00DE; B = 16'h00FB; #100;
A = 16'h00DE; B = 16'h00FC; #100;
A = 16'h00DE; B = 16'h00FD; #100;
A = 16'h00DE; B = 16'h00FE; #100;
A = 16'h00DE; B = 16'h00FF; #100;
A = 16'h00DF; B = 16'h000; #100;
A = 16'h00DF; B = 16'h001; #100;
A = 16'h00DF; B = 16'h002; #100;
A = 16'h00DF; B = 16'h003; #100;
A = 16'h00DF; B = 16'h004; #100;
A = 16'h00DF; B = 16'h005; #100;
A = 16'h00DF; B = 16'h006; #100;
A = 16'h00DF; B = 16'h007; #100;
A = 16'h00DF; B = 16'h008; #100;
A = 16'h00DF; B = 16'h009; #100;
A = 16'h00DF; B = 16'h00A; #100;
A = 16'h00DF; B = 16'h00B; #100;
A = 16'h00DF; B = 16'h00C; #100;
A = 16'h00DF; B = 16'h00D; #100;
A = 16'h00DF; B = 16'h00E; #100;
A = 16'h00DF; B = 16'h00F; #100;
A = 16'h00DF; B = 16'h0010; #100;
A = 16'h00DF; B = 16'h0011; #100;
A = 16'h00DF; B = 16'h0012; #100;
A = 16'h00DF; B = 16'h0013; #100;
A = 16'h00DF; B = 16'h0014; #100;
A = 16'h00DF; B = 16'h0015; #100;
A = 16'h00DF; B = 16'h0016; #100;
A = 16'h00DF; B = 16'h0017; #100;
A = 16'h00DF; B = 16'h0018; #100;
A = 16'h00DF; B = 16'h0019; #100;
A = 16'h00DF; B = 16'h001A; #100;
A = 16'h00DF; B = 16'h001B; #100;
A = 16'h00DF; B = 16'h001C; #100;
A = 16'h00DF; B = 16'h001D; #100;
A = 16'h00DF; B = 16'h001E; #100;
A = 16'h00DF; B = 16'h001F; #100;
A = 16'h00DF; B = 16'h0020; #100;
A = 16'h00DF; B = 16'h0021; #100;
A = 16'h00DF; B = 16'h0022; #100;
A = 16'h00DF; B = 16'h0023; #100;
A = 16'h00DF; B = 16'h0024; #100;
A = 16'h00DF; B = 16'h0025; #100;
A = 16'h00DF; B = 16'h0026; #100;
A = 16'h00DF; B = 16'h0027; #100;
A = 16'h00DF; B = 16'h0028; #100;
A = 16'h00DF; B = 16'h0029; #100;
A = 16'h00DF; B = 16'h002A; #100;
A = 16'h00DF; B = 16'h002B; #100;
A = 16'h00DF; B = 16'h002C; #100;
A = 16'h00DF; B = 16'h002D; #100;
A = 16'h00DF; B = 16'h002E; #100;
A = 16'h00DF; B = 16'h002F; #100;
A = 16'h00DF; B = 16'h0030; #100;
A = 16'h00DF; B = 16'h0031; #100;
A = 16'h00DF; B = 16'h0032; #100;
A = 16'h00DF; B = 16'h0033; #100;
A = 16'h00DF; B = 16'h0034; #100;
A = 16'h00DF; B = 16'h0035; #100;
A = 16'h00DF; B = 16'h0036; #100;
A = 16'h00DF; B = 16'h0037; #100;
A = 16'h00DF; B = 16'h0038; #100;
A = 16'h00DF; B = 16'h0039; #100;
A = 16'h00DF; B = 16'h003A; #100;
A = 16'h00DF; B = 16'h003B; #100;
A = 16'h00DF; B = 16'h003C; #100;
A = 16'h00DF; B = 16'h003D; #100;
A = 16'h00DF; B = 16'h003E; #100;
A = 16'h00DF; B = 16'h003F; #100;
A = 16'h00DF; B = 16'h0040; #100;
A = 16'h00DF; B = 16'h0041; #100;
A = 16'h00DF; B = 16'h0042; #100;
A = 16'h00DF; B = 16'h0043; #100;
A = 16'h00DF; B = 16'h0044; #100;
A = 16'h00DF; B = 16'h0045; #100;
A = 16'h00DF; B = 16'h0046; #100;
A = 16'h00DF; B = 16'h0047; #100;
A = 16'h00DF; B = 16'h0048; #100;
A = 16'h00DF; B = 16'h0049; #100;
A = 16'h00DF; B = 16'h004A; #100;
A = 16'h00DF; B = 16'h004B; #100;
A = 16'h00DF; B = 16'h004C; #100;
A = 16'h00DF; B = 16'h004D; #100;
A = 16'h00DF; B = 16'h004E; #100;
A = 16'h00DF; B = 16'h004F; #100;
A = 16'h00DF; B = 16'h0050; #100;
A = 16'h00DF; B = 16'h0051; #100;
A = 16'h00DF; B = 16'h0052; #100;
A = 16'h00DF; B = 16'h0053; #100;
A = 16'h00DF; B = 16'h0054; #100;
A = 16'h00DF; B = 16'h0055; #100;
A = 16'h00DF; B = 16'h0056; #100;
A = 16'h00DF; B = 16'h0057; #100;
A = 16'h00DF; B = 16'h0058; #100;
A = 16'h00DF; B = 16'h0059; #100;
A = 16'h00DF; B = 16'h005A; #100;
A = 16'h00DF; B = 16'h005B; #100;
A = 16'h00DF; B = 16'h005C; #100;
A = 16'h00DF; B = 16'h005D; #100;
A = 16'h00DF; B = 16'h005E; #100;
A = 16'h00DF; B = 16'h005F; #100;
A = 16'h00DF; B = 16'h0060; #100;
A = 16'h00DF; B = 16'h0061; #100;
A = 16'h00DF; B = 16'h0062; #100;
A = 16'h00DF; B = 16'h0063; #100;
A = 16'h00DF; B = 16'h0064; #100;
A = 16'h00DF; B = 16'h0065; #100;
A = 16'h00DF; B = 16'h0066; #100;
A = 16'h00DF; B = 16'h0067; #100;
A = 16'h00DF; B = 16'h0068; #100;
A = 16'h00DF; B = 16'h0069; #100;
A = 16'h00DF; B = 16'h006A; #100;
A = 16'h00DF; B = 16'h006B; #100;
A = 16'h00DF; B = 16'h006C; #100;
A = 16'h00DF; B = 16'h006D; #100;
A = 16'h00DF; B = 16'h006E; #100;
A = 16'h00DF; B = 16'h006F; #100;
A = 16'h00DF; B = 16'h0070; #100;
A = 16'h00DF; B = 16'h0071; #100;
A = 16'h00DF; B = 16'h0072; #100;
A = 16'h00DF; B = 16'h0073; #100;
A = 16'h00DF; B = 16'h0074; #100;
A = 16'h00DF; B = 16'h0075; #100;
A = 16'h00DF; B = 16'h0076; #100;
A = 16'h00DF; B = 16'h0077; #100;
A = 16'h00DF; B = 16'h0078; #100;
A = 16'h00DF; B = 16'h0079; #100;
A = 16'h00DF; B = 16'h007A; #100;
A = 16'h00DF; B = 16'h007B; #100;
A = 16'h00DF; B = 16'h007C; #100;
A = 16'h00DF; B = 16'h007D; #100;
A = 16'h00DF; B = 16'h007E; #100;
A = 16'h00DF; B = 16'h007F; #100;
A = 16'h00DF; B = 16'h0080; #100;
A = 16'h00DF; B = 16'h0081; #100;
A = 16'h00DF; B = 16'h0082; #100;
A = 16'h00DF; B = 16'h0083; #100;
A = 16'h00DF; B = 16'h0084; #100;
A = 16'h00DF; B = 16'h0085; #100;
A = 16'h00DF; B = 16'h0086; #100;
A = 16'h00DF; B = 16'h0087; #100;
A = 16'h00DF; B = 16'h0088; #100;
A = 16'h00DF; B = 16'h0089; #100;
A = 16'h00DF; B = 16'h008A; #100;
A = 16'h00DF; B = 16'h008B; #100;
A = 16'h00DF; B = 16'h008C; #100;
A = 16'h00DF; B = 16'h008D; #100;
A = 16'h00DF; B = 16'h008E; #100;
A = 16'h00DF; B = 16'h008F; #100;
A = 16'h00DF; B = 16'h0090; #100;
A = 16'h00DF; B = 16'h0091; #100;
A = 16'h00DF; B = 16'h0092; #100;
A = 16'h00DF; B = 16'h0093; #100;
A = 16'h00DF; B = 16'h0094; #100;
A = 16'h00DF; B = 16'h0095; #100;
A = 16'h00DF; B = 16'h0096; #100;
A = 16'h00DF; B = 16'h0097; #100;
A = 16'h00DF; B = 16'h0098; #100;
A = 16'h00DF; B = 16'h0099; #100;
A = 16'h00DF; B = 16'h009A; #100;
A = 16'h00DF; B = 16'h009B; #100;
A = 16'h00DF; B = 16'h009C; #100;
A = 16'h00DF; B = 16'h009D; #100;
A = 16'h00DF; B = 16'h009E; #100;
A = 16'h00DF; B = 16'h009F; #100;
A = 16'h00DF; B = 16'h00A0; #100;
A = 16'h00DF; B = 16'h00A1; #100;
A = 16'h00DF; B = 16'h00A2; #100;
A = 16'h00DF; B = 16'h00A3; #100;
A = 16'h00DF; B = 16'h00A4; #100;
A = 16'h00DF; B = 16'h00A5; #100;
A = 16'h00DF; B = 16'h00A6; #100;
A = 16'h00DF; B = 16'h00A7; #100;
A = 16'h00DF; B = 16'h00A8; #100;
A = 16'h00DF; B = 16'h00A9; #100;
A = 16'h00DF; B = 16'h00AA; #100;
A = 16'h00DF; B = 16'h00AB; #100;
A = 16'h00DF; B = 16'h00AC; #100;
A = 16'h00DF; B = 16'h00AD; #100;
A = 16'h00DF; B = 16'h00AE; #100;
A = 16'h00DF; B = 16'h00AF; #100;
A = 16'h00DF; B = 16'h00B0; #100;
A = 16'h00DF; B = 16'h00B1; #100;
A = 16'h00DF; B = 16'h00B2; #100;
A = 16'h00DF; B = 16'h00B3; #100;
A = 16'h00DF; B = 16'h00B4; #100;
A = 16'h00DF; B = 16'h00B5; #100;
A = 16'h00DF; B = 16'h00B6; #100;
A = 16'h00DF; B = 16'h00B7; #100;
A = 16'h00DF; B = 16'h00B8; #100;
A = 16'h00DF; B = 16'h00B9; #100;
A = 16'h00DF; B = 16'h00BA; #100;
A = 16'h00DF; B = 16'h00BB; #100;
A = 16'h00DF; B = 16'h00BC; #100;
A = 16'h00DF; B = 16'h00BD; #100;
A = 16'h00DF; B = 16'h00BE; #100;
A = 16'h00DF; B = 16'h00BF; #100;
A = 16'h00DF; B = 16'h00C0; #100;
A = 16'h00DF; B = 16'h00C1; #100;
A = 16'h00DF; B = 16'h00C2; #100;
A = 16'h00DF; B = 16'h00C3; #100;
A = 16'h00DF; B = 16'h00C4; #100;
A = 16'h00DF; B = 16'h00C5; #100;
A = 16'h00DF; B = 16'h00C6; #100;
A = 16'h00DF; B = 16'h00C7; #100;
A = 16'h00DF; B = 16'h00C8; #100;
A = 16'h00DF; B = 16'h00C9; #100;
A = 16'h00DF; B = 16'h00CA; #100;
A = 16'h00DF; B = 16'h00CB; #100;
A = 16'h00DF; B = 16'h00CC; #100;
A = 16'h00DF; B = 16'h00CD; #100;
A = 16'h00DF; B = 16'h00CE; #100;
A = 16'h00DF; B = 16'h00CF; #100;
A = 16'h00DF; B = 16'h00D0; #100;
A = 16'h00DF; B = 16'h00D1; #100;
A = 16'h00DF; B = 16'h00D2; #100;
A = 16'h00DF; B = 16'h00D3; #100;
A = 16'h00DF; B = 16'h00D4; #100;
A = 16'h00DF; B = 16'h00D5; #100;
A = 16'h00DF; B = 16'h00D6; #100;
A = 16'h00DF; B = 16'h00D7; #100;
A = 16'h00DF; B = 16'h00D8; #100;
A = 16'h00DF; B = 16'h00D9; #100;
A = 16'h00DF; B = 16'h00DA; #100;
A = 16'h00DF; B = 16'h00DB; #100;
A = 16'h00DF; B = 16'h00DC; #100;
A = 16'h00DF; B = 16'h00DD; #100;
A = 16'h00DF; B = 16'h00DE; #100;
A = 16'h00DF; B = 16'h00DF; #100;
A = 16'h00DF; B = 16'h00E0; #100;
A = 16'h00DF; B = 16'h00E1; #100;
A = 16'h00DF; B = 16'h00E2; #100;
A = 16'h00DF; B = 16'h00E3; #100;
A = 16'h00DF; B = 16'h00E4; #100;
A = 16'h00DF; B = 16'h00E5; #100;
A = 16'h00DF; B = 16'h00E6; #100;
A = 16'h00DF; B = 16'h00E7; #100;
A = 16'h00DF; B = 16'h00E8; #100;
A = 16'h00DF; B = 16'h00E9; #100;
A = 16'h00DF; B = 16'h00EA; #100;
A = 16'h00DF; B = 16'h00EB; #100;
A = 16'h00DF; B = 16'h00EC; #100;
A = 16'h00DF; B = 16'h00ED; #100;
A = 16'h00DF; B = 16'h00EE; #100;
A = 16'h00DF; B = 16'h00EF; #100;
A = 16'h00DF; B = 16'h00F0; #100;
A = 16'h00DF; B = 16'h00F1; #100;
A = 16'h00DF; B = 16'h00F2; #100;
A = 16'h00DF; B = 16'h00F3; #100;
A = 16'h00DF; B = 16'h00F4; #100;
A = 16'h00DF; B = 16'h00F5; #100;
A = 16'h00DF; B = 16'h00F6; #100;
A = 16'h00DF; B = 16'h00F7; #100;
A = 16'h00DF; B = 16'h00F8; #100;
A = 16'h00DF; B = 16'h00F9; #100;
A = 16'h00DF; B = 16'h00FA; #100;
A = 16'h00DF; B = 16'h00FB; #100;
A = 16'h00DF; B = 16'h00FC; #100;
A = 16'h00DF; B = 16'h00FD; #100;
A = 16'h00DF; B = 16'h00FE; #100;
A = 16'h00DF; B = 16'h00FF; #100;
A = 16'h00E0; B = 16'h000; #100;
A = 16'h00E0; B = 16'h001; #100;
A = 16'h00E0; B = 16'h002; #100;
A = 16'h00E0; B = 16'h003; #100;
A = 16'h00E0; B = 16'h004; #100;
A = 16'h00E0; B = 16'h005; #100;
A = 16'h00E0; B = 16'h006; #100;
A = 16'h00E0; B = 16'h007; #100;
A = 16'h00E0; B = 16'h008; #100;
A = 16'h00E0; B = 16'h009; #100;
A = 16'h00E0; B = 16'h00A; #100;
A = 16'h00E0; B = 16'h00B; #100;
A = 16'h00E0; B = 16'h00C; #100;
A = 16'h00E0; B = 16'h00D; #100;
A = 16'h00E0; B = 16'h00E; #100;
A = 16'h00E0; B = 16'h00F; #100;
A = 16'h00E0; B = 16'h0010; #100;
A = 16'h00E0; B = 16'h0011; #100;
A = 16'h00E0; B = 16'h0012; #100;
A = 16'h00E0; B = 16'h0013; #100;
A = 16'h00E0; B = 16'h0014; #100;
A = 16'h00E0; B = 16'h0015; #100;
A = 16'h00E0; B = 16'h0016; #100;
A = 16'h00E0; B = 16'h0017; #100;
A = 16'h00E0; B = 16'h0018; #100;
A = 16'h00E0; B = 16'h0019; #100;
A = 16'h00E0; B = 16'h001A; #100;
A = 16'h00E0; B = 16'h001B; #100;
A = 16'h00E0; B = 16'h001C; #100;
A = 16'h00E0; B = 16'h001D; #100;
A = 16'h00E0; B = 16'h001E; #100;
A = 16'h00E0; B = 16'h001F; #100;
A = 16'h00E0; B = 16'h0020; #100;
A = 16'h00E0; B = 16'h0021; #100;
A = 16'h00E0; B = 16'h0022; #100;
A = 16'h00E0; B = 16'h0023; #100;
A = 16'h00E0; B = 16'h0024; #100;
A = 16'h00E0; B = 16'h0025; #100;
A = 16'h00E0; B = 16'h0026; #100;
A = 16'h00E0; B = 16'h0027; #100;
A = 16'h00E0; B = 16'h0028; #100;
A = 16'h00E0; B = 16'h0029; #100;
A = 16'h00E0; B = 16'h002A; #100;
A = 16'h00E0; B = 16'h002B; #100;
A = 16'h00E0; B = 16'h002C; #100;
A = 16'h00E0; B = 16'h002D; #100;
A = 16'h00E0; B = 16'h002E; #100;
A = 16'h00E0; B = 16'h002F; #100;
A = 16'h00E0; B = 16'h0030; #100;
A = 16'h00E0; B = 16'h0031; #100;
A = 16'h00E0; B = 16'h0032; #100;
A = 16'h00E0; B = 16'h0033; #100;
A = 16'h00E0; B = 16'h0034; #100;
A = 16'h00E0; B = 16'h0035; #100;
A = 16'h00E0; B = 16'h0036; #100;
A = 16'h00E0; B = 16'h0037; #100;
A = 16'h00E0; B = 16'h0038; #100;
A = 16'h00E0; B = 16'h0039; #100;
A = 16'h00E0; B = 16'h003A; #100;
A = 16'h00E0; B = 16'h003B; #100;
A = 16'h00E0; B = 16'h003C; #100;
A = 16'h00E0; B = 16'h003D; #100;
A = 16'h00E0; B = 16'h003E; #100;
A = 16'h00E0; B = 16'h003F; #100;
A = 16'h00E0; B = 16'h0040; #100;
A = 16'h00E0; B = 16'h0041; #100;
A = 16'h00E0; B = 16'h0042; #100;
A = 16'h00E0; B = 16'h0043; #100;
A = 16'h00E0; B = 16'h0044; #100;
A = 16'h00E0; B = 16'h0045; #100;
A = 16'h00E0; B = 16'h0046; #100;
A = 16'h00E0; B = 16'h0047; #100;
A = 16'h00E0; B = 16'h0048; #100;
A = 16'h00E0; B = 16'h0049; #100;
A = 16'h00E0; B = 16'h004A; #100;
A = 16'h00E0; B = 16'h004B; #100;
A = 16'h00E0; B = 16'h004C; #100;
A = 16'h00E0; B = 16'h004D; #100;
A = 16'h00E0; B = 16'h004E; #100;
A = 16'h00E0; B = 16'h004F; #100;
A = 16'h00E0; B = 16'h0050; #100;
A = 16'h00E0; B = 16'h0051; #100;
A = 16'h00E0; B = 16'h0052; #100;
A = 16'h00E0; B = 16'h0053; #100;
A = 16'h00E0; B = 16'h0054; #100;
A = 16'h00E0; B = 16'h0055; #100;
A = 16'h00E0; B = 16'h0056; #100;
A = 16'h00E0; B = 16'h0057; #100;
A = 16'h00E0; B = 16'h0058; #100;
A = 16'h00E0; B = 16'h0059; #100;
A = 16'h00E0; B = 16'h005A; #100;
A = 16'h00E0; B = 16'h005B; #100;
A = 16'h00E0; B = 16'h005C; #100;
A = 16'h00E0; B = 16'h005D; #100;
A = 16'h00E0; B = 16'h005E; #100;
A = 16'h00E0; B = 16'h005F; #100;
A = 16'h00E0; B = 16'h0060; #100;
A = 16'h00E0; B = 16'h0061; #100;
A = 16'h00E0; B = 16'h0062; #100;
A = 16'h00E0; B = 16'h0063; #100;
A = 16'h00E0; B = 16'h0064; #100;
A = 16'h00E0; B = 16'h0065; #100;
A = 16'h00E0; B = 16'h0066; #100;
A = 16'h00E0; B = 16'h0067; #100;
A = 16'h00E0; B = 16'h0068; #100;
A = 16'h00E0; B = 16'h0069; #100;
A = 16'h00E0; B = 16'h006A; #100;
A = 16'h00E0; B = 16'h006B; #100;
A = 16'h00E0; B = 16'h006C; #100;
A = 16'h00E0; B = 16'h006D; #100;
A = 16'h00E0; B = 16'h006E; #100;
A = 16'h00E0; B = 16'h006F; #100;
A = 16'h00E0; B = 16'h0070; #100;
A = 16'h00E0; B = 16'h0071; #100;
A = 16'h00E0; B = 16'h0072; #100;
A = 16'h00E0; B = 16'h0073; #100;
A = 16'h00E0; B = 16'h0074; #100;
A = 16'h00E0; B = 16'h0075; #100;
A = 16'h00E0; B = 16'h0076; #100;
A = 16'h00E0; B = 16'h0077; #100;
A = 16'h00E0; B = 16'h0078; #100;
A = 16'h00E0; B = 16'h0079; #100;
A = 16'h00E0; B = 16'h007A; #100;
A = 16'h00E0; B = 16'h007B; #100;
A = 16'h00E0; B = 16'h007C; #100;
A = 16'h00E0; B = 16'h007D; #100;
A = 16'h00E0; B = 16'h007E; #100;
A = 16'h00E0; B = 16'h007F; #100;
A = 16'h00E0; B = 16'h0080; #100;
A = 16'h00E0; B = 16'h0081; #100;
A = 16'h00E0; B = 16'h0082; #100;
A = 16'h00E0; B = 16'h0083; #100;
A = 16'h00E0; B = 16'h0084; #100;
A = 16'h00E0; B = 16'h0085; #100;
A = 16'h00E0; B = 16'h0086; #100;
A = 16'h00E0; B = 16'h0087; #100;
A = 16'h00E0; B = 16'h0088; #100;
A = 16'h00E0; B = 16'h0089; #100;
A = 16'h00E0; B = 16'h008A; #100;
A = 16'h00E0; B = 16'h008B; #100;
A = 16'h00E0; B = 16'h008C; #100;
A = 16'h00E0; B = 16'h008D; #100;
A = 16'h00E0; B = 16'h008E; #100;
A = 16'h00E0; B = 16'h008F; #100;
A = 16'h00E0; B = 16'h0090; #100;
A = 16'h00E0; B = 16'h0091; #100;
A = 16'h00E0; B = 16'h0092; #100;
A = 16'h00E0; B = 16'h0093; #100;
A = 16'h00E0; B = 16'h0094; #100;
A = 16'h00E0; B = 16'h0095; #100;
A = 16'h00E0; B = 16'h0096; #100;
A = 16'h00E0; B = 16'h0097; #100;
A = 16'h00E0; B = 16'h0098; #100;
A = 16'h00E0; B = 16'h0099; #100;
A = 16'h00E0; B = 16'h009A; #100;
A = 16'h00E0; B = 16'h009B; #100;
A = 16'h00E0; B = 16'h009C; #100;
A = 16'h00E0; B = 16'h009D; #100;
A = 16'h00E0; B = 16'h009E; #100;
A = 16'h00E0; B = 16'h009F; #100;
A = 16'h00E0; B = 16'h00A0; #100;
A = 16'h00E0; B = 16'h00A1; #100;
A = 16'h00E0; B = 16'h00A2; #100;
A = 16'h00E0; B = 16'h00A3; #100;
A = 16'h00E0; B = 16'h00A4; #100;
A = 16'h00E0; B = 16'h00A5; #100;
A = 16'h00E0; B = 16'h00A6; #100;
A = 16'h00E0; B = 16'h00A7; #100;
A = 16'h00E0; B = 16'h00A8; #100;
A = 16'h00E0; B = 16'h00A9; #100;
A = 16'h00E0; B = 16'h00AA; #100;
A = 16'h00E0; B = 16'h00AB; #100;
A = 16'h00E0; B = 16'h00AC; #100;
A = 16'h00E0; B = 16'h00AD; #100;
A = 16'h00E0; B = 16'h00AE; #100;
A = 16'h00E0; B = 16'h00AF; #100;
A = 16'h00E0; B = 16'h00B0; #100;
A = 16'h00E0; B = 16'h00B1; #100;
A = 16'h00E0; B = 16'h00B2; #100;
A = 16'h00E0; B = 16'h00B3; #100;
A = 16'h00E0; B = 16'h00B4; #100;
A = 16'h00E0; B = 16'h00B5; #100;
A = 16'h00E0; B = 16'h00B6; #100;
A = 16'h00E0; B = 16'h00B7; #100;
A = 16'h00E0; B = 16'h00B8; #100;
A = 16'h00E0; B = 16'h00B9; #100;
A = 16'h00E0; B = 16'h00BA; #100;
A = 16'h00E0; B = 16'h00BB; #100;
A = 16'h00E0; B = 16'h00BC; #100;
A = 16'h00E0; B = 16'h00BD; #100;
A = 16'h00E0; B = 16'h00BE; #100;
A = 16'h00E0; B = 16'h00BF; #100;
A = 16'h00E0; B = 16'h00C0; #100;
A = 16'h00E0; B = 16'h00C1; #100;
A = 16'h00E0; B = 16'h00C2; #100;
A = 16'h00E0; B = 16'h00C3; #100;
A = 16'h00E0; B = 16'h00C4; #100;
A = 16'h00E0; B = 16'h00C5; #100;
A = 16'h00E0; B = 16'h00C6; #100;
A = 16'h00E0; B = 16'h00C7; #100;
A = 16'h00E0; B = 16'h00C8; #100;
A = 16'h00E0; B = 16'h00C9; #100;
A = 16'h00E0; B = 16'h00CA; #100;
A = 16'h00E0; B = 16'h00CB; #100;
A = 16'h00E0; B = 16'h00CC; #100;
A = 16'h00E0; B = 16'h00CD; #100;
A = 16'h00E0; B = 16'h00CE; #100;
A = 16'h00E0; B = 16'h00CF; #100;
A = 16'h00E0; B = 16'h00D0; #100;
A = 16'h00E0; B = 16'h00D1; #100;
A = 16'h00E0; B = 16'h00D2; #100;
A = 16'h00E0; B = 16'h00D3; #100;
A = 16'h00E0; B = 16'h00D4; #100;
A = 16'h00E0; B = 16'h00D5; #100;
A = 16'h00E0; B = 16'h00D6; #100;
A = 16'h00E0; B = 16'h00D7; #100;
A = 16'h00E0; B = 16'h00D8; #100;
A = 16'h00E0; B = 16'h00D9; #100;
A = 16'h00E0; B = 16'h00DA; #100;
A = 16'h00E0; B = 16'h00DB; #100;
A = 16'h00E0; B = 16'h00DC; #100;
A = 16'h00E0; B = 16'h00DD; #100;
A = 16'h00E0; B = 16'h00DE; #100;
A = 16'h00E0; B = 16'h00DF; #100;
A = 16'h00E0; B = 16'h00E0; #100;
A = 16'h00E0; B = 16'h00E1; #100;
A = 16'h00E0; B = 16'h00E2; #100;
A = 16'h00E0; B = 16'h00E3; #100;
A = 16'h00E0; B = 16'h00E4; #100;
A = 16'h00E0; B = 16'h00E5; #100;
A = 16'h00E0; B = 16'h00E6; #100;
A = 16'h00E0; B = 16'h00E7; #100;
A = 16'h00E0; B = 16'h00E8; #100;
A = 16'h00E0; B = 16'h00E9; #100;
A = 16'h00E0; B = 16'h00EA; #100;
A = 16'h00E0; B = 16'h00EB; #100;
A = 16'h00E0; B = 16'h00EC; #100;
A = 16'h00E0; B = 16'h00ED; #100;
A = 16'h00E0; B = 16'h00EE; #100;
A = 16'h00E0; B = 16'h00EF; #100;
A = 16'h00E0; B = 16'h00F0; #100;
A = 16'h00E0; B = 16'h00F1; #100;
A = 16'h00E0; B = 16'h00F2; #100;
A = 16'h00E0; B = 16'h00F3; #100;
A = 16'h00E0; B = 16'h00F4; #100;
A = 16'h00E0; B = 16'h00F5; #100;
A = 16'h00E0; B = 16'h00F6; #100;
A = 16'h00E0; B = 16'h00F7; #100;
A = 16'h00E0; B = 16'h00F8; #100;
A = 16'h00E0; B = 16'h00F9; #100;
A = 16'h00E0; B = 16'h00FA; #100;
A = 16'h00E0; B = 16'h00FB; #100;
A = 16'h00E0; B = 16'h00FC; #100;
A = 16'h00E0; B = 16'h00FD; #100;
A = 16'h00E0; B = 16'h00FE; #100;
A = 16'h00E0; B = 16'h00FF; #100;
A = 16'h00E1; B = 16'h000; #100;
A = 16'h00E1; B = 16'h001; #100;
A = 16'h00E1; B = 16'h002; #100;
A = 16'h00E1; B = 16'h003; #100;
A = 16'h00E1; B = 16'h004; #100;
A = 16'h00E1; B = 16'h005; #100;
A = 16'h00E1; B = 16'h006; #100;
A = 16'h00E1; B = 16'h007; #100;
A = 16'h00E1; B = 16'h008; #100;
A = 16'h00E1; B = 16'h009; #100;
A = 16'h00E1; B = 16'h00A; #100;
A = 16'h00E1; B = 16'h00B; #100;
A = 16'h00E1; B = 16'h00C; #100;
A = 16'h00E1; B = 16'h00D; #100;
A = 16'h00E1; B = 16'h00E; #100;
A = 16'h00E1; B = 16'h00F; #100;
A = 16'h00E1; B = 16'h0010; #100;
A = 16'h00E1; B = 16'h0011; #100;
A = 16'h00E1; B = 16'h0012; #100;
A = 16'h00E1; B = 16'h0013; #100;
A = 16'h00E1; B = 16'h0014; #100;
A = 16'h00E1; B = 16'h0015; #100;
A = 16'h00E1; B = 16'h0016; #100;
A = 16'h00E1; B = 16'h0017; #100;
A = 16'h00E1; B = 16'h0018; #100;
A = 16'h00E1; B = 16'h0019; #100;
A = 16'h00E1; B = 16'h001A; #100;
A = 16'h00E1; B = 16'h001B; #100;
A = 16'h00E1; B = 16'h001C; #100;
A = 16'h00E1; B = 16'h001D; #100;
A = 16'h00E1; B = 16'h001E; #100;
A = 16'h00E1; B = 16'h001F; #100;
A = 16'h00E1; B = 16'h0020; #100;
A = 16'h00E1; B = 16'h0021; #100;
A = 16'h00E1; B = 16'h0022; #100;
A = 16'h00E1; B = 16'h0023; #100;
A = 16'h00E1; B = 16'h0024; #100;
A = 16'h00E1; B = 16'h0025; #100;
A = 16'h00E1; B = 16'h0026; #100;
A = 16'h00E1; B = 16'h0027; #100;
A = 16'h00E1; B = 16'h0028; #100;
A = 16'h00E1; B = 16'h0029; #100;
A = 16'h00E1; B = 16'h002A; #100;
A = 16'h00E1; B = 16'h002B; #100;
A = 16'h00E1; B = 16'h002C; #100;
A = 16'h00E1; B = 16'h002D; #100;
A = 16'h00E1; B = 16'h002E; #100;
A = 16'h00E1; B = 16'h002F; #100;
A = 16'h00E1; B = 16'h0030; #100;
A = 16'h00E1; B = 16'h0031; #100;
A = 16'h00E1; B = 16'h0032; #100;
A = 16'h00E1; B = 16'h0033; #100;
A = 16'h00E1; B = 16'h0034; #100;
A = 16'h00E1; B = 16'h0035; #100;
A = 16'h00E1; B = 16'h0036; #100;
A = 16'h00E1; B = 16'h0037; #100;
A = 16'h00E1; B = 16'h0038; #100;
A = 16'h00E1; B = 16'h0039; #100;
A = 16'h00E1; B = 16'h003A; #100;
A = 16'h00E1; B = 16'h003B; #100;
A = 16'h00E1; B = 16'h003C; #100;
A = 16'h00E1; B = 16'h003D; #100;
A = 16'h00E1; B = 16'h003E; #100;
A = 16'h00E1; B = 16'h003F; #100;
A = 16'h00E1; B = 16'h0040; #100;
A = 16'h00E1; B = 16'h0041; #100;
A = 16'h00E1; B = 16'h0042; #100;
A = 16'h00E1; B = 16'h0043; #100;
A = 16'h00E1; B = 16'h0044; #100;
A = 16'h00E1; B = 16'h0045; #100;
A = 16'h00E1; B = 16'h0046; #100;
A = 16'h00E1; B = 16'h0047; #100;
A = 16'h00E1; B = 16'h0048; #100;
A = 16'h00E1; B = 16'h0049; #100;
A = 16'h00E1; B = 16'h004A; #100;
A = 16'h00E1; B = 16'h004B; #100;
A = 16'h00E1; B = 16'h004C; #100;
A = 16'h00E1; B = 16'h004D; #100;
A = 16'h00E1; B = 16'h004E; #100;
A = 16'h00E1; B = 16'h004F; #100;
A = 16'h00E1; B = 16'h0050; #100;
A = 16'h00E1; B = 16'h0051; #100;
A = 16'h00E1; B = 16'h0052; #100;
A = 16'h00E1; B = 16'h0053; #100;
A = 16'h00E1; B = 16'h0054; #100;
A = 16'h00E1; B = 16'h0055; #100;
A = 16'h00E1; B = 16'h0056; #100;
A = 16'h00E1; B = 16'h0057; #100;
A = 16'h00E1; B = 16'h0058; #100;
A = 16'h00E1; B = 16'h0059; #100;
A = 16'h00E1; B = 16'h005A; #100;
A = 16'h00E1; B = 16'h005B; #100;
A = 16'h00E1; B = 16'h005C; #100;
A = 16'h00E1; B = 16'h005D; #100;
A = 16'h00E1; B = 16'h005E; #100;
A = 16'h00E1; B = 16'h005F; #100;
A = 16'h00E1; B = 16'h0060; #100;
A = 16'h00E1; B = 16'h0061; #100;
A = 16'h00E1; B = 16'h0062; #100;
A = 16'h00E1; B = 16'h0063; #100;
A = 16'h00E1; B = 16'h0064; #100;
A = 16'h00E1; B = 16'h0065; #100;
A = 16'h00E1; B = 16'h0066; #100;
A = 16'h00E1; B = 16'h0067; #100;
A = 16'h00E1; B = 16'h0068; #100;
A = 16'h00E1; B = 16'h0069; #100;
A = 16'h00E1; B = 16'h006A; #100;
A = 16'h00E1; B = 16'h006B; #100;
A = 16'h00E1; B = 16'h006C; #100;
A = 16'h00E1; B = 16'h006D; #100;
A = 16'h00E1; B = 16'h006E; #100;
A = 16'h00E1; B = 16'h006F; #100;
A = 16'h00E1; B = 16'h0070; #100;
A = 16'h00E1; B = 16'h0071; #100;
A = 16'h00E1; B = 16'h0072; #100;
A = 16'h00E1; B = 16'h0073; #100;
A = 16'h00E1; B = 16'h0074; #100;
A = 16'h00E1; B = 16'h0075; #100;
A = 16'h00E1; B = 16'h0076; #100;
A = 16'h00E1; B = 16'h0077; #100;
A = 16'h00E1; B = 16'h0078; #100;
A = 16'h00E1; B = 16'h0079; #100;
A = 16'h00E1; B = 16'h007A; #100;
A = 16'h00E1; B = 16'h007B; #100;
A = 16'h00E1; B = 16'h007C; #100;
A = 16'h00E1; B = 16'h007D; #100;
A = 16'h00E1; B = 16'h007E; #100;
A = 16'h00E1; B = 16'h007F; #100;
A = 16'h00E1; B = 16'h0080; #100;
A = 16'h00E1; B = 16'h0081; #100;
A = 16'h00E1; B = 16'h0082; #100;
A = 16'h00E1; B = 16'h0083; #100;
A = 16'h00E1; B = 16'h0084; #100;
A = 16'h00E1; B = 16'h0085; #100;
A = 16'h00E1; B = 16'h0086; #100;
A = 16'h00E1; B = 16'h0087; #100;
A = 16'h00E1; B = 16'h0088; #100;
A = 16'h00E1; B = 16'h0089; #100;
A = 16'h00E1; B = 16'h008A; #100;
A = 16'h00E1; B = 16'h008B; #100;
A = 16'h00E1; B = 16'h008C; #100;
A = 16'h00E1; B = 16'h008D; #100;
A = 16'h00E1; B = 16'h008E; #100;
A = 16'h00E1; B = 16'h008F; #100;
A = 16'h00E1; B = 16'h0090; #100;
A = 16'h00E1; B = 16'h0091; #100;
A = 16'h00E1; B = 16'h0092; #100;
A = 16'h00E1; B = 16'h0093; #100;
A = 16'h00E1; B = 16'h0094; #100;
A = 16'h00E1; B = 16'h0095; #100;
A = 16'h00E1; B = 16'h0096; #100;
A = 16'h00E1; B = 16'h0097; #100;
A = 16'h00E1; B = 16'h0098; #100;
A = 16'h00E1; B = 16'h0099; #100;
A = 16'h00E1; B = 16'h009A; #100;
A = 16'h00E1; B = 16'h009B; #100;
A = 16'h00E1; B = 16'h009C; #100;
A = 16'h00E1; B = 16'h009D; #100;
A = 16'h00E1; B = 16'h009E; #100;
A = 16'h00E1; B = 16'h009F; #100;
A = 16'h00E1; B = 16'h00A0; #100;
A = 16'h00E1; B = 16'h00A1; #100;
A = 16'h00E1; B = 16'h00A2; #100;
A = 16'h00E1; B = 16'h00A3; #100;
A = 16'h00E1; B = 16'h00A4; #100;
A = 16'h00E1; B = 16'h00A5; #100;
A = 16'h00E1; B = 16'h00A6; #100;
A = 16'h00E1; B = 16'h00A7; #100;
A = 16'h00E1; B = 16'h00A8; #100;
A = 16'h00E1; B = 16'h00A9; #100;
A = 16'h00E1; B = 16'h00AA; #100;
A = 16'h00E1; B = 16'h00AB; #100;
A = 16'h00E1; B = 16'h00AC; #100;
A = 16'h00E1; B = 16'h00AD; #100;
A = 16'h00E1; B = 16'h00AE; #100;
A = 16'h00E1; B = 16'h00AF; #100;
A = 16'h00E1; B = 16'h00B0; #100;
A = 16'h00E1; B = 16'h00B1; #100;
A = 16'h00E1; B = 16'h00B2; #100;
A = 16'h00E1; B = 16'h00B3; #100;
A = 16'h00E1; B = 16'h00B4; #100;
A = 16'h00E1; B = 16'h00B5; #100;
A = 16'h00E1; B = 16'h00B6; #100;
A = 16'h00E1; B = 16'h00B7; #100;
A = 16'h00E1; B = 16'h00B8; #100;
A = 16'h00E1; B = 16'h00B9; #100;
A = 16'h00E1; B = 16'h00BA; #100;
A = 16'h00E1; B = 16'h00BB; #100;
A = 16'h00E1; B = 16'h00BC; #100;
A = 16'h00E1; B = 16'h00BD; #100;
A = 16'h00E1; B = 16'h00BE; #100;
A = 16'h00E1; B = 16'h00BF; #100;
A = 16'h00E1; B = 16'h00C0; #100;
A = 16'h00E1; B = 16'h00C1; #100;
A = 16'h00E1; B = 16'h00C2; #100;
A = 16'h00E1; B = 16'h00C3; #100;
A = 16'h00E1; B = 16'h00C4; #100;
A = 16'h00E1; B = 16'h00C5; #100;
A = 16'h00E1; B = 16'h00C6; #100;
A = 16'h00E1; B = 16'h00C7; #100;
A = 16'h00E1; B = 16'h00C8; #100;
A = 16'h00E1; B = 16'h00C9; #100;
A = 16'h00E1; B = 16'h00CA; #100;
A = 16'h00E1; B = 16'h00CB; #100;
A = 16'h00E1; B = 16'h00CC; #100;
A = 16'h00E1; B = 16'h00CD; #100;
A = 16'h00E1; B = 16'h00CE; #100;
A = 16'h00E1; B = 16'h00CF; #100;
A = 16'h00E1; B = 16'h00D0; #100;
A = 16'h00E1; B = 16'h00D1; #100;
A = 16'h00E1; B = 16'h00D2; #100;
A = 16'h00E1; B = 16'h00D3; #100;
A = 16'h00E1; B = 16'h00D4; #100;
A = 16'h00E1; B = 16'h00D5; #100;
A = 16'h00E1; B = 16'h00D6; #100;
A = 16'h00E1; B = 16'h00D7; #100;
A = 16'h00E1; B = 16'h00D8; #100;
A = 16'h00E1; B = 16'h00D9; #100;
A = 16'h00E1; B = 16'h00DA; #100;
A = 16'h00E1; B = 16'h00DB; #100;
A = 16'h00E1; B = 16'h00DC; #100;
A = 16'h00E1; B = 16'h00DD; #100;
A = 16'h00E1; B = 16'h00DE; #100;
A = 16'h00E1; B = 16'h00DF; #100;
A = 16'h00E1; B = 16'h00E0; #100;
A = 16'h00E1; B = 16'h00E1; #100;
A = 16'h00E1; B = 16'h00E2; #100;
A = 16'h00E1; B = 16'h00E3; #100;
A = 16'h00E1; B = 16'h00E4; #100;
A = 16'h00E1; B = 16'h00E5; #100;
A = 16'h00E1; B = 16'h00E6; #100;
A = 16'h00E1; B = 16'h00E7; #100;
A = 16'h00E1; B = 16'h00E8; #100;
A = 16'h00E1; B = 16'h00E9; #100;
A = 16'h00E1; B = 16'h00EA; #100;
A = 16'h00E1; B = 16'h00EB; #100;
A = 16'h00E1; B = 16'h00EC; #100;
A = 16'h00E1; B = 16'h00ED; #100;
A = 16'h00E1; B = 16'h00EE; #100;
A = 16'h00E1; B = 16'h00EF; #100;
A = 16'h00E1; B = 16'h00F0; #100;
A = 16'h00E1; B = 16'h00F1; #100;
A = 16'h00E1; B = 16'h00F2; #100;
A = 16'h00E1; B = 16'h00F3; #100;
A = 16'h00E1; B = 16'h00F4; #100;
A = 16'h00E1; B = 16'h00F5; #100;
A = 16'h00E1; B = 16'h00F6; #100;
A = 16'h00E1; B = 16'h00F7; #100;
A = 16'h00E1; B = 16'h00F8; #100;
A = 16'h00E1; B = 16'h00F9; #100;
A = 16'h00E1; B = 16'h00FA; #100;
A = 16'h00E1; B = 16'h00FB; #100;
A = 16'h00E1; B = 16'h00FC; #100;
A = 16'h00E1; B = 16'h00FD; #100;
A = 16'h00E1; B = 16'h00FE; #100;
A = 16'h00E1; B = 16'h00FF; #100;
A = 16'h00E2; B = 16'h000; #100;
A = 16'h00E2; B = 16'h001; #100;
A = 16'h00E2; B = 16'h002; #100;
A = 16'h00E2; B = 16'h003; #100;
A = 16'h00E2; B = 16'h004; #100;
A = 16'h00E2; B = 16'h005; #100;
A = 16'h00E2; B = 16'h006; #100;
A = 16'h00E2; B = 16'h007; #100;
A = 16'h00E2; B = 16'h008; #100;
A = 16'h00E2; B = 16'h009; #100;
A = 16'h00E2; B = 16'h00A; #100;
A = 16'h00E2; B = 16'h00B; #100;
A = 16'h00E2; B = 16'h00C; #100;
A = 16'h00E2; B = 16'h00D; #100;
A = 16'h00E2; B = 16'h00E; #100;
A = 16'h00E2; B = 16'h00F; #100;
A = 16'h00E2; B = 16'h0010; #100;
A = 16'h00E2; B = 16'h0011; #100;
A = 16'h00E2; B = 16'h0012; #100;
A = 16'h00E2; B = 16'h0013; #100;
A = 16'h00E2; B = 16'h0014; #100;
A = 16'h00E2; B = 16'h0015; #100;
A = 16'h00E2; B = 16'h0016; #100;
A = 16'h00E2; B = 16'h0017; #100;
A = 16'h00E2; B = 16'h0018; #100;
A = 16'h00E2; B = 16'h0019; #100;
A = 16'h00E2; B = 16'h001A; #100;
A = 16'h00E2; B = 16'h001B; #100;
A = 16'h00E2; B = 16'h001C; #100;
A = 16'h00E2; B = 16'h001D; #100;
A = 16'h00E2; B = 16'h001E; #100;
A = 16'h00E2; B = 16'h001F; #100;
A = 16'h00E2; B = 16'h0020; #100;
A = 16'h00E2; B = 16'h0021; #100;
A = 16'h00E2; B = 16'h0022; #100;
A = 16'h00E2; B = 16'h0023; #100;
A = 16'h00E2; B = 16'h0024; #100;
A = 16'h00E2; B = 16'h0025; #100;
A = 16'h00E2; B = 16'h0026; #100;
A = 16'h00E2; B = 16'h0027; #100;
A = 16'h00E2; B = 16'h0028; #100;
A = 16'h00E2; B = 16'h0029; #100;
A = 16'h00E2; B = 16'h002A; #100;
A = 16'h00E2; B = 16'h002B; #100;
A = 16'h00E2; B = 16'h002C; #100;
A = 16'h00E2; B = 16'h002D; #100;
A = 16'h00E2; B = 16'h002E; #100;
A = 16'h00E2; B = 16'h002F; #100;
A = 16'h00E2; B = 16'h0030; #100;
A = 16'h00E2; B = 16'h0031; #100;
A = 16'h00E2; B = 16'h0032; #100;
A = 16'h00E2; B = 16'h0033; #100;
A = 16'h00E2; B = 16'h0034; #100;
A = 16'h00E2; B = 16'h0035; #100;
A = 16'h00E2; B = 16'h0036; #100;
A = 16'h00E2; B = 16'h0037; #100;
A = 16'h00E2; B = 16'h0038; #100;
A = 16'h00E2; B = 16'h0039; #100;
A = 16'h00E2; B = 16'h003A; #100;
A = 16'h00E2; B = 16'h003B; #100;
A = 16'h00E2; B = 16'h003C; #100;
A = 16'h00E2; B = 16'h003D; #100;
A = 16'h00E2; B = 16'h003E; #100;
A = 16'h00E2; B = 16'h003F; #100;
A = 16'h00E2; B = 16'h0040; #100;
A = 16'h00E2; B = 16'h0041; #100;
A = 16'h00E2; B = 16'h0042; #100;
A = 16'h00E2; B = 16'h0043; #100;
A = 16'h00E2; B = 16'h0044; #100;
A = 16'h00E2; B = 16'h0045; #100;
A = 16'h00E2; B = 16'h0046; #100;
A = 16'h00E2; B = 16'h0047; #100;
A = 16'h00E2; B = 16'h0048; #100;
A = 16'h00E2; B = 16'h0049; #100;
A = 16'h00E2; B = 16'h004A; #100;
A = 16'h00E2; B = 16'h004B; #100;
A = 16'h00E2; B = 16'h004C; #100;
A = 16'h00E2; B = 16'h004D; #100;
A = 16'h00E2; B = 16'h004E; #100;
A = 16'h00E2; B = 16'h004F; #100;
A = 16'h00E2; B = 16'h0050; #100;
A = 16'h00E2; B = 16'h0051; #100;
A = 16'h00E2; B = 16'h0052; #100;
A = 16'h00E2; B = 16'h0053; #100;
A = 16'h00E2; B = 16'h0054; #100;
A = 16'h00E2; B = 16'h0055; #100;
A = 16'h00E2; B = 16'h0056; #100;
A = 16'h00E2; B = 16'h0057; #100;
A = 16'h00E2; B = 16'h0058; #100;
A = 16'h00E2; B = 16'h0059; #100;
A = 16'h00E2; B = 16'h005A; #100;
A = 16'h00E2; B = 16'h005B; #100;
A = 16'h00E2; B = 16'h005C; #100;
A = 16'h00E2; B = 16'h005D; #100;
A = 16'h00E2; B = 16'h005E; #100;
A = 16'h00E2; B = 16'h005F; #100;
A = 16'h00E2; B = 16'h0060; #100;
A = 16'h00E2; B = 16'h0061; #100;
A = 16'h00E2; B = 16'h0062; #100;
A = 16'h00E2; B = 16'h0063; #100;
A = 16'h00E2; B = 16'h0064; #100;
A = 16'h00E2; B = 16'h0065; #100;
A = 16'h00E2; B = 16'h0066; #100;
A = 16'h00E2; B = 16'h0067; #100;
A = 16'h00E2; B = 16'h0068; #100;
A = 16'h00E2; B = 16'h0069; #100;
A = 16'h00E2; B = 16'h006A; #100;
A = 16'h00E2; B = 16'h006B; #100;
A = 16'h00E2; B = 16'h006C; #100;
A = 16'h00E2; B = 16'h006D; #100;
A = 16'h00E2; B = 16'h006E; #100;
A = 16'h00E2; B = 16'h006F; #100;
A = 16'h00E2; B = 16'h0070; #100;
A = 16'h00E2; B = 16'h0071; #100;
A = 16'h00E2; B = 16'h0072; #100;
A = 16'h00E2; B = 16'h0073; #100;
A = 16'h00E2; B = 16'h0074; #100;
A = 16'h00E2; B = 16'h0075; #100;
A = 16'h00E2; B = 16'h0076; #100;
A = 16'h00E2; B = 16'h0077; #100;
A = 16'h00E2; B = 16'h0078; #100;
A = 16'h00E2; B = 16'h0079; #100;
A = 16'h00E2; B = 16'h007A; #100;
A = 16'h00E2; B = 16'h007B; #100;
A = 16'h00E2; B = 16'h007C; #100;
A = 16'h00E2; B = 16'h007D; #100;
A = 16'h00E2; B = 16'h007E; #100;
A = 16'h00E2; B = 16'h007F; #100;
A = 16'h00E2; B = 16'h0080; #100;
A = 16'h00E2; B = 16'h0081; #100;
A = 16'h00E2; B = 16'h0082; #100;
A = 16'h00E2; B = 16'h0083; #100;
A = 16'h00E2; B = 16'h0084; #100;
A = 16'h00E2; B = 16'h0085; #100;
A = 16'h00E2; B = 16'h0086; #100;
A = 16'h00E2; B = 16'h0087; #100;
A = 16'h00E2; B = 16'h0088; #100;
A = 16'h00E2; B = 16'h0089; #100;
A = 16'h00E2; B = 16'h008A; #100;
A = 16'h00E2; B = 16'h008B; #100;
A = 16'h00E2; B = 16'h008C; #100;
A = 16'h00E2; B = 16'h008D; #100;
A = 16'h00E2; B = 16'h008E; #100;
A = 16'h00E2; B = 16'h008F; #100;
A = 16'h00E2; B = 16'h0090; #100;
A = 16'h00E2; B = 16'h0091; #100;
A = 16'h00E2; B = 16'h0092; #100;
A = 16'h00E2; B = 16'h0093; #100;
A = 16'h00E2; B = 16'h0094; #100;
A = 16'h00E2; B = 16'h0095; #100;
A = 16'h00E2; B = 16'h0096; #100;
A = 16'h00E2; B = 16'h0097; #100;
A = 16'h00E2; B = 16'h0098; #100;
A = 16'h00E2; B = 16'h0099; #100;
A = 16'h00E2; B = 16'h009A; #100;
A = 16'h00E2; B = 16'h009B; #100;
A = 16'h00E2; B = 16'h009C; #100;
A = 16'h00E2; B = 16'h009D; #100;
A = 16'h00E2; B = 16'h009E; #100;
A = 16'h00E2; B = 16'h009F; #100;
A = 16'h00E2; B = 16'h00A0; #100;
A = 16'h00E2; B = 16'h00A1; #100;
A = 16'h00E2; B = 16'h00A2; #100;
A = 16'h00E2; B = 16'h00A3; #100;
A = 16'h00E2; B = 16'h00A4; #100;
A = 16'h00E2; B = 16'h00A5; #100;
A = 16'h00E2; B = 16'h00A6; #100;
A = 16'h00E2; B = 16'h00A7; #100;
A = 16'h00E2; B = 16'h00A8; #100;
A = 16'h00E2; B = 16'h00A9; #100;
A = 16'h00E2; B = 16'h00AA; #100;
A = 16'h00E2; B = 16'h00AB; #100;
A = 16'h00E2; B = 16'h00AC; #100;
A = 16'h00E2; B = 16'h00AD; #100;
A = 16'h00E2; B = 16'h00AE; #100;
A = 16'h00E2; B = 16'h00AF; #100;
A = 16'h00E2; B = 16'h00B0; #100;
A = 16'h00E2; B = 16'h00B1; #100;
A = 16'h00E2; B = 16'h00B2; #100;
A = 16'h00E2; B = 16'h00B3; #100;
A = 16'h00E2; B = 16'h00B4; #100;
A = 16'h00E2; B = 16'h00B5; #100;
A = 16'h00E2; B = 16'h00B6; #100;
A = 16'h00E2; B = 16'h00B7; #100;
A = 16'h00E2; B = 16'h00B8; #100;
A = 16'h00E2; B = 16'h00B9; #100;
A = 16'h00E2; B = 16'h00BA; #100;
A = 16'h00E2; B = 16'h00BB; #100;
A = 16'h00E2; B = 16'h00BC; #100;
A = 16'h00E2; B = 16'h00BD; #100;
A = 16'h00E2; B = 16'h00BE; #100;
A = 16'h00E2; B = 16'h00BF; #100;
A = 16'h00E2; B = 16'h00C0; #100;
A = 16'h00E2; B = 16'h00C1; #100;
A = 16'h00E2; B = 16'h00C2; #100;
A = 16'h00E2; B = 16'h00C3; #100;
A = 16'h00E2; B = 16'h00C4; #100;
A = 16'h00E2; B = 16'h00C5; #100;
A = 16'h00E2; B = 16'h00C6; #100;
A = 16'h00E2; B = 16'h00C7; #100;
A = 16'h00E2; B = 16'h00C8; #100;
A = 16'h00E2; B = 16'h00C9; #100;
A = 16'h00E2; B = 16'h00CA; #100;
A = 16'h00E2; B = 16'h00CB; #100;
A = 16'h00E2; B = 16'h00CC; #100;
A = 16'h00E2; B = 16'h00CD; #100;
A = 16'h00E2; B = 16'h00CE; #100;
A = 16'h00E2; B = 16'h00CF; #100;
A = 16'h00E2; B = 16'h00D0; #100;
A = 16'h00E2; B = 16'h00D1; #100;
A = 16'h00E2; B = 16'h00D2; #100;
A = 16'h00E2; B = 16'h00D3; #100;
A = 16'h00E2; B = 16'h00D4; #100;
A = 16'h00E2; B = 16'h00D5; #100;
A = 16'h00E2; B = 16'h00D6; #100;
A = 16'h00E2; B = 16'h00D7; #100;
A = 16'h00E2; B = 16'h00D8; #100;
A = 16'h00E2; B = 16'h00D9; #100;
A = 16'h00E2; B = 16'h00DA; #100;
A = 16'h00E2; B = 16'h00DB; #100;
A = 16'h00E2; B = 16'h00DC; #100;
A = 16'h00E2; B = 16'h00DD; #100;
A = 16'h00E2; B = 16'h00DE; #100;
A = 16'h00E2; B = 16'h00DF; #100;
A = 16'h00E2; B = 16'h00E0; #100;
A = 16'h00E2; B = 16'h00E1; #100;
A = 16'h00E2; B = 16'h00E2; #100;
A = 16'h00E2; B = 16'h00E3; #100;
A = 16'h00E2; B = 16'h00E4; #100;
A = 16'h00E2; B = 16'h00E5; #100;
A = 16'h00E2; B = 16'h00E6; #100;
A = 16'h00E2; B = 16'h00E7; #100;
A = 16'h00E2; B = 16'h00E8; #100;
A = 16'h00E2; B = 16'h00E9; #100;
A = 16'h00E2; B = 16'h00EA; #100;
A = 16'h00E2; B = 16'h00EB; #100;
A = 16'h00E2; B = 16'h00EC; #100;
A = 16'h00E2; B = 16'h00ED; #100;
A = 16'h00E2; B = 16'h00EE; #100;
A = 16'h00E2; B = 16'h00EF; #100;
A = 16'h00E2; B = 16'h00F0; #100;
A = 16'h00E2; B = 16'h00F1; #100;
A = 16'h00E2; B = 16'h00F2; #100;
A = 16'h00E2; B = 16'h00F3; #100;
A = 16'h00E2; B = 16'h00F4; #100;
A = 16'h00E2; B = 16'h00F5; #100;
A = 16'h00E2; B = 16'h00F6; #100;
A = 16'h00E2; B = 16'h00F7; #100;
A = 16'h00E2; B = 16'h00F8; #100;
A = 16'h00E2; B = 16'h00F9; #100;
A = 16'h00E2; B = 16'h00FA; #100;
A = 16'h00E2; B = 16'h00FB; #100;
A = 16'h00E2; B = 16'h00FC; #100;
A = 16'h00E2; B = 16'h00FD; #100;
A = 16'h00E2; B = 16'h00FE; #100;
A = 16'h00E2; B = 16'h00FF; #100;
A = 16'h00E3; B = 16'h000; #100;
A = 16'h00E3; B = 16'h001; #100;
A = 16'h00E3; B = 16'h002; #100;
A = 16'h00E3; B = 16'h003; #100;
A = 16'h00E3; B = 16'h004; #100;
A = 16'h00E3; B = 16'h005; #100;
A = 16'h00E3; B = 16'h006; #100;
A = 16'h00E3; B = 16'h007; #100;
A = 16'h00E3; B = 16'h008; #100;
A = 16'h00E3; B = 16'h009; #100;
A = 16'h00E3; B = 16'h00A; #100;
A = 16'h00E3; B = 16'h00B; #100;
A = 16'h00E3; B = 16'h00C; #100;
A = 16'h00E3; B = 16'h00D; #100;
A = 16'h00E3; B = 16'h00E; #100;
A = 16'h00E3; B = 16'h00F; #100;
A = 16'h00E3; B = 16'h0010; #100;
A = 16'h00E3; B = 16'h0011; #100;
A = 16'h00E3; B = 16'h0012; #100;
A = 16'h00E3; B = 16'h0013; #100;
A = 16'h00E3; B = 16'h0014; #100;
A = 16'h00E3; B = 16'h0015; #100;
A = 16'h00E3; B = 16'h0016; #100;
A = 16'h00E3; B = 16'h0017; #100;
A = 16'h00E3; B = 16'h0018; #100;
A = 16'h00E3; B = 16'h0019; #100;
A = 16'h00E3; B = 16'h001A; #100;
A = 16'h00E3; B = 16'h001B; #100;
A = 16'h00E3; B = 16'h001C; #100;
A = 16'h00E3; B = 16'h001D; #100;
A = 16'h00E3; B = 16'h001E; #100;
A = 16'h00E3; B = 16'h001F; #100;
A = 16'h00E3; B = 16'h0020; #100;
A = 16'h00E3; B = 16'h0021; #100;
A = 16'h00E3; B = 16'h0022; #100;
A = 16'h00E3; B = 16'h0023; #100;
A = 16'h00E3; B = 16'h0024; #100;
A = 16'h00E3; B = 16'h0025; #100;
A = 16'h00E3; B = 16'h0026; #100;
A = 16'h00E3; B = 16'h0027; #100;
A = 16'h00E3; B = 16'h0028; #100;
A = 16'h00E3; B = 16'h0029; #100;
A = 16'h00E3; B = 16'h002A; #100;
A = 16'h00E3; B = 16'h002B; #100;
A = 16'h00E3; B = 16'h002C; #100;
A = 16'h00E3; B = 16'h002D; #100;
A = 16'h00E3; B = 16'h002E; #100;
A = 16'h00E3; B = 16'h002F; #100;
A = 16'h00E3; B = 16'h0030; #100;
A = 16'h00E3; B = 16'h0031; #100;
A = 16'h00E3; B = 16'h0032; #100;
A = 16'h00E3; B = 16'h0033; #100;
A = 16'h00E3; B = 16'h0034; #100;
A = 16'h00E3; B = 16'h0035; #100;
A = 16'h00E3; B = 16'h0036; #100;
A = 16'h00E3; B = 16'h0037; #100;
A = 16'h00E3; B = 16'h0038; #100;
A = 16'h00E3; B = 16'h0039; #100;
A = 16'h00E3; B = 16'h003A; #100;
A = 16'h00E3; B = 16'h003B; #100;
A = 16'h00E3; B = 16'h003C; #100;
A = 16'h00E3; B = 16'h003D; #100;
A = 16'h00E3; B = 16'h003E; #100;
A = 16'h00E3; B = 16'h003F; #100;
A = 16'h00E3; B = 16'h0040; #100;
A = 16'h00E3; B = 16'h0041; #100;
A = 16'h00E3; B = 16'h0042; #100;
A = 16'h00E3; B = 16'h0043; #100;
A = 16'h00E3; B = 16'h0044; #100;
A = 16'h00E3; B = 16'h0045; #100;
A = 16'h00E3; B = 16'h0046; #100;
A = 16'h00E3; B = 16'h0047; #100;
A = 16'h00E3; B = 16'h0048; #100;
A = 16'h00E3; B = 16'h0049; #100;
A = 16'h00E3; B = 16'h004A; #100;
A = 16'h00E3; B = 16'h004B; #100;
A = 16'h00E3; B = 16'h004C; #100;
A = 16'h00E3; B = 16'h004D; #100;
A = 16'h00E3; B = 16'h004E; #100;
A = 16'h00E3; B = 16'h004F; #100;
A = 16'h00E3; B = 16'h0050; #100;
A = 16'h00E3; B = 16'h0051; #100;
A = 16'h00E3; B = 16'h0052; #100;
A = 16'h00E3; B = 16'h0053; #100;
A = 16'h00E3; B = 16'h0054; #100;
A = 16'h00E3; B = 16'h0055; #100;
A = 16'h00E3; B = 16'h0056; #100;
A = 16'h00E3; B = 16'h0057; #100;
A = 16'h00E3; B = 16'h0058; #100;
A = 16'h00E3; B = 16'h0059; #100;
A = 16'h00E3; B = 16'h005A; #100;
A = 16'h00E3; B = 16'h005B; #100;
A = 16'h00E3; B = 16'h005C; #100;
A = 16'h00E3; B = 16'h005D; #100;
A = 16'h00E3; B = 16'h005E; #100;
A = 16'h00E3; B = 16'h005F; #100;
A = 16'h00E3; B = 16'h0060; #100;
A = 16'h00E3; B = 16'h0061; #100;
A = 16'h00E3; B = 16'h0062; #100;
A = 16'h00E3; B = 16'h0063; #100;
A = 16'h00E3; B = 16'h0064; #100;
A = 16'h00E3; B = 16'h0065; #100;
A = 16'h00E3; B = 16'h0066; #100;
A = 16'h00E3; B = 16'h0067; #100;
A = 16'h00E3; B = 16'h0068; #100;
A = 16'h00E3; B = 16'h0069; #100;
A = 16'h00E3; B = 16'h006A; #100;
A = 16'h00E3; B = 16'h006B; #100;
A = 16'h00E3; B = 16'h006C; #100;
A = 16'h00E3; B = 16'h006D; #100;
A = 16'h00E3; B = 16'h006E; #100;
A = 16'h00E3; B = 16'h006F; #100;
A = 16'h00E3; B = 16'h0070; #100;
A = 16'h00E3; B = 16'h0071; #100;
A = 16'h00E3; B = 16'h0072; #100;
A = 16'h00E3; B = 16'h0073; #100;
A = 16'h00E3; B = 16'h0074; #100;
A = 16'h00E3; B = 16'h0075; #100;
A = 16'h00E3; B = 16'h0076; #100;
A = 16'h00E3; B = 16'h0077; #100;
A = 16'h00E3; B = 16'h0078; #100;
A = 16'h00E3; B = 16'h0079; #100;
A = 16'h00E3; B = 16'h007A; #100;
A = 16'h00E3; B = 16'h007B; #100;
A = 16'h00E3; B = 16'h007C; #100;
A = 16'h00E3; B = 16'h007D; #100;
A = 16'h00E3; B = 16'h007E; #100;
A = 16'h00E3; B = 16'h007F; #100;
A = 16'h00E3; B = 16'h0080; #100;
A = 16'h00E3; B = 16'h0081; #100;
A = 16'h00E3; B = 16'h0082; #100;
A = 16'h00E3; B = 16'h0083; #100;
A = 16'h00E3; B = 16'h0084; #100;
A = 16'h00E3; B = 16'h0085; #100;
A = 16'h00E3; B = 16'h0086; #100;
A = 16'h00E3; B = 16'h0087; #100;
A = 16'h00E3; B = 16'h0088; #100;
A = 16'h00E3; B = 16'h0089; #100;
A = 16'h00E3; B = 16'h008A; #100;
A = 16'h00E3; B = 16'h008B; #100;
A = 16'h00E3; B = 16'h008C; #100;
A = 16'h00E3; B = 16'h008D; #100;
A = 16'h00E3; B = 16'h008E; #100;
A = 16'h00E3; B = 16'h008F; #100;
A = 16'h00E3; B = 16'h0090; #100;
A = 16'h00E3; B = 16'h0091; #100;
A = 16'h00E3; B = 16'h0092; #100;
A = 16'h00E3; B = 16'h0093; #100;
A = 16'h00E3; B = 16'h0094; #100;
A = 16'h00E3; B = 16'h0095; #100;
A = 16'h00E3; B = 16'h0096; #100;
A = 16'h00E3; B = 16'h0097; #100;
A = 16'h00E3; B = 16'h0098; #100;
A = 16'h00E3; B = 16'h0099; #100;
A = 16'h00E3; B = 16'h009A; #100;
A = 16'h00E3; B = 16'h009B; #100;
A = 16'h00E3; B = 16'h009C; #100;
A = 16'h00E3; B = 16'h009D; #100;
A = 16'h00E3; B = 16'h009E; #100;
A = 16'h00E3; B = 16'h009F; #100;
A = 16'h00E3; B = 16'h00A0; #100;
A = 16'h00E3; B = 16'h00A1; #100;
A = 16'h00E3; B = 16'h00A2; #100;
A = 16'h00E3; B = 16'h00A3; #100;
A = 16'h00E3; B = 16'h00A4; #100;
A = 16'h00E3; B = 16'h00A5; #100;
A = 16'h00E3; B = 16'h00A6; #100;
A = 16'h00E3; B = 16'h00A7; #100;
A = 16'h00E3; B = 16'h00A8; #100;
A = 16'h00E3; B = 16'h00A9; #100;
A = 16'h00E3; B = 16'h00AA; #100;
A = 16'h00E3; B = 16'h00AB; #100;
A = 16'h00E3; B = 16'h00AC; #100;
A = 16'h00E3; B = 16'h00AD; #100;
A = 16'h00E3; B = 16'h00AE; #100;
A = 16'h00E3; B = 16'h00AF; #100;
A = 16'h00E3; B = 16'h00B0; #100;
A = 16'h00E3; B = 16'h00B1; #100;
A = 16'h00E3; B = 16'h00B2; #100;
A = 16'h00E3; B = 16'h00B3; #100;
A = 16'h00E3; B = 16'h00B4; #100;
A = 16'h00E3; B = 16'h00B5; #100;
A = 16'h00E3; B = 16'h00B6; #100;
A = 16'h00E3; B = 16'h00B7; #100;
A = 16'h00E3; B = 16'h00B8; #100;
A = 16'h00E3; B = 16'h00B9; #100;
A = 16'h00E3; B = 16'h00BA; #100;
A = 16'h00E3; B = 16'h00BB; #100;
A = 16'h00E3; B = 16'h00BC; #100;
A = 16'h00E3; B = 16'h00BD; #100;
A = 16'h00E3; B = 16'h00BE; #100;
A = 16'h00E3; B = 16'h00BF; #100;
A = 16'h00E3; B = 16'h00C0; #100;
A = 16'h00E3; B = 16'h00C1; #100;
A = 16'h00E3; B = 16'h00C2; #100;
A = 16'h00E3; B = 16'h00C3; #100;
A = 16'h00E3; B = 16'h00C4; #100;
A = 16'h00E3; B = 16'h00C5; #100;
A = 16'h00E3; B = 16'h00C6; #100;
A = 16'h00E3; B = 16'h00C7; #100;
A = 16'h00E3; B = 16'h00C8; #100;
A = 16'h00E3; B = 16'h00C9; #100;
A = 16'h00E3; B = 16'h00CA; #100;
A = 16'h00E3; B = 16'h00CB; #100;
A = 16'h00E3; B = 16'h00CC; #100;
A = 16'h00E3; B = 16'h00CD; #100;
A = 16'h00E3; B = 16'h00CE; #100;
A = 16'h00E3; B = 16'h00CF; #100;
A = 16'h00E3; B = 16'h00D0; #100;
A = 16'h00E3; B = 16'h00D1; #100;
A = 16'h00E3; B = 16'h00D2; #100;
A = 16'h00E3; B = 16'h00D3; #100;
A = 16'h00E3; B = 16'h00D4; #100;
A = 16'h00E3; B = 16'h00D5; #100;
A = 16'h00E3; B = 16'h00D6; #100;
A = 16'h00E3; B = 16'h00D7; #100;
A = 16'h00E3; B = 16'h00D8; #100;
A = 16'h00E3; B = 16'h00D9; #100;
A = 16'h00E3; B = 16'h00DA; #100;
A = 16'h00E3; B = 16'h00DB; #100;
A = 16'h00E3; B = 16'h00DC; #100;
A = 16'h00E3; B = 16'h00DD; #100;
A = 16'h00E3; B = 16'h00DE; #100;
A = 16'h00E3; B = 16'h00DF; #100;
A = 16'h00E3; B = 16'h00E0; #100;
A = 16'h00E3; B = 16'h00E1; #100;
A = 16'h00E3; B = 16'h00E2; #100;
A = 16'h00E3; B = 16'h00E3; #100;
A = 16'h00E3; B = 16'h00E4; #100;
A = 16'h00E3; B = 16'h00E5; #100;
A = 16'h00E3; B = 16'h00E6; #100;
A = 16'h00E3; B = 16'h00E7; #100;
A = 16'h00E3; B = 16'h00E8; #100;
A = 16'h00E3; B = 16'h00E9; #100;
A = 16'h00E3; B = 16'h00EA; #100;
A = 16'h00E3; B = 16'h00EB; #100;
A = 16'h00E3; B = 16'h00EC; #100;
A = 16'h00E3; B = 16'h00ED; #100;
A = 16'h00E3; B = 16'h00EE; #100;
A = 16'h00E3; B = 16'h00EF; #100;
A = 16'h00E3; B = 16'h00F0; #100;
A = 16'h00E3; B = 16'h00F1; #100;
A = 16'h00E3; B = 16'h00F2; #100;
A = 16'h00E3; B = 16'h00F3; #100;
A = 16'h00E3; B = 16'h00F4; #100;
A = 16'h00E3; B = 16'h00F5; #100;
A = 16'h00E3; B = 16'h00F6; #100;
A = 16'h00E3; B = 16'h00F7; #100;
A = 16'h00E3; B = 16'h00F8; #100;
A = 16'h00E3; B = 16'h00F9; #100;
A = 16'h00E3; B = 16'h00FA; #100;
A = 16'h00E3; B = 16'h00FB; #100;
A = 16'h00E3; B = 16'h00FC; #100;
A = 16'h00E3; B = 16'h00FD; #100;
A = 16'h00E3; B = 16'h00FE; #100;
A = 16'h00E3; B = 16'h00FF; #100;
A = 16'h00E4; B = 16'h000; #100;
A = 16'h00E4; B = 16'h001; #100;
A = 16'h00E4; B = 16'h002; #100;
A = 16'h00E4; B = 16'h003; #100;
A = 16'h00E4; B = 16'h004; #100;
A = 16'h00E4; B = 16'h005; #100;
A = 16'h00E4; B = 16'h006; #100;
A = 16'h00E4; B = 16'h007; #100;
A = 16'h00E4; B = 16'h008; #100;
A = 16'h00E4; B = 16'h009; #100;
A = 16'h00E4; B = 16'h00A; #100;
A = 16'h00E4; B = 16'h00B; #100;
A = 16'h00E4; B = 16'h00C; #100;
A = 16'h00E4; B = 16'h00D; #100;
A = 16'h00E4; B = 16'h00E; #100;
A = 16'h00E4; B = 16'h00F; #100;
A = 16'h00E4; B = 16'h0010; #100;
A = 16'h00E4; B = 16'h0011; #100;
A = 16'h00E4; B = 16'h0012; #100;
A = 16'h00E4; B = 16'h0013; #100;
A = 16'h00E4; B = 16'h0014; #100;
A = 16'h00E4; B = 16'h0015; #100;
A = 16'h00E4; B = 16'h0016; #100;
A = 16'h00E4; B = 16'h0017; #100;
A = 16'h00E4; B = 16'h0018; #100;
A = 16'h00E4; B = 16'h0019; #100;
A = 16'h00E4; B = 16'h001A; #100;
A = 16'h00E4; B = 16'h001B; #100;
A = 16'h00E4; B = 16'h001C; #100;
A = 16'h00E4; B = 16'h001D; #100;
A = 16'h00E4; B = 16'h001E; #100;
A = 16'h00E4; B = 16'h001F; #100;
A = 16'h00E4; B = 16'h0020; #100;
A = 16'h00E4; B = 16'h0021; #100;
A = 16'h00E4; B = 16'h0022; #100;
A = 16'h00E4; B = 16'h0023; #100;
A = 16'h00E4; B = 16'h0024; #100;
A = 16'h00E4; B = 16'h0025; #100;
A = 16'h00E4; B = 16'h0026; #100;
A = 16'h00E4; B = 16'h0027; #100;
A = 16'h00E4; B = 16'h0028; #100;
A = 16'h00E4; B = 16'h0029; #100;
A = 16'h00E4; B = 16'h002A; #100;
A = 16'h00E4; B = 16'h002B; #100;
A = 16'h00E4; B = 16'h002C; #100;
A = 16'h00E4; B = 16'h002D; #100;
A = 16'h00E4; B = 16'h002E; #100;
A = 16'h00E4; B = 16'h002F; #100;
A = 16'h00E4; B = 16'h0030; #100;
A = 16'h00E4; B = 16'h0031; #100;
A = 16'h00E4; B = 16'h0032; #100;
A = 16'h00E4; B = 16'h0033; #100;
A = 16'h00E4; B = 16'h0034; #100;
A = 16'h00E4; B = 16'h0035; #100;
A = 16'h00E4; B = 16'h0036; #100;
A = 16'h00E4; B = 16'h0037; #100;
A = 16'h00E4; B = 16'h0038; #100;
A = 16'h00E4; B = 16'h0039; #100;
A = 16'h00E4; B = 16'h003A; #100;
A = 16'h00E4; B = 16'h003B; #100;
A = 16'h00E4; B = 16'h003C; #100;
A = 16'h00E4; B = 16'h003D; #100;
A = 16'h00E4; B = 16'h003E; #100;
A = 16'h00E4; B = 16'h003F; #100;
A = 16'h00E4; B = 16'h0040; #100;
A = 16'h00E4; B = 16'h0041; #100;
A = 16'h00E4; B = 16'h0042; #100;
A = 16'h00E4; B = 16'h0043; #100;
A = 16'h00E4; B = 16'h0044; #100;
A = 16'h00E4; B = 16'h0045; #100;
A = 16'h00E4; B = 16'h0046; #100;
A = 16'h00E4; B = 16'h0047; #100;
A = 16'h00E4; B = 16'h0048; #100;
A = 16'h00E4; B = 16'h0049; #100;
A = 16'h00E4; B = 16'h004A; #100;
A = 16'h00E4; B = 16'h004B; #100;
A = 16'h00E4; B = 16'h004C; #100;
A = 16'h00E4; B = 16'h004D; #100;
A = 16'h00E4; B = 16'h004E; #100;
A = 16'h00E4; B = 16'h004F; #100;
A = 16'h00E4; B = 16'h0050; #100;
A = 16'h00E4; B = 16'h0051; #100;
A = 16'h00E4; B = 16'h0052; #100;
A = 16'h00E4; B = 16'h0053; #100;
A = 16'h00E4; B = 16'h0054; #100;
A = 16'h00E4; B = 16'h0055; #100;
A = 16'h00E4; B = 16'h0056; #100;
A = 16'h00E4; B = 16'h0057; #100;
A = 16'h00E4; B = 16'h0058; #100;
A = 16'h00E4; B = 16'h0059; #100;
A = 16'h00E4; B = 16'h005A; #100;
A = 16'h00E4; B = 16'h005B; #100;
A = 16'h00E4; B = 16'h005C; #100;
A = 16'h00E4; B = 16'h005D; #100;
A = 16'h00E4; B = 16'h005E; #100;
A = 16'h00E4; B = 16'h005F; #100;
A = 16'h00E4; B = 16'h0060; #100;
A = 16'h00E4; B = 16'h0061; #100;
A = 16'h00E4; B = 16'h0062; #100;
A = 16'h00E4; B = 16'h0063; #100;
A = 16'h00E4; B = 16'h0064; #100;
A = 16'h00E4; B = 16'h0065; #100;
A = 16'h00E4; B = 16'h0066; #100;
A = 16'h00E4; B = 16'h0067; #100;
A = 16'h00E4; B = 16'h0068; #100;
A = 16'h00E4; B = 16'h0069; #100;
A = 16'h00E4; B = 16'h006A; #100;
A = 16'h00E4; B = 16'h006B; #100;
A = 16'h00E4; B = 16'h006C; #100;
A = 16'h00E4; B = 16'h006D; #100;
A = 16'h00E4; B = 16'h006E; #100;
A = 16'h00E4; B = 16'h006F; #100;
A = 16'h00E4; B = 16'h0070; #100;
A = 16'h00E4; B = 16'h0071; #100;
A = 16'h00E4; B = 16'h0072; #100;
A = 16'h00E4; B = 16'h0073; #100;
A = 16'h00E4; B = 16'h0074; #100;
A = 16'h00E4; B = 16'h0075; #100;
A = 16'h00E4; B = 16'h0076; #100;
A = 16'h00E4; B = 16'h0077; #100;
A = 16'h00E4; B = 16'h0078; #100;
A = 16'h00E4; B = 16'h0079; #100;
A = 16'h00E4; B = 16'h007A; #100;
A = 16'h00E4; B = 16'h007B; #100;
A = 16'h00E4; B = 16'h007C; #100;
A = 16'h00E4; B = 16'h007D; #100;
A = 16'h00E4; B = 16'h007E; #100;
A = 16'h00E4; B = 16'h007F; #100;
A = 16'h00E4; B = 16'h0080; #100;
A = 16'h00E4; B = 16'h0081; #100;
A = 16'h00E4; B = 16'h0082; #100;
A = 16'h00E4; B = 16'h0083; #100;
A = 16'h00E4; B = 16'h0084; #100;
A = 16'h00E4; B = 16'h0085; #100;
A = 16'h00E4; B = 16'h0086; #100;
A = 16'h00E4; B = 16'h0087; #100;
A = 16'h00E4; B = 16'h0088; #100;
A = 16'h00E4; B = 16'h0089; #100;
A = 16'h00E4; B = 16'h008A; #100;
A = 16'h00E4; B = 16'h008B; #100;
A = 16'h00E4; B = 16'h008C; #100;
A = 16'h00E4; B = 16'h008D; #100;
A = 16'h00E4; B = 16'h008E; #100;
A = 16'h00E4; B = 16'h008F; #100;
A = 16'h00E4; B = 16'h0090; #100;
A = 16'h00E4; B = 16'h0091; #100;
A = 16'h00E4; B = 16'h0092; #100;
A = 16'h00E4; B = 16'h0093; #100;
A = 16'h00E4; B = 16'h0094; #100;
A = 16'h00E4; B = 16'h0095; #100;
A = 16'h00E4; B = 16'h0096; #100;
A = 16'h00E4; B = 16'h0097; #100;
A = 16'h00E4; B = 16'h0098; #100;
A = 16'h00E4; B = 16'h0099; #100;
A = 16'h00E4; B = 16'h009A; #100;
A = 16'h00E4; B = 16'h009B; #100;
A = 16'h00E4; B = 16'h009C; #100;
A = 16'h00E4; B = 16'h009D; #100;
A = 16'h00E4; B = 16'h009E; #100;
A = 16'h00E4; B = 16'h009F; #100;
A = 16'h00E4; B = 16'h00A0; #100;
A = 16'h00E4; B = 16'h00A1; #100;
A = 16'h00E4; B = 16'h00A2; #100;
A = 16'h00E4; B = 16'h00A3; #100;
A = 16'h00E4; B = 16'h00A4; #100;
A = 16'h00E4; B = 16'h00A5; #100;
A = 16'h00E4; B = 16'h00A6; #100;
A = 16'h00E4; B = 16'h00A7; #100;
A = 16'h00E4; B = 16'h00A8; #100;
A = 16'h00E4; B = 16'h00A9; #100;
A = 16'h00E4; B = 16'h00AA; #100;
A = 16'h00E4; B = 16'h00AB; #100;
A = 16'h00E4; B = 16'h00AC; #100;
A = 16'h00E4; B = 16'h00AD; #100;
A = 16'h00E4; B = 16'h00AE; #100;
A = 16'h00E4; B = 16'h00AF; #100;
A = 16'h00E4; B = 16'h00B0; #100;
A = 16'h00E4; B = 16'h00B1; #100;
A = 16'h00E4; B = 16'h00B2; #100;
A = 16'h00E4; B = 16'h00B3; #100;
A = 16'h00E4; B = 16'h00B4; #100;
A = 16'h00E4; B = 16'h00B5; #100;
A = 16'h00E4; B = 16'h00B6; #100;
A = 16'h00E4; B = 16'h00B7; #100;
A = 16'h00E4; B = 16'h00B8; #100;
A = 16'h00E4; B = 16'h00B9; #100;
A = 16'h00E4; B = 16'h00BA; #100;
A = 16'h00E4; B = 16'h00BB; #100;
A = 16'h00E4; B = 16'h00BC; #100;
A = 16'h00E4; B = 16'h00BD; #100;
A = 16'h00E4; B = 16'h00BE; #100;
A = 16'h00E4; B = 16'h00BF; #100;
A = 16'h00E4; B = 16'h00C0; #100;
A = 16'h00E4; B = 16'h00C1; #100;
A = 16'h00E4; B = 16'h00C2; #100;
A = 16'h00E4; B = 16'h00C3; #100;
A = 16'h00E4; B = 16'h00C4; #100;
A = 16'h00E4; B = 16'h00C5; #100;
A = 16'h00E4; B = 16'h00C6; #100;
A = 16'h00E4; B = 16'h00C7; #100;
A = 16'h00E4; B = 16'h00C8; #100;
A = 16'h00E4; B = 16'h00C9; #100;
A = 16'h00E4; B = 16'h00CA; #100;
A = 16'h00E4; B = 16'h00CB; #100;
A = 16'h00E4; B = 16'h00CC; #100;
A = 16'h00E4; B = 16'h00CD; #100;
A = 16'h00E4; B = 16'h00CE; #100;
A = 16'h00E4; B = 16'h00CF; #100;
A = 16'h00E4; B = 16'h00D0; #100;
A = 16'h00E4; B = 16'h00D1; #100;
A = 16'h00E4; B = 16'h00D2; #100;
A = 16'h00E4; B = 16'h00D3; #100;
A = 16'h00E4; B = 16'h00D4; #100;
A = 16'h00E4; B = 16'h00D5; #100;
A = 16'h00E4; B = 16'h00D6; #100;
A = 16'h00E4; B = 16'h00D7; #100;
A = 16'h00E4; B = 16'h00D8; #100;
A = 16'h00E4; B = 16'h00D9; #100;
A = 16'h00E4; B = 16'h00DA; #100;
A = 16'h00E4; B = 16'h00DB; #100;
A = 16'h00E4; B = 16'h00DC; #100;
A = 16'h00E4; B = 16'h00DD; #100;
A = 16'h00E4; B = 16'h00DE; #100;
A = 16'h00E4; B = 16'h00DF; #100;
A = 16'h00E4; B = 16'h00E0; #100;
A = 16'h00E4; B = 16'h00E1; #100;
A = 16'h00E4; B = 16'h00E2; #100;
A = 16'h00E4; B = 16'h00E3; #100;
A = 16'h00E4; B = 16'h00E4; #100;
A = 16'h00E4; B = 16'h00E5; #100;
A = 16'h00E4; B = 16'h00E6; #100;
A = 16'h00E4; B = 16'h00E7; #100;
A = 16'h00E4; B = 16'h00E8; #100;
A = 16'h00E4; B = 16'h00E9; #100;
A = 16'h00E4; B = 16'h00EA; #100;
A = 16'h00E4; B = 16'h00EB; #100;
A = 16'h00E4; B = 16'h00EC; #100;
A = 16'h00E4; B = 16'h00ED; #100;
A = 16'h00E4; B = 16'h00EE; #100;
A = 16'h00E4; B = 16'h00EF; #100;
A = 16'h00E4; B = 16'h00F0; #100;
A = 16'h00E4; B = 16'h00F1; #100;
A = 16'h00E4; B = 16'h00F2; #100;
A = 16'h00E4; B = 16'h00F3; #100;
A = 16'h00E4; B = 16'h00F4; #100;
A = 16'h00E4; B = 16'h00F5; #100;
A = 16'h00E4; B = 16'h00F6; #100;
A = 16'h00E4; B = 16'h00F7; #100;
A = 16'h00E4; B = 16'h00F8; #100;
A = 16'h00E4; B = 16'h00F9; #100;
A = 16'h00E4; B = 16'h00FA; #100;
A = 16'h00E4; B = 16'h00FB; #100;
A = 16'h00E4; B = 16'h00FC; #100;
A = 16'h00E4; B = 16'h00FD; #100;
A = 16'h00E4; B = 16'h00FE; #100;
A = 16'h00E4; B = 16'h00FF; #100;
A = 16'h00E5; B = 16'h000; #100;
A = 16'h00E5; B = 16'h001; #100;
A = 16'h00E5; B = 16'h002; #100;
A = 16'h00E5; B = 16'h003; #100;
A = 16'h00E5; B = 16'h004; #100;
A = 16'h00E5; B = 16'h005; #100;
A = 16'h00E5; B = 16'h006; #100;
A = 16'h00E5; B = 16'h007; #100;
A = 16'h00E5; B = 16'h008; #100;
A = 16'h00E5; B = 16'h009; #100;
A = 16'h00E5; B = 16'h00A; #100;
A = 16'h00E5; B = 16'h00B; #100;
A = 16'h00E5; B = 16'h00C; #100;
A = 16'h00E5; B = 16'h00D; #100;
A = 16'h00E5; B = 16'h00E; #100;
A = 16'h00E5; B = 16'h00F; #100;
A = 16'h00E5; B = 16'h0010; #100;
A = 16'h00E5; B = 16'h0011; #100;
A = 16'h00E5; B = 16'h0012; #100;
A = 16'h00E5; B = 16'h0013; #100;
A = 16'h00E5; B = 16'h0014; #100;
A = 16'h00E5; B = 16'h0015; #100;
A = 16'h00E5; B = 16'h0016; #100;
A = 16'h00E5; B = 16'h0017; #100;
A = 16'h00E5; B = 16'h0018; #100;
A = 16'h00E5; B = 16'h0019; #100;
A = 16'h00E5; B = 16'h001A; #100;
A = 16'h00E5; B = 16'h001B; #100;
A = 16'h00E5; B = 16'h001C; #100;
A = 16'h00E5; B = 16'h001D; #100;
A = 16'h00E5; B = 16'h001E; #100;
A = 16'h00E5; B = 16'h001F; #100;
A = 16'h00E5; B = 16'h0020; #100;
A = 16'h00E5; B = 16'h0021; #100;
A = 16'h00E5; B = 16'h0022; #100;
A = 16'h00E5; B = 16'h0023; #100;
A = 16'h00E5; B = 16'h0024; #100;
A = 16'h00E5; B = 16'h0025; #100;
A = 16'h00E5; B = 16'h0026; #100;
A = 16'h00E5; B = 16'h0027; #100;
A = 16'h00E5; B = 16'h0028; #100;
A = 16'h00E5; B = 16'h0029; #100;
A = 16'h00E5; B = 16'h002A; #100;
A = 16'h00E5; B = 16'h002B; #100;
A = 16'h00E5; B = 16'h002C; #100;
A = 16'h00E5; B = 16'h002D; #100;
A = 16'h00E5; B = 16'h002E; #100;
A = 16'h00E5; B = 16'h002F; #100;
A = 16'h00E5; B = 16'h0030; #100;
A = 16'h00E5; B = 16'h0031; #100;
A = 16'h00E5; B = 16'h0032; #100;
A = 16'h00E5; B = 16'h0033; #100;
A = 16'h00E5; B = 16'h0034; #100;
A = 16'h00E5; B = 16'h0035; #100;
A = 16'h00E5; B = 16'h0036; #100;
A = 16'h00E5; B = 16'h0037; #100;
A = 16'h00E5; B = 16'h0038; #100;
A = 16'h00E5; B = 16'h0039; #100;
A = 16'h00E5; B = 16'h003A; #100;
A = 16'h00E5; B = 16'h003B; #100;
A = 16'h00E5; B = 16'h003C; #100;
A = 16'h00E5; B = 16'h003D; #100;
A = 16'h00E5; B = 16'h003E; #100;
A = 16'h00E5; B = 16'h003F; #100;
A = 16'h00E5; B = 16'h0040; #100;
A = 16'h00E5; B = 16'h0041; #100;
A = 16'h00E5; B = 16'h0042; #100;
A = 16'h00E5; B = 16'h0043; #100;
A = 16'h00E5; B = 16'h0044; #100;
A = 16'h00E5; B = 16'h0045; #100;
A = 16'h00E5; B = 16'h0046; #100;
A = 16'h00E5; B = 16'h0047; #100;
A = 16'h00E5; B = 16'h0048; #100;
A = 16'h00E5; B = 16'h0049; #100;
A = 16'h00E5; B = 16'h004A; #100;
A = 16'h00E5; B = 16'h004B; #100;
A = 16'h00E5; B = 16'h004C; #100;
A = 16'h00E5; B = 16'h004D; #100;
A = 16'h00E5; B = 16'h004E; #100;
A = 16'h00E5; B = 16'h004F; #100;
A = 16'h00E5; B = 16'h0050; #100;
A = 16'h00E5; B = 16'h0051; #100;
A = 16'h00E5; B = 16'h0052; #100;
A = 16'h00E5; B = 16'h0053; #100;
A = 16'h00E5; B = 16'h0054; #100;
A = 16'h00E5; B = 16'h0055; #100;
A = 16'h00E5; B = 16'h0056; #100;
A = 16'h00E5; B = 16'h0057; #100;
A = 16'h00E5; B = 16'h0058; #100;
A = 16'h00E5; B = 16'h0059; #100;
A = 16'h00E5; B = 16'h005A; #100;
A = 16'h00E5; B = 16'h005B; #100;
A = 16'h00E5; B = 16'h005C; #100;
A = 16'h00E5; B = 16'h005D; #100;
A = 16'h00E5; B = 16'h005E; #100;
A = 16'h00E5; B = 16'h005F; #100;
A = 16'h00E5; B = 16'h0060; #100;
A = 16'h00E5; B = 16'h0061; #100;
A = 16'h00E5; B = 16'h0062; #100;
A = 16'h00E5; B = 16'h0063; #100;
A = 16'h00E5; B = 16'h0064; #100;
A = 16'h00E5; B = 16'h0065; #100;
A = 16'h00E5; B = 16'h0066; #100;
A = 16'h00E5; B = 16'h0067; #100;
A = 16'h00E5; B = 16'h0068; #100;
A = 16'h00E5; B = 16'h0069; #100;
A = 16'h00E5; B = 16'h006A; #100;
A = 16'h00E5; B = 16'h006B; #100;
A = 16'h00E5; B = 16'h006C; #100;
A = 16'h00E5; B = 16'h006D; #100;
A = 16'h00E5; B = 16'h006E; #100;
A = 16'h00E5; B = 16'h006F; #100;
A = 16'h00E5; B = 16'h0070; #100;
A = 16'h00E5; B = 16'h0071; #100;
A = 16'h00E5; B = 16'h0072; #100;
A = 16'h00E5; B = 16'h0073; #100;
A = 16'h00E5; B = 16'h0074; #100;
A = 16'h00E5; B = 16'h0075; #100;
A = 16'h00E5; B = 16'h0076; #100;
A = 16'h00E5; B = 16'h0077; #100;
A = 16'h00E5; B = 16'h0078; #100;
A = 16'h00E5; B = 16'h0079; #100;
A = 16'h00E5; B = 16'h007A; #100;
A = 16'h00E5; B = 16'h007B; #100;
A = 16'h00E5; B = 16'h007C; #100;
A = 16'h00E5; B = 16'h007D; #100;
A = 16'h00E5; B = 16'h007E; #100;
A = 16'h00E5; B = 16'h007F; #100;
A = 16'h00E5; B = 16'h0080; #100;
A = 16'h00E5; B = 16'h0081; #100;
A = 16'h00E5; B = 16'h0082; #100;
A = 16'h00E5; B = 16'h0083; #100;
A = 16'h00E5; B = 16'h0084; #100;
A = 16'h00E5; B = 16'h0085; #100;
A = 16'h00E5; B = 16'h0086; #100;
A = 16'h00E5; B = 16'h0087; #100;
A = 16'h00E5; B = 16'h0088; #100;
A = 16'h00E5; B = 16'h0089; #100;
A = 16'h00E5; B = 16'h008A; #100;
A = 16'h00E5; B = 16'h008B; #100;
A = 16'h00E5; B = 16'h008C; #100;
A = 16'h00E5; B = 16'h008D; #100;
A = 16'h00E5; B = 16'h008E; #100;
A = 16'h00E5; B = 16'h008F; #100;
A = 16'h00E5; B = 16'h0090; #100;
A = 16'h00E5; B = 16'h0091; #100;
A = 16'h00E5; B = 16'h0092; #100;
A = 16'h00E5; B = 16'h0093; #100;
A = 16'h00E5; B = 16'h0094; #100;
A = 16'h00E5; B = 16'h0095; #100;
A = 16'h00E5; B = 16'h0096; #100;
A = 16'h00E5; B = 16'h0097; #100;
A = 16'h00E5; B = 16'h0098; #100;
A = 16'h00E5; B = 16'h0099; #100;
A = 16'h00E5; B = 16'h009A; #100;
A = 16'h00E5; B = 16'h009B; #100;
A = 16'h00E5; B = 16'h009C; #100;
A = 16'h00E5; B = 16'h009D; #100;
A = 16'h00E5; B = 16'h009E; #100;
A = 16'h00E5; B = 16'h009F; #100;
A = 16'h00E5; B = 16'h00A0; #100;
A = 16'h00E5; B = 16'h00A1; #100;
A = 16'h00E5; B = 16'h00A2; #100;
A = 16'h00E5; B = 16'h00A3; #100;
A = 16'h00E5; B = 16'h00A4; #100;
A = 16'h00E5; B = 16'h00A5; #100;
A = 16'h00E5; B = 16'h00A6; #100;
A = 16'h00E5; B = 16'h00A7; #100;
A = 16'h00E5; B = 16'h00A8; #100;
A = 16'h00E5; B = 16'h00A9; #100;
A = 16'h00E5; B = 16'h00AA; #100;
A = 16'h00E5; B = 16'h00AB; #100;
A = 16'h00E5; B = 16'h00AC; #100;
A = 16'h00E5; B = 16'h00AD; #100;
A = 16'h00E5; B = 16'h00AE; #100;
A = 16'h00E5; B = 16'h00AF; #100;
A = 16'h00E5; B = 16'h00B0; #100;
A = 16'h00E5; B = 16'h00B1; #100;
A = 16'h00E5; B = 16'h00B2; #100;
A = 16'h00E5; B = 16'h00B3; #100;
A = 16'h00E5; B = 16'h00B4; #100;
A = 16'h00E5; B = 16'h00B5; #100;
A = 16'h00E5; B = 16'h00B6; #100;
A = 16'h00E5; B = 16'h00B7; #100;
A = 16'h00E5; B = 16'h00B8; #100;
A = 16'h00E5; B = 16'h00B9; #100;
A = 16'h00E5; B = 16'h00BA; #100;
A = 16'h00E5; B = 16'h00BB; #100;
A = 16'h00E5; B = 16'h00BC; #100;
A = 16'h00E5; B = 16'h00BD; #100;
A = 16'h00E5; B = 16'h00BE; #100;
A = 16'h00E5; B = 16'h00BF; #100;
A = 16'h00E5; B = 16'h00C0; #100;
A = 16'h00E5; B = 16'h00C1; #100;
A = 16'h00E5; B = 16'h00C2; #100;
A = 16'h00E5; B = 16'h00C3; #100;
A = 16'h00E5; B = 16'h00C4; #100;
A = 16'h00E5; B = 16'h00C5; #100;
A = 16'h00E5; B = 16'h00C6; #100;
A = 16'h00E5; B = 16'h00C7; #100;
A = 16'h00E5; B = 16'h00C8; #100;
A = 16'h00E5; B = 16'h00C9; #100;
A = 16'h00E5; B = 16'h00CA; #100;
A = 16'h00E5; B = 16'h00CB; #100;
A = 16'h00E5; B = 16'h00CC; #100;
A = 16'h00E5; B = 16'h00CD; #100;
A = 16'h00E5; B = 16'h00CE; #100;
A = 16'h00E5; B = 16'h00CF; #100;
A = 16'h00E5; B = 16'h00D0; #100;
A = 16'h00E5; B = 16'h00D1; #100;
A = 16'h00E5; B = 16'h00D2; #100;
A = 16'h00E5; B = 16'h00D3; #100;
A = 16'h00E5; B = 16'h00D4; #100;
A = 16'h00E5; B = 16'h00D5; #100;
A = 16'h00E5; B = 16'h00D6; #100;
A = 16'h00E5; B = 16'h00D7; #100;
A = 16'h00E5; B = 16'h00D8; #100;
A = 16'h00E5; B = 16'h00D9; #100;
A = 16'h00E5; B = 16'h00DA; #100;
A = 16'h00E5; B = 16'h00DB; #100;
A = 16'h00E5; B = 16'h00DC; #100;
A = 16'h00E5; B = 16'h00DD; #100;
A = 16'h00E5; B = 16'h00DE; #100;
A = 16'h00E5; B = 16'h00DF; #100;
A = 16'h00E5; B = 16'h00E0; #100;
A = 16'h00E5; B = 16'h00E1; #100;
A = 16'h00E5; B = 16'h00E2; #100;
A = 16'h00E5; B = 16'h00E3; #100;
A = 16'h00E5; B = 16'h00E4; #100;
A = 16'h00E5; B = 16'h00E5; #100;
A = 16'h00E5; B = 16'h00E6; #100;
A = 16'h00E5; B = 16'h00E7; #100;
A = 16'h00E5; B = 16'h00E8; #100;
A = 16'h00E5; B = 16'h00E9; #100;
A = 16'h00E5; B = 16'h00EA; #100;
A = 16'h00E5; B = 16'h00EB; #100;
A = 16'h00E5; B = 16'h00EC; #100;
A = 16'h00E5; B = 16'h00ED; #100;
A = 16'h00E5; B = 16'h00EE; #100;
A = 16'h00E5; B = 16'h00EF; #100;
A = 16'h00E5; B = 16'h00F0; #100;
A = 16'h00E5; B = 16'h00F1; #100;
A = 16'h00E5; B = 16'h00F2; #100;
A = 16'h00E5; B = 16'h00F3; #100;
A = 16'h00E5; B = 16'h00F4; #100;
A = 16'h00E5; B = 16'h00F5; #100;
A = 16'h00E5; B = 16'h00F6; #100;
A = 16'h00E5; B = 16'h00F7; #100;
A = 16'h00E5; B = 16'h00F8; #100;
A = 16'h00E5; B = 16'h00F9; #100;
A = 16'h00E5; B = 16'h00FA; #100;
A = 16'h00E5; B = 16'h00FB; #100;
A = 16'h00E5; B = 16'h00FC; #100;
A = 16'h00E5; B = 16'h00FD; #100;
A = 16'h00E5; B = 16'h00FE; #100;
A = 16'h00E5; B = 16'h00FF; #100;
A = 16'h00E6; B = 16'h000; #100;
A = 16'h00E6; B = 16'h001; #100;
A = 16'h00E6; B = 16'h002; #100;
A = 16'h00E6; B = 16'h003; #100;
A = 16'h00E6; B = 16'h004; #100;
A = 16'h00E6; B = 16'h005; #100;
A = 16'h00E6; B = 16'h006; #100;
A = 16'h00E6; B = 16'h007; #100;
A = 16'h00E6; B = 16'h008; #100;
A = 16'h00E6; B = 16'h009; #100;
A = 16'h00E6; B = 16'h00A; #100;
A = 16'h00E6; B = 16'h00B; #100;
A = 16'h00E6; B = 16'h00C; #100;
A = 16'h00E6; B = 16'h00D; #100;
A = 16'h00E6; B = 16'h00E; #100;
A = 16'h00E6; B = 16'h00F; #100;
A = 16'h00E6; B = 16'h0010; #100;
A = 16'h00E6; B = 16'h0011; #100;
A = 16'h00E6; B = 16'h0012; #100;
A = 16'h00E6; B = 16'h0013; #100;
A = 16'h00E6; B = 16'h0014; #100;
A = 16'h00E6; B = 16'h0015; #100;
A = 16'h00E6; B = 16'h0016; #100;
A = 16'h00E6; B = 16'h0017; #100;
A = 16'h00E6; B = 16'h0018; #100;
A = 16'h00E6; B = 16'h0019; #100;
A = 16'h00E6; B = 16'h001A; #100;
A = 16'h00E6; B = 16'h001B; #100;
A = 16'h00E6; B = 16'h001C; #100;
A = 16'h00E6; B = 16'h001D; #100;
A = 16'h00E6; B = 16'h001E; #100;
A = 16'h00E6; B = 16'h001F; #100;
A = 16'h00E6; B = 16'h0020; #100;
A = 16'h00E6; B = 16'h0021; #100;
A = 16'h00E6; B = 16'h0022; #100;
A = 16'h00E6; B = 16'h0023; #100;
A = 16'h00E6; B = 16'h0024; #100;
A = 16'h00E6; B = 16'h0025; #100;
A = 16'h00E6; B = 16'h0026; #100;
A = 16'h00E6; B = 16'h0027; #100;
A = 16'h00E6; B = 16'h0028; #100;
A = 16'h00E6; B = 16'h0029; #100;
A = 16'h00E6; B = 16'h002A; #100;
A = 16'h00E6; B = 16'h002B; #100;
A = 16'h00E6; B = 16'h002C; #100;
A = 16'h00E6; B = 16'h002D; #100;
A = 16'h00E6; B = 16'h002E; #100;
A = 16'h00E6; B = 16'h002F; #100;
A = 16'h00E6; B = 16'h0030; #100;
A = 16'h00E6; B = 16'h0031; #100;
A = 16'h00E6; B = 16'h0032; #100;
A = 16'h00E6; B = 16'h0033; #100;
A = 16'h00E6; B = 16'h0034; #100;
A = 16'h00E6; B = 16'h0035; #100;
A = 16'h00E6; B = 16'h0036; #100;
A = 16'h00E6; B = 16'h0037; #100;
A = 16'h00E6; B = 16'h0038; #100;
A = 16'h00E6; B = 16'h0039; #100;
A = 16'h00E6; B = 16'h003A; #100;
A = 16'h00E6; B = 16'h003B; #100;
A = 16'h00E6; B = 16'h003C; #100;
A = 16'h00E6; B = 16'h003D; #100;
A = 16'h00E6; B = 16'h003E; #100;
A = 16'h00E6; B = 16'h003F; #100;
A = 16'h00E6; B = 16'h0040; #100;
A = 16'h00E6; B = 16'h0041; #100;
A = 16'h00E6; B = 16'h0042; #100;
A = 16'h00E6; B = 16'h0043; #100;
A = 16'h00E6; B = 16'h0044; #100;
A = 16'h00E6; B = 16'h0045; #100;
A = 16'h00E6; B = 16'h0046; #100;
A = 16'h00E6; B = 16'h0047; #100;
A = 16'h00E6; B = 16'h0048; #100;
A = 16'h00E6; B = 16'h0049; #100;
A = 16'h00E6; B = 16'h004A; #100;
A = 16'h00E6; B = 16'h004B; #100;
A = 16'h00E6; B = 16'h004C; #100;
A = 16'h00E6; B = 16'h004D; #100;
A = 16'h00E6; B = 16'h004E; #100;
A = 16'h00E6; B = 16'h004F; #100;
A = 16'h00E6; B = 16'h0050; #100;
A = 16'h00E6; B = 16'h0051; #100;
A = 16'h00E6; B = 16'h0052; #100;
A = 16'h00E6; B = 16'h0053; #100;
A = 16'h00E6; B = 16'h0054; #100;
A = 16'h00E6; B = 16'h0055; #100;
A = 16'h00E6; B = 16'h0056; #100;
A = 16'h00E6; B = 16'h0057; #100;
A = 16'h00E6; B = 16'h0058; #100;
A = 16'h00E6; B = 16'h0059; #100;
A = 16'h00E6; B = 16'h005A; #100;
A = 16'h00E6; B = 16'h005B; #100;
A = 16'h00E6; B = 16'h005C; #100;
A = 16'h00E6; B = 16'h005D; #100;
A = 16'h00E6; B = 16'h005E; #100;
A = 16'h00E6; B = 16'h005F; #100;
A = 16'h00E6; B = 16'h0060; #100;
A = 16'h00E6; B = 16'h0061; #100;
A = 16'h00E6; B = 16'h0062; #100;
A = 16'h00E6; B = 16'h0063; #100;
A = 16'h00E6; B = 16'h0064; #100;
A = 16'h00E6; B = 16'h0065; #100;
A = 16'h00E6; B = 16'h0066; #100;
A = 16'h00E6; B = 16'h0067; #100;
A = 16'h00E6; B = 16'h0068; #100;
A = 16'h00E6; B = 16'h0069; #100;
A = 16'h00E6; B = 16'h006A; #100;
A = 16'h00E6; B = 16'h006B; #100;
A = 16'h00E6; B = 16'h006C; #100;
A = 16'h00E6; B = 16'h006D; #100;
A = 16'h00E6; B = 16'h006E; #100;
A = 16'h00E6; B = 16'h006F; #100;
A = 16'h00E6; B = 16'h0070; #100;
A = 16'h00E6; B = 16'h0071; #100;
A = 16'h00E6; B = 16'h0072; #100;
A = 16'h00E6; B = 16'h0073; #100;
A = 16'h00E6; B = 16'h0074; #100;
A = 16'h00E6; B = 16'h0075; #100;
A = 16'h00E6; B = 16'h0076; #100;
A = 16'h00E6; B = 16'h0077; #100;
A = 16'h00E6; B = 16'h0078; #100;
A = 16'h00E6; B = 16'h0079; #100;
A = 16'h00E6; B = 16'h007A; #100;
A = 16'h00E6; B = 16'h007B; #100;
A = 16'h00E6; B = 16'h007C; #100;
A = 16'h00E6; B = 16'h007D; #100;
A = 16'h00E6; B = 16'h007E; #100;
A = 16'h00E6; B = 16'h007F; #100;
A = 16'h00E6; B = 16'h0080; #100;
A = 16'h00E6; B = 16'h0081; #100;
A = 16'h00E6; B = 16'h0082; #100;
A = 16'h00E6; B = 16'h0083; #100;
A = 16'h00E6; B = 16'h0084; #100;
A = 16'h00E6; B = 16'h0085; #100;
A = 16'h00E6; B = 16'h0086; #100;
A = 16'h00E6; B = 16'h0087; #100;
A = 16'h00E6; B = 16'h0088; #100;
A = 16'h00E6; B = 16'h0089; #100;
A = 16'h00E6; B = 16'h008A; #100;
A = 16'h00E6; B = 16'h008B; #100;
A = 16'h00E6; B = 16'h008C; #100;
A = 16'h00E6; B = 16'h008D; #100;
A = 16'h00E6; B = 16'h008E; #100;
A = 16'h00E6; B = 16'h008F; #100;
A = 16'h00E6; B = 16'h0090; #100;
A = 16'h00E6; B = 16'h0091; #100;
A = 16'h00E6; B = 16'h0092; #100;
A = 16'h00E6; B = 16'h0093; #100;
A = 16'h00E6; B = 16'h0094; #100;
A = 16'h00E6; B = 16'h0095; #100;
A = 16'h00E6; B = 16'h0096; #100;
A = 16'h00E6; B = 16'h0097; #100;
A = 16'h00E6; B = 16'h0098; #100;
A = 16'h00E6; B = 16'h0099; #100;
A = 16'h00E6; B = 16'h009A; #100;
A = 16'h00E6; B = 16'h009B; #100;
A = 16'h00E6; B = 16'h009C; #100;
A = 16'h00E6; B = 16'h009D; #100;
A = 16'h00E6; B = 16'h009E; #100;
A = 16'h00E6; B = 16'h009F; #100;
A = 16'h00E6; B = 16'h00A0; #100;
A = 16'h00E6; B = 16'h00A1; #100;
A = 16'h00E6; B = 16'h00A2; #100;
A = 16'h00E6; B = 16'h00A3; #100;
A = 16'h00E6; B = 16'h00A4; #100;
A = 16'h00E6; B = 16'h00A5; #100;
A = 16'h00E6; B = 16'h00A6; #100;
A = 16'h00E6; B = 16'h00A7; #100;
A = 16'h00E6; B = 16'h00A8; #100;
A = 16'h00E6; B = 16'h00A9; #100;
A = 16'h00E6; B = 16'h00AA; #100;
A = 16'h00E6; B = 16'h00AB; #100;
A = 16'h00E6; B = 16'h00AC; #100;
A = 16'h00E6; B = 16'h00AD; #100;
A = 16'h00E6; B = 16'h00AE; #100;
A = 16'h00E6; B = 16'h00AF; #100;
A = 16'h00E6; B = 16'h00B0; #100;
A = 16'h00E6; B = 16'h00B1; #100;
A = 16'h00E6; B = 16'h00B2; #100;
A = 16'h00E6; B = 16'h00B3; #100;
A = 16'h00E6; B = 16'h00B4; #100;
A = 16'h00E6; B = 16'h00B5; #100;
A = 16'h00E6; B = 16'h00B6; #100;
A = 16'h00E6; B = 16'h00B7; #100;
A = 16'h00E6; B = 16'h00B8; #100;
A = 16'h00E6; B = 16'h00B9; #100;
A = 16'h00E6; B = 16'h00BA; #100;
A = 16'h00E6; B = 16'h00BB; #100;
A = 16'h00E6; B = 16'h00BC; #100;
A = 16'h00E6; B = 16'h00BD; #100;
A = 16'h00E6; B = 16'h00BE; #100;
A = 16'h00E6; B = 16'h00BF; #100;
A = 16'h00E6; B = 16'h00C0; #100;
A = 16'h00E6; B = 16'h00C1; #100;
A = 16'h00E6; B = 16'h00C2; #100;
A = 16'h00E6; B = 16'h00C3; #100;
A = 16'h00E6; B = 16'h00C4; #100;
A = 16'h00E6; B = 16'h00C5; #100;
A = 16'h00E6; B = 16'h00C6; #100;
A = 16'h00E6; B = 16'h00C7; #100;
A = 16'h00E6; B = 16'h00C8; #100;
A = 16'h00E6; B = 16'h00C9; #100;
A = 16'h00E6; B = 16'h00CA; #100;
A = 16'h00E6; B = 16'h00CB; #100;
A = 16'h00E6; B = 16'h00CC; #100;
A = 16'h00E6; B = 16'h00CD; #100;
A = 16'h00E6; B = 16'h00CE; #100;
A = 16'h00E6; B = 16'h00CF; #100;
A = 16'h00E6; B = 16'h00D0; #100;
A = 16'h00E6; B = 16'h00D1; #100;
A = 16'h00E6; B = 16'h00D2; #100;
A = 16'h00E6; B = 16'h00D3; #100;
A = 16'h00E6; B = 16'h00D4; #100;
A = 16'h00E6; B = 16'h00D5; #100;
A = 16'h00E6; B = 16'h00D6; #100;
A = 16'h00E6; B = 16'h00D7; #100;
A = 16'h00E6; B = 16'h00D8; #100;
A = 16'h00E6; B = 16'h00D9; #100;
A = 16'h00E6; B = 16'h00DA; #100;
A = 16'h00E6; B = 16'h00DB; #100;
A = 16'h00E6; B = 16'h00DC; #100;
A = 16'h00E6; B = 16'h00DD; #100;
A = 16'h00E6; B = 16'h00DE; #100;
A = 16'h00E6; B = 16'h00DF; #100;
A = 16'h00E6; B = 16'h00E0; #100;
A = 16'h00E6; B = 16'h00E1; #100;
A = 16'h00E6; B = 16'h00E2; #100;
A = 16'h00E6; B = 16'h00E3; #100;
A = 16'h00E6; B = 16'h00E4; #100;
A = 16'h00E6; B = 16'h00E5; #100;
A = 16'h00E6; B = 16'h00E6; #100;
A = 16'h00E6; B = 16'h00E7; #100;
A = 16'h00E6; B = 16'h00E8; #100;
A = 16'h00E6; B = 16'h00E9; #100;
A = 16'h00E6; B = 16'h00EA; #100;
A = 16'h00E6; B = 16'h00EB; #100;
A = 16'h00E6; B = 16'h00EC; #100;
A = 16'h00E6; B = 16'h00ED; #100;
A = 16'h00E6; B = 16'h00EE; #100;
A = 16'h00E6; B = 16'h00EF; #100;
A = 16'h00E6; B = 16'h00F0; #100;
A = 16'h00E6; B = 16'h00F1; #100;
A = 16'h00E6; B = 16'h00F2; #100;
A = 16'h00E6; B = 16'h00F3; #100;
A = 16'h00E6; B = 16'h00F4; #100;
A = 16'h00E6; B = 16'h00F5; #100;
A = 16'h00E6; B = 16'h00F6; #100;
A = 16'h00E6; B = 16'h00F7; #100;
A = 16'h00E6; B = 16'h00F8; #100;
A = 16'h00E6; B = 16'h00F9; #100;
A = 16'h00E6; B = 16'h00FA; #100;
A = 16'h00E6; B = 16'h00FB; #100;
A = 16'h00E6; B = 16'h00FC; #100;
A = 16'h00E6; B = 16'h00FD; #100;
A = 16'h00E6; B = 16'h00FE; #100;
A = 16'h00E6; B = 16'h00FF; #100;
A = 16'h00E7; B = 16'h000; #100;
A = 16'h00E7; B = 16'h001; #100;
A = 16'h00E7; B = 16'h002; #100;
A = 16'h00E7; B = 16'h003; #100;
A = 16'h00E7; B = 16'h004; #100;
A = 16'h00E7; B = 16'h005; #100;
A = 16'h00E7; B = 16'h006; #100;
A = 16'h00E7; B = 16'h007; #100;
A = 16'h00E7; B = 16'h008; #100;
A = 16'h00E7; B = 16'h009; #100;
A = 16'h00E7; B = 16'h00A; #100;
A = 16'h00E7; B = 16'h00B; #100;
A = 16'h00E7; B = 16'h00C; #100;
A = 16'h00E7; B = 16'h00D; #100;
A = 16'h00E7; B = 16'h00E; #100;
A = 16'h00E7; B = 16'h00F; #100;
A = 16'h00E7; B = 16'h0010; #100;
A = 16'h00E7; B = 16'h0011; #100;
A = 16'h00E7; B = 16'h0012; #100;
A = 16'h00E7; B = 16'h0013; #100;
A = 16'h00E7; B = 16'h0014; #100;
A = 16'h00E7; B = 16'h0015; #100;
A = 16'h00E7; B = 16'h0016; #100;
A = 16'h00E7; B = 16'h0017; #100;
A = 16'h00E7; B = 16'h0018; #100;
A = 16'h00E7; B = 16'h0019; #100;
A = 16'h00E7; B = 16'h001A; #100;
A = 16'h00E7; B = 16'h001B; #100;
A = 16'h00E7; B = 16'h001C; #100;
A = 16'h00E7; B = 16'h001D; #100;
A = 16'h00E7; B = 16'h001E; #100;
A = 16'h00E7; B = 16'h001F; #100;
A = 16'h00E7; B = 16'h0020; #100;
A = 16'h00E7; B = 16'h0021; #100;
A = 16'h00E7; B = 16'h0022; #100;
A = 16'h00E7; B = 16'h0023; #100;
A = 16'h00E7; B = 16'h0024; #100;
A = 16'h00E7; B = 16'h0025; #100;
A = 16'h00E7; B = 16'h0026; #100;
A = 16'h00E7; B = 16'h0027; #100;
A = 16'h00E7; B = 16'h0028; #100;
A = 16'h00E7; B = 16'h0029; #100;
A = 16'h00E7; B = 16'h002A; #100;
A = 16'h00E7; B = 16'h002B; #100;
A = 16'h00E7; B = 16'h002C; #100;
A = 16'h00E7; B = 16'h002D; #100;
A = 16'h00E7; B = 16'h002E; #100;
A = 16'h00E7; B = 16'h002F; #100;
A = 16'h00E7; B = 16'h0030; #100;
A = 16'h00E7; B = 16'h0031; #100;
A = 16'h00E7; B = 16'h0032; #100;
A = 16'h00E7; B = 16'h0033; #100;
A = 16'h00E7; B = 16'h0034; #100;
A = 16'h00E7; B = 16'h0035; #100;
A = 16'h00E7; B = 16'h0036; #100;
A = 16'h00E7; B = 16'h0037; #100;
A = 16'h00E7; B = 16'h0038; #100;
A = 16'h00E7; B = 16'h0039; #100;
A = 16'h00E7; B = 16'h003A; #100;
A = 16'h00E7; B = 16'h003B; #100;
A = 16'h00E7; B = 16'h003C; #100;
A = 16'h00E7; B = 16'h003D; #100;
A = 16'h00E7; B = 16'h003E; #100;
A = 16'h00E7; B = 16'h003F; #100;
A = 16'h00E7; B = 16'h0040; #100;
A = 16'h00E7; B = 16'h0041; #100;
A = 16'h00E7; B = 16'h0042; #100;
A = 16'h00E7; B = 16'h0043; #100;
A = 16'h00E7; B = 16'h0044; #100;
A = 16'h00E7; B = 16'h0045; #100;
A = 16'h00E7; B = 16'h0046; #100;
A = 16'h00E7; B = 16'h0047; #100;
A = 16'h00E7; B = 16'h0048; #100;
A = 16'h00E7; B = 16'h0049; #100;
A = 16'h00E7; B = 16'h004A; #100;
A = 16'h00E7; B = 16'h004B; #100;
A = 16'h00E7; B = 16'h004C; #100;
A = 16'h00E7; B = 16'h004D; #100;
A = 16'h00E7; B = 16'h004E; #100;
A = 16'h00E7; B = 16'h004F; #100;
A = 16'h00E7; B = 16'h0050; #100;
A = 16'h00E7; B = 16'h0051; #100;
A = 16'h00E7; B = 16'h0052; #100;
A = 16'h00E7; B = 16'h0053; #100;
A = 16'h00E7; B = 16'h0054; #100;
A = 16'h00E7; B = 16'h0055; #100;
A = 16'h00E7; B = 16'h0056; #100;
A = 16'h00E7; B = 16'h0057; #100;
A = 16'h00E7; B = 16'h0058; #100;
A = 16'h00E7; B = 16'h0059; #100;
A = 16'h00E7; B = 16'h005A; #100;
A = 16'h00E7; B = 16'h005B; #100;
A = 16'h00E7; B = 16'h005C; #100;
A = 16'h00E7; B = 16'h005D; #100;
A = 16'h00E7; B = 16'h005E; #100;
A = 16'h00E7; B = 16'h005F; #100;
A = 16'h00E7; B = 16'h0060; #100;
A = 16'h00E7; B = 16'h0061; #100;
A = 16'h00E7; B = 16'h0062; #100;
A = 16'h00E7; B = 16'h0063; #100;
A = 16'h00E7; B = 16'h0064; #100;
A = 16'h00E7; B = 16'h0065; #100;
A = 16'h00E7; B = 16'h0066; #100;
A = 16'h00E7; B = 16'h0067; #100;
A = 16'h00E7; B = 16'h0068; #100;
A = 16'h00E7; B = 16'h0069; #100;
A = 16'h00E7; B = 16'h006A; #100;
A = 16'h00E7; B = 16'h006B; #100;
A = 16'h00E7; B = 16'h006C; #100;
A = 16'h00E7; B = 16'h006D; #100;
A = 16'h00E7; B = 16'h006E; #100;
A = 16'h00E7; B = 16'h006F; #100;
A = 16'h00E7; B = 16'h0070; #100;
A = 16'h00E7; B = 16'h0071; #100;
A = 16'h00E7; B = 16'h0072; #100;
A = 16'h00E7; B = 16'h0073; #100;
A = 16'h00E7; B = 16'h0074; #100;
A = 16'h00E7; B = 16'h0075; #100;
A = 16'h00E7; B = 16'h0076; #100;
A = 16'h00E7; B = 16'h0077; #100;
A = 16'h00E7; B = 16'h0078; #100;
A = 16'h00E7; B = 16'h0079; #100;
A = 16'h00E7; B = 16'h007A; #100;
A = 16'h00E7; B = 16'h007B; #100;
A = 16'h00E7; B = 16'h007C; #100;
A = 16'h00E7; B = 16'h007D; #100;
A = 16'h00E7; B = 16'h007E; #100;
A = 16'h00E7; B = 16'h007F; #100;
A = 16'h00E7; B = 16'h0080; #100;
A = 16'h00E7; B = 16'h0081; #100;
A = 16'h00E7; B = 16'h0082; #100;
A = 16'h00E7; B = 16'h0083; #100;
A = 16'h00E7; B = 16'h0084; #100;
A = 16'h00E7; B = 16'h0085; #100;
A = 16'h00E7; B = 16'h0086; #100;
A = 16'h00E7; B = 16'h0087; #100;
A = 16'h00E7; B = 16'h0088; #100;
A = 16'h00E7; B = 16'h0089; #100;
A = 16'h00E7; B = 16'h008A; #100;
A = 16'h00E7; B = 16'h008B; #100;
A = 16'h00E7; B = 16'h008C; #100;
A = 16'h00E7; B = 16'h008D; #100;
A = 16'h00E7; B = 16'h008E; #100;
A = 16'h00E7; B = 16'h008F; #100;
A = 16'h00E7; B = 16'h0090; #100;
A = 16'h00E7; B = 16'h0091; #100;
A = 16'h00E7; B = 16'h0092; #100;
A = 16'h00E7; B = 16'h0093; #100;
A = 16'h00E7; B = 16'h0094; #100;
A = 16'h00E7; B = 16'h0095; #100;
A = 16'h00E7; B = 16'h0096; #100;
A = 16'h00E7; B = 16'h0097; #100;
A = 16'h00E7; B = 16'h0098; #100;
A = 16'h00E7; B = 16'h0099; #100;
A = 16'h00E7; B = 16'h009A; #100;
A = 16'h00E7; B = 16'h009B; #100;
A = 16'h00E7; B = 16'h009C; #100;
A = 16'h00E7; B = 16'h009D; #100;
A = 16'h00E7; B = 16'h009E; #100;
A = 16'h00E7; B = 16'h009F; #100;
A = 16'h00E7; B = 16'h00A0; #100;
A = 16'h00E7; B = 16'h00A1; #100;
A = 16'h00E7; B = 16'h00A2; #100;
A = 16'h00E7; B = 16'h00A3; #100;
A = 16'h00E7; B = 16'h00A4; #100;
A = 16'h00E7; B = 16'h00A5; #100;
A = 16'h00E7; B = 16'h00A6; #100;
A = 16'h00E7; B = 16'h00A7; #100;
A = 16'h00E7; B = 16'h00A8; #100;
A = 16'h00E7; B = 16'h00A9; #100;
A = 16'h00E7; B = 16'h00AA; #100;
A = 16'h00E7; B = 16'h00AB; #100;
A = 16'h00E7; B = 16'h00AC; #100;
A = 16'h00E7; B = 16'h00AD; #100;
A = 16'h00E7; B = 16'h00AE; #100;
A = 16'h00E7; B = 16'h00AF; #100;
A = 16'h00E7; B = 16'h00B0; #100;
A = 16'h00E7; B = 16'h00B1; #100;
A = 16'h00E7; B = 16'h00B2; #100;
A = 16'h00E7; B = 16'h00B3; #100;
A = 16'h00E7; B = 16'h00B4; #100;
A = 16'h00E7; B = 16'h00B5; #100;
A = 16'h00E7; B = 16'h00B6; #100;
A = 16'h00E7; B = 16'h00B7; #100;
A = 16'h00E7; B = 16'h00B8; #100;
A = 16'h00E7; B = 16'h00B9; #100;
A = 16'h00E7; B = 16'h00BA; #100;
A = 16'h00E7; B = 16'h00BB; #100;
A = 16'h00E7; B = 16'h00BC; #100;
A = 16'h00E7; B = 16'h00BD; #100;
A = 16'h00E7; B = 16'h00BE; #100;
A = 16'h00E7; B = 16'h00BF; #100;
A = 16'h00E7; B = 16'h00C0; #100;
A = 16'h00E7; B = 16'h00C1; #100;
A = 16'h00E7; B = 16'h00C2; #100;
A = 16'h00E7; B = 16'h00C3; #100;
A = 16'h00E7; B = 16'h00C4; #100;
A = 16'h00E7; B = 16'h00C5; #100;
A = 16'h00E7; B = 16'h00C6; #100;
A = 16'h00E7; B = 16'h00C7; #100;
A = 16'h00E7; B = 16'h00C8; #100;
A = 16'h00E7; B = 16'h00C9; #100;
A = 16'h00E7; B = 16'h00CA; #100;
A = 16'h00E7; B = 16'h00CB; #100;
A = 16'h00E7; B = 16'h00CC; #100;
A = 16'h00E7; B = 16'h00CD; #100;
A = 16'h00E7; B = 16'h00CE; #100;
A = 16'h00E7; B = 16'h00CF; #100;
A = 16'h00E7; B = 16'h00D0; #100;
A = 16'h00E7; B = 16'h00D1; #100;
A = 16'h00E7; B = 16'h00D2; #100;
A = 16'h00E7; B = 16'h00D3; #100;
A = 16'h00E7; B = 16'h00D4; #100;
A = 16'h00E7; B = 16'h00D5; #100;
A = 16'h00E7; B = 16'h00D6; #100;
A = 16'h00E7; B = 16'h00D7; #100;
A = 16'h00E7; B = 16'h00D8; #100;
A = 16'h00E7; B = 16'h00D9; #100;
A = 16'h00E7; B = 16'h00DA; #100;
A = 16'h00E7; B = 16'h00DB; #100;
A = 16'h00E7; B = 16'h00DC; #100;
A = 16'h00E7; B = 16'h00DD; #100;
A = 16'h00E7; B = 16'h00DE; #100;
A = 16'h00E7; B = 16'h00DF; #100;
A = 16'h00E7; B = 16'h00E0; #100;
A = 16'h00E7; B = 16'h00E1; #100;
A = 16'h00E7; B = 16'h00E2; #100;
A = 16'h00E7; B = 16'h00E3; #100;
A = 16'h00E7; B = 16'h00E4; #100;
A = 16'h00E7; B = 16'h00E5; #100;
A = 16'h00E7; B = 16'h00E6; #100;
A = 16'h00E7; B = 16'h00E7; #100;
A = 16'h00E7; B = 16'h00E8; #100;
A = 16'h00E7; B = 16'h00E9; #100;
A = 16'h00E7; B = 16'h00EA; #100;
A = 16'h00E7; B = 16'h00EB; #100;
A = 16'h00E7; B = 16'h00EC; #100;
A = 16'h00E7; B = 16'h00ED; #100;
A = 16'h00E7; B = 16'h00EE; #100;
A = 16'h00E7; B = 16'h00EF; #100;
A = 16'h00E7; B = 16'h00F0; #100;
A = 16'h00E7; B = 16'h00F1; #100;
A = 16'h00E7; B = 16'h00F2; #100;
A = 16'h00E7; B = 16'h00F3; #100;
A = 16'h00E7; B = 16'h00F4; #100;
A = 16'h00E7; B = 16'h00F5; #100;
A = 16'h00E7; B = 16'h00F6; #100;
A = 16'h00E7; B = 16'h00F7; #100;
A = 16'h00E7; B = 16'h00F8; #100;
A = 16'h00E7; B = 16'h00F9; #100;
A = 16'h00E7; B = 16'h00FA; #100;
A = 16'h00E7; B = 16'h00FB; #100;
A = 16'h00E7; B = 16'h00FC; #100;
A = 16'h00E7; B = 16'h00FD; #100;
A = 16'h00E7; B = 16'h00FE; #100;
A = 16'h00E7; B = 16'h00FF; #100;
A = 16'h00E8; B = 16'h000; #100;
A = 16'h00E8; B = 16'h001; #100;
A = 16'h00E8; B = 16'h002; #100;
A = 16'h00E8; B = 16'h003; #100;
A = 16'h00E8; B = 16'h004; #100;
A = 16'h00E8; B = 16'h005; #100;
A = 16'h00E8; B = 16'h006; #100;
A = 16'h00E8; B = 16'h007; #100;
A = 16'h00E8; B = 16'h008; #100;
A = 16'h00E8; B = 16'h009; #100;
A = 16'h00E8; B = 16'h00A; #100;
A = 16'h00E8; B = 16'h00B; #100;
A = 16'h00E8; B = 16'h00C; #100;
A = 16'h00E8; B = 16'h00D; #100;
A = 16'h00E8; B = 16'h00E; #100;
A = 16'h00E8; B = 16'h00F; #100;
A = 16'h00E8; B = 16'h0010; #100;
A = 16'h00E8; B = 16'h0011; #100;
A = 16'h00E8; B = 16'h0012; #100;
A = 16'h00E8; B = 16'h0013; #100;
A = 16'h00E8; B = 16'h0014; #100;
A = 16'h00E8; B = 16'h0015; #100;
A = 16'h00E8; B = 16'h0016; #100;
A = 16'h00E8; B = 16'h0017; #100;
A = 16'h00E8; B = 16'h0018; #100;
A = 16'h00E8; B = 16'h0019; #100;
A = 16'h00E8; B = 16'h001A; #100;
A = 16'h00E8; B = 16'h001B; #100;
A = 16'h00E8; B = 16'h001C; #100;
A = 16'h00E8; B = 16'h001D; #100;
A = 16'h00E8; B = 16'h001E; #100;
A = 16'h00E8; B = 16'h001F; #100;
A = 16'h00E8; B = 16'h0020; #100;
A = 16'h00E8; B = 16'h0021; #100;
A = 16'h00E8; B = 16'h0022; #100;
A = 16'h00E8; B = 16'h0023; #100;
A = 16'h00E8; B = 16'h0024; #100;
A = 16'h00E8; B = 16'h0025; #100;
A = 16'h00E8; B = 16'h0026; #100;
A = 16'h00E8; B = 16'h0027; #100;
A = 16'h00E8; B = 16'h0028; #100;
A = 16'h00E8; B = 16'h0029; #100;
A = 16'h00E8; B = 16'h002A; #100;
A = 16'h00E8; B = 16'h002B; #100;
A = 16'h00E8; B = 16'h002C; #100;
A = 16'h00E8; B = 16'h002D; #100;
A = 16'h00E8; B = 16'h002E; #100;
A = 16'h00E8; B = 16'h002F; #100;
A = 16'h00E8; B = 16'h0030; #100;
A = 16'h00E8; B = 16'h0031; #100;
A = 16'h00E8; B = 16'h0032; #100;
A = 16'h00E8; B = 16'h0033; #100;
A = 16'h00E8; B = 16'h0034; #100;
A = 16'h00E8; B = 16'h0035; #100;
A = 16'h00E8; B = 16'h0036; #100;
A = 16'h00E8; B = 16'h0037; #100;
A = 16'h00E8; B = 16'h0038; #100;
A = 16'h00E8; B = 16'h0039; #100;
A = 16'h00E8; B = 16'h003A; #100;
A = 16'h00E8; B = 16'h003B; #100;
A = 16'h00E8; B = 16'h003C; #100;
A = 16'h00E8; B = 16'h003D; #100;
A = 16'h00E8; B = 16'h003E; #100;
A = 16'h00E8; B = 16'h003F; #100;
A = 16'h00E8; B = 16'h0040; #100;
A = 16'h00E8; B = 16'h0041; #100;
A = 16'h00E8; B = 16'h0042; #100;
A = 16'h00E8; B = 16'h0043; #100;
A = 16'h00E8; B = 16'h0044; #100;
A = 16'h00E8; B = 16'h0045; #100;
A = 16'h00E8; B = 16'h0046; #100;
A = 16'h00E8; B = 16'h0047; #100;
A = 16'h00E8; B = 16'h0048; #100;
A = 16'h00E8; B = 16'h0049; #100;
A = 16'h00E8; B = 16'h004A; #100;
A = 16'h00E8; B = 16'h004B; #100;
A = 16'h00E8; B = 16'h004C; #100;
A = 16'h00E8; B = 16'h004D; #100;
A = 16'h00E8; B = 16'h004E; #100;
A = 16'h00E8; B = 16'h004F; #100;
A = 16'h00E8; B = 16'h0050; #100;
A = 16'h00E8; B = 16'h0051; #100;
A = 16'h00E8; B = 16'h0052; #100;
A = 16'h00E8; B = 16'h0053; #100;
A = 16'h00E8; B = 16'h0054; #100;
A = 16'h00E8; B = 16'h0055; #100;
A = 16'h00E8; B = 16'h0056; #100;
A = 16'h00E8; B = 16'h0057; #100;
A = 16'h00E8; B = 16'h0058; #100;
A = 16'h00E8; B = 16'h0059; #100;
A = 16'h00E8; B = 16'h005A; #100;
A = 16'h00E8; B = 16'h005B; #100;
A = 16'h00E8; B = 16'h005C; #100;
A = 16'h00E8; B = 16'h005D; #100;
A = 16'h00E8; B = 16'h005E; #100;
A = 16'h00E8; B = 16'h005F; #100;
A = 16'h00E8; B = 16'h0060; #100;
A = 16'h00E8; B = 16'h0061; #100;
A = 16'h00E8; B = 16'h0062; #100;
A = 16'h00E8; B = 16'h0063; #100;
A = 16'h00E8; B = 16'h0064; #100;
A = 16'h00E8; B = 16'h0065; #100;
A = 16'h00E8; B = 16'h0066; #100;
A = 16'h00E8; B = 16'h0067; #100;
A = 16'h00E8; B = 16'h0068; #100;
A = 16'h00E8; B = 16'h0069; #100;
A = 16'h00E8; B = 16'h006A; #100;
A = 16'h00E8; B = 16'h006B; #100;
A = 16'h00E8; B = 16'h006C; #100;
A = 16'h00E8; B = 16'h006D; #100;
A = 16'h00E8; B = 16'h006E; #100;
A = 16'h00E8; B = 16'h006F; #100;
A = 16'h00E8; B = 16'h0070; #100;
A = 16'h00E8; B = 16'h0071; #100;
A = 16'h00E8; B = 16'h0072; #100;
A = 16'h00E8; B = 16'h0073; #100;
A = 16'h00E8; B = 16'h0074; #100;
A = 16'h00E8; B = 16'h0075; #100;
A = 16'h00E8; B = 16'h0076; #100;
A = 16'h00E8; B = 16'h0077; #100;
A = 16'h00E8; B = 16'h0078; #100;
A = 16'h00E8; B = 16'h0079; #100;
A = 16'h00E8; B = 16'h007A; #100;
A = 16'h00E8; B = 16'h007B; #100;
A = 16'h00E8; B = 16'h007C; #100;
A = 16'h00E8; B = 16'h007D; #100;
A = 16'h00E8; B = 16'h007E; #100;
A = 16'h00E8; B = 16'h007F; #100;
A = 16'h00E8; B = 16'h0080; #100;
A = 16'h00E8; B = 16'h0081; #100;
A = 16'h00E8; B = 16'h0082; #100;
A = 16'h00E8; B = 16'h0083; #100;
A = 16'h00E8; B = 16'h0084; #100;
A = 16'h00E8; B = 16'h0085; #100;
A = 16'h00E8; B = 16'h0086; #100;
A = 16'h00E8; B = 16'h0087; #100;
A = 16'h00E8; B = 16'h0088; #100;
A = 16'h00E8; B = 16'h0089; #100;
A = 16'h00E8; B = 16'h008A; #100;
A = 16'h00E8; B = 16'h008B; #100;
A = 16'h00E8; B = 16'h008C; #100;
A = 16'h00E8; B = 16'h008D; #100;
A = 16'h00E8; B = 16'h008E; #100;
A = 16'h00E8; B = 16'h008F; #100;
A = 16'h00E8; B = 16'h0090; #100;
A = 16'h00E8; B = 16'h0091; #100;
A = 16'h00E8; B = 16'h0092; #100;
A = 16'h00E8; B = 16'h0093; #100;
A = 16'h00E8; B = 16'h0094; #100;
A = 16'h00E8; B = 16'h0095; #100;
A = 16'h00E8; B = 16'h0096; #100;
A = 16'h00E8; B = 16'h0097; #100;
A = 16'h00E8; B = 16'h0098; #100;
A = 16'h00E8; B = 16'h0099; #100;
A = 16'h00E8; B = 16'h009A; #100;
A = 16'h00E8; B = 16'h009B; #100;
A = 16'h00E8; B = 16'h009C; #100;
A = 16'h00E8; B = 16'h009D; #100;
A = 16'h00E8; B = 16'h009E; #100;
A = 16'h00E8; B = 16'h009F; #100;
A = 16'h00E8; B = 16'h00A0; #100;
A = 16'h00E8; B = 16'h00A1; #100;
A = 16'h00E8; B = 16'h00A2; #100;
A = 16'h00E8; B = 16'h00A3; #100;
A = 16'h00E8; B = 16'h00A4; #100;
A = 16'h00E8; B = 16'h00A5; #100;
A = 16'h00E8; B = 16'h00A6; #100;
A = 16'h00E8; B = 16'h00A7; #100;
A = 16'h00E8; B = 16'h00A8; #100;
A = 16'h00E8; B = 16'h00A9; #100;
A = 16'h00E8; B = 16'h00AA; #100;
A = 16'h00E8; B = 16'h00AB; #100;
A = 16'h00E8; B = 16'h00AC; #100;
A = 16'h00E8; B = 16'h00AD; #100;
A = 16'h00E8; B = 16'h00AE; #100;
A = 16'h00E8; B = 16'h00AF; #100;
A = 16'h00E8; B = 16'h00B0; #100;
A = 16'h00E8; B = 16'h00B1; #100;
A = 16'h00E8; B = 16'h00B2; #100;
A = 16'h00E8; B = 16'h00B3; #100;
A = 16'h00E8; B = 16'h00B4; #100;
A = 16'h00E8; B = 16'h00B5; #100;
A = 16'h00E8; B = 16'h00B6; #100;
A = 16'h00E8; B = 16'h00B7; #100;
A = 16'h00E8; B = 16'h00B8; #100;
A = 16'h00E8; B = 16'h00B9; #100;
A = 16'h00E8; B = 16'h00BA; #100;
A = 16'h00E8; B = 16'h00BB; #100;
A = 16'h00E8; B = 16'h00BC; #100;
A = 16'h00E8; B = 16'h00BD; #100;
A = 16'h00E8; B = 16'h00BE; #100;
A = 16'h00E8; B = 16'h00BF; #100;
A = 16'h00E8; B = 16'h00C0; #100;
A = 16'h00E8; B = 16'h00C1; #100;
A = 16'h00E8; B = 16'h00C2; #100;
A = 16'h00E8; B = 16'h00C3; #100;
A = 16'h00E8; B = 16'h00C4; #100;
A = 16'h00E8; B = 16'h00C5; #100;
A = 16'h00E8; B = 16'h00C6; #100;
A = 16'h00E8; B = 16'h00C7; #100;
A = 16'h00E8; B = 16'h00C8; #100;
A = 16'h00E8; B = 16'h00C9; #100;
A = 16'h00E8; B = 16'h00CA; #100;
A = 16'h00E8; B = 16'h00CB; #100;
A = 16'h00E8; B = 16'h00CC; #100;
A = 16'h00E8; B = 16'h00CD; #100;
A = 16'h00E8; B = 16'h00CE; #100;
A = 16'h00E8; B = 16'h00CF; #100;
A = 16'h00E8; B = 16'h00D0; #100;
A = 16'h00E8; B = 16'h00D1; #100;
A = 16'h00E8; B = 16'h00D2; #100;
A = 16'h00E8; B = 16'h00D3; #100;
A = 16'h00E8; B = 16'h00D4; #100;
A = 16'h00E8; B = 16'h00D5; #100;
A = 16'h00E8; B = 16'h00D6; #100;
A = 16'h00E8; B = 16'h00D7; #100;
A = 16'h00E8; B = 16'h00D8; #100;
A = 16'h00E8; B = 16'h00D9; #100;
A = 16'h00E8; B = 16'h00DA; #100;
A = 16'h00E8; B = 16'h00DB; #100;
A = 16'h00E8; B = 16'h00DC; #100;
A = 16'h00E8; B = 16'h00DD; #100;
A = 16'h00E8; B = 16'h00DE; #100;
A = 16'h00E8; B = 16'h00DF; #100;
A = 16'h00E8; B = 16'h00E0; #100;
A = 16'h00E8; B = 16'h00E1; #100;
A = 16'h00E8; B = 16'h00E2; #100;
A = 16'h00E8; B = 16'h00E3; #100;
A = 16'h00E8; B = 16'h00E4; #100;
A = 16'h00E8; B = 16'h00E5; #100;
A = 16'h00E8; B = 16'h00E6; #100;
A = 16'h00E8; B = 16'h00E7; #100;
A = 16'h00E8; B = 16'h00E8; #100;
A = 16'h00E8; B = 16'h00E9; #100;
A = 16'h00E8; B = 16'h00EA; #100;
A = 16'h00E8; B = 16'h00EB; #100;
A = 16'h00E8; B = 16'h00EC; #100;
A = 16'h00E8; B = 16'h00ED; #100;
A = 16'h00E8; B = 16'h00EE; #100;
A = 16'h00E8; B = 16'h00EF; #100;
A = 16'h00E8; B = 16'h00F0; #100;
A = 16'h00E8; B = 16'h00F1; #100;
A = 16'h00E8; B = 16'h00F2; #100;
A = 16'h00E8; B = 16'h00F3; #100;
A = 16'h00E8; B = 16'h00F4; #100;
A = 16'h00E8; B = 16'h00F5; #100;
A = 16'h00E8; B = 16'h00F6; #100;
A = 16'h00E8; B = 16'h00F7; #100;
A = 16'h00E8; B = 16'h00F8; #100;
A = 16'h00E8; B = 16'h00F9; #100;
A = 16'h00E8; B = 16'h00FA; #100;
A = 16'h00E8; B = 16'h00FB; #100;
A = 16'h00E8; B = 16'h00FC; #100;
A = 16'h00E8; B = 16'h00FD; #100;
A = 16'h00E8; B = 16'h00FE; #100;
A = 16'h00E8; B = 16'h00FF; #100;
A = 16'h00E9; B = 16'h000; #100;
A = 16'h00E9; B = 16'h001; #100;
A = 16'h00E9; B = 16'h002; #100;
A = 16'h00E9; B = 16'h003; #100;
A = 16'h00E9; B = 16'h004; #100;
A = 16'h00E9; B = 16'h005; #100;
A = 16'h00E9; B = 16'h006; #100;
A = 16'h00E9; B = 16'h007; #100;
A = 16'h00E9; B = 16'h008; #100;
A = 16'h00E9; B = 16'h009; #100;
A = 16'h00E9; B = 16'h00A; #100;
A = 16'h00E9; B = 16'h00B; #100;
A = 16'h00E9; B = 16'h00C; #100;
A = 16'h00E9; B = 16'h00D; #100;
A = 16'h00E9; B = 16'h00E; #100;
A = 16'h00E9; B = 16'h00F; #100;
A = 16'h00E9; B = 16'h0010; #100;
A = 16'h00E9; B = 16'h0011; #100;
A = 16'h00E9; B = 16'h0012; #100;
A = 16'h00E9; B = 16'h0013; #100;
A = 16'h00E9; B = 16'h0014; #100;
A = 16'h00E9; B = 16'h0015; #100;
A = 16'h00E9; B = 16'h0016; #100;
A = 16'h00E9; B = 16'h0017; #100;
A = 16'h00E9; B = 16'h0018; #100;
A = 16'h00E9; B = 16'h0019; #100;
A = 16'h00E9; B = 16'h001A; #100;
A = 16'h00E9; B = 16'h001B; #100;
A = 16'h00E9; B = 16'h001C; #100;
A = 16'h00E9; B = 16'h001D; #100;
A = 16'h00E9; B = 16'h001E; #100;
A = 16'h00E9; B = 16'h001F; #100;
A = 16'h00E9; B = 16'h0020; #100;
A = 16'h00E9; B = 16'h0021; #100;
A = 16'h00E9; B = 16'h0022; #100;
A = 16'h00E9; B = 16'h0023; #100;
A = 16'h00E9; B = 16'h0024; #100;
A = 16'h00E9; B = 16'h0025; #100;
A = 16'h00E9; B = 16'h0026; #100;
A = 16'h00E9; B = 16'h0027; #100;
A = 16'h00E9; B = 16'h0028; #100;
A = 16'h00E9; B = 16'h0029; #100;
A = 16'h00E9; B = 16'h002A; #100;
A = 16'h00E9; B = 16'h002B; #100;
A = 16'h00E9; B = 16'h002C; #100;
A = 16'h00E9; B = 16'h002D; #100;
A = 16'h00E9; B = 16'h002E; #100;
A = 16'h00E9; B = 16'h002F; #100;
A = 16'h00E9; B = 16'h0030; #100;
A = 16'h00E9; B = 16'h0031; #100;
A = 16'h00E9; B = 16'h0032; #100;
A = 16'h00E9; B = 16'h0033; #100;
A = 16'h00E9; B = 16'h0034; #100;
A = 16'h00E9; B = 16'h0035; #100;
A = 16'h00E9; B = 16'h0036; #100;
A = 16'h00E9; B = 16'h0037; #100;
A = 16'h00E9; B = 16'h0038; #100;
A = 16'h00E9; B = 16'h0039; #100;
A = 16'h00E9; B = 16'h003A; #100;
A = 16'h00E9; B = 16'h003B; #100;
A = 16'h00E9; B = 16'h003C; #100;
A = 16'h00E9; B = 16'h003D; #100;
A = 16'h00E9; B = 16'h003E; #100;
A = 16'h00E9; B = 16'h003F; #100;
A = 16'h00E9; B = 16'h0040; #100;
A = 16'h00E9; B = 16'h0041; #100;
A = 16'h00E9; B = 16'h0042; #100;
A = 16'h00E9; B = 16'h0043; #100;
A = 16'h00E9; B = 16'h0044; #100;
A = 16'h00E9; B = 16'h0045; #100;
A = 16'h00E9; B = 16'h0046; #100;
A = 16'h00E9; B = 16'h0047; #100;
A = 16'h00E9; B = 16'h0048; #100;
A = 16'h00E9; B = 16'h0049; #100;
A = 16'h00E9; B = 16'h004A; #100;
A = 16'h00E9; B = 16'h004B; #100;
A = 16'h00E9; B = 16'h004C; #100;
A = 16'h00E9; B = 16'h004D; #100;
A = 16'h00E9; B = 16'h004E; #100;
A = 16'h00E9; B = 16'h004F; #100;
A = 16'h00E9; B = 16'h0050; #100;
A = 16'h00E9; B = 16'h0051; #100;
A = 16'h00E9; B = 16'h0052; #100;
A = 16'h00E9; B = 16'h0053; #100;
A = 16'h00E9; B = 16'h0054; #100;
A = 16'h00E9; B = 16'h0055; #100;
A = 16'h00E9; B = 16'h0056; #100;
A = 16'h00E9; B = 16'h0057; #100;
A = 16'h00E9; B = 16'h0058; #100;
A = 16'h00E9; B = 16'h0059; #100;
A = 16'h00E9; B = 16'h005A; #100;
A = 16'h00E9; B = 16'h005B; #100;
A = 16'h00E9; B = 16'h005C; #100;
A = 16'h00E9; B = 16'h005D; #100;
A = 16'h00E9; B = 16'h005E; #100;
A = 16'h00E9; B = 16'h005F; #100;
A = 16'h00E9; B = 16'h0060; #100;
A = 16'h00E9; B = 16'h0061; #100;
A = 16'h00E9; B = 16'h0062; #100;
A = 16'h00E9; B = 16'h0063; #100;
A = 16'h00E9; B = 16'h0064; #100;
A = 16'h00E9; B = 16'h0065; #100;
A = 16'h00E9; B = 16'h0066; #100;
A = 16'h00E9; B = 16'h0067; #100;
A = 16'h00E9; B = 16'h0068; #100;
A = 16'h00E9; B = 16'h0069; #100;
A = 16'h00E9; B = 16'h006A; #100;
A = 16'h00E9; B = 16'h006B; #100;
A = 16'h00E9; B = 16'h006C; #100;
A = 16'h00E9; B = 16'h006D; #100;
A = 16'h00E9; B = 16'h006E; #100;
A = 16'h00E9; B = 16'h006F; #100;
A = 16'h00E9; B = 16'h0070; #100;
A = 16'h00E9; B = 16'h0071; #100;
A = 16'h00E9; B = 16'h0072; #100;
A = 16'h00E9; B = 16'h0073; #100;
A = 16'h00E9; B = 16'h0074; #100;
A = 16'h00E9; B = 16'h0075; #100;
A = 16'h00E9; B = 16'h0076; #100;
A = 16'h00E9; B = 16'h0077; #100;
A = 16'h00E9; B = 16'h0078; #100;
A = 16'h00E9; B = 16'h0079; #100;
A = 16'h00E9; B = 16'h007A; #100;
A = 16'h00E9; B = 16'h007B; #100;
A = 16'h00E9; B = 16'h007C; #100;
A = 16'h00E9; B = 16'h007D; #100;
A = 16'h00E9; B = 16'h007E; #100;
A = 16'h00E9; B = 16'h007F; #100;
A = 16'h00E9; B = 16'h0080; #100;
A = 16'h00E9; B = 16'h0081; #100;
A = 16'h00E9; B = 16'h0082; #100;
A = 16'h00E9; B = 16'h0083; #100;
A = 16'h00E9; B = 16'h0084; #100;
A = 16'h00E9; B = 16'h0085; #100;
A = 16'h00E9; B = 16'h0086; #100;
A = 16'h00E9; B = 16'h0087; #100;
A = 16'h00E9; B = 16'h0088; #100;
A = 16'h00E9; B = 16'h0089; #100;
A = 16'h00E9; B = 16'h008A; #100;
A = 16'h00E9; B = 16'h008B; #100;
A = 16'h00E9; B = 16'h008C; #100;
A = 16'h00E9; B = 16'h008D; #100;
A = 16'h00E9; B = 16'h008E; #100;
A = 16'h00E9; B = 16'h008F; #100;
A = 16'h00E9; B = 16'h0090; #100;
A = 16'h00E9; B = 16'h0091; #100;
A = 16'h00E9; B = 16'h0092; #100;
A = 16'h00E9; B = 16'h0093; #100;
A = 16'h00E9; B = 16'h0094; #100;
A = 16'h00E9; B = 16'h0095; #100;
A = 16'h00E9; B = 16'h0096; #100;
A = 16'h00E9; B = 16'h0097; #100;
A = 16'h00E9; B = 16'h0098; #100;
A = 16'h00E9; B = 16'h0099; #100;
A = 16'h00E9; B = 16'h009A; #100;
A = 16'h00E9; B = 16'h009B; #100;
A = 16'h00E9; B = 16'h009C; #100;
A = 16'h00E9; B = 16'h009D; #100;
A = 16'h00E9; B = 16'h009E; #100;
A = 16'h00E9; B = 16'h009F; #100;
A = 16'h00E9; B = 16'h00A0; #100;
A = 16'h00E9; B = 16'h00A1; #100;
A = 16'h00E9; B = 16'h00A2; #100;
A = 16'h00E9; B = 16'h00A3; #100;
A = 16'h00E9; B = 16'h00A4; #100;
A = 16'h00E9; B = 16'h00A5; #100;
A = 16'h00E9; B = 16'h00A6; #100;
A = 16'h00E9; B = 16'h00A7; #100;
A = 16'h00E9; B = 16'h00A8; #100;
A = 16'h00E9; B = 16'h00A9; #100;
A = 16'h00E9; B = 16'h00AA; #100;
A = 16'h00E9; B = 16'h00AB; #100;
A = 16'h00E9; B = 16'h00AC; #100;
A = 16'h00E9; B = 16'h00AD; #100;
A = 16'h00E9; B = 16'h00AE; #100;
A = 16'h00E9; B = 16'h00AF; #100;
A = 16'h00E9; B = 16'h00B0; #100;
A = 16'h00E9; B = 16'h00B1; #100;
A = 16'h00E9; B = 16'h00B2; #100;
A = 16'h00E9; B = 16'h00B3; #100;
A = 16'h00E9; B = 16'h00B4; #100;
A = 16'h00E9; B = 16'h00B5; #100;
A = 16'h00E9; B = 16'h00B6; #100;
A = 16'h00E9; B = 16'h00B7; #100;
A = 16'h00E9; B = 16'h00B8; #100;
A = 16'h00E9; B = 16'h00B9; #100;
A = 16'h00E9; B = 16'h00BA; #100;
A = 16'h00E9; B = 16'h00BB; #100;
A = 16'h00E9; B = 16'h00BC; #100;
A = 16'h00E9; B = 16'h00BD; #100;
A = 16'h00E9; B = 16'h00BE; #100;
A = 16'h00E9; B = 16'h00BF; #100;
A = 16'h00E9; B = 16'h00C0; #100;
A = 16'h00E9; B = 16'h00C1; #100;
A = 16'h00E9; B = 16'h00C2; #100;
A = 16'h00E9; B = 16'h00C3; #100;
A = 16'h00E9; B = 16'h00C4; #100;
A = 16'h00E9; B = 16'h00C5; #100;
A = 16'h00E9; B = 16'h00C6; #100;
A = 16'h00E9; B = 16'h00C7; #100;
A = 16'h00E9; B = 16'h00C8; #100;
A = 16'h00E9; B = 16'h00C9; #100;
A = 16'h00E9; B = 16'h00CA; #100;
A = 16'h00E9; B = 16'h00CB; #100;
A = 16'h00E9; B = 16'h00CC; #100;
A = 16'h00E9; B = 16'h00CD; #100;
A = 16'h00E9; B = 16'h00CE; #100;
A = 16'h00E9; B = 16'h00CF; #100;
A = 16'h00E9; B = 16'h00D0; #100;
A = 16'h00E9; B = 16'h00D1; #100;
A = 16'h00E9; B = 16'h00D2; #100;
A = 16'h00E9; B = 16'h00D3; #100;
A = 16'h00E9; B = 16'h00D4; #100;
A = 16'h00E9; B = 16'h00D5; #100;
A = 16'h00E9; B = 16'h00D6; #100;
A = 16'h00E9; B = 16'h00D7; #100;
A = 16'h00E9; B = 16'h00D8; #100;
A = 16'h00E9; B = 16'h00D9; #100;
A = 16'h00E9; B = 16'h00DA; #100;
A = 16'h00E9; B = 16'h00DB; #100;
A = 16'h00E9; B = 16'h00DC; #100;
A = 16'h00E9; B = 16'h00DD; #100;
A = 16'h00E9; B = 16'h00DE; #100;
A = 16'h00E9; B = 16'h00DF; #100;
A = 16'h00E9; B = 16'h00E0; #100;
A = 16'h00E9; B = 16'h00E1; #100;
A = 16'h00E9; B = 16'h00E2; #100;
A = 16'h00E9; B = 16'h00E3; #100;
A = 16'h00E9; B = 16'h00E4; #100;
A = 16'h00E9; B = 16'h00E5; #100;
A = 16'h00E9; B = 16'h00E6; #100;
A = 16'h00E9; B = 16'h00E7; #100;
A = 16'h00E9; B = 16'h00E8; #100;
A = 16'h00E9; B = 16'h00E9; #100;
A = 16'h00E9; B = 16'h00EA; #100;
A = 16'h00E9; B = 16'h00EB; #100;
A = 16'h00E9; B = 16'h00EC; #100;
A = 16'h00E9; B = 16'h00ED; #100;
A = 16'h00E9; B = 16'h00EE; #100;
A = 16'h00E9; B = 16'h00EF; #100;
A = 16'h00E9; B = 16'h00F0; #100;
A = 16'h00E9; B = 16'h00F1; #100;
A = 16'h00E9; B = 16'h00F2; #100;
A = 16'h00E9; B = 16'h00F3; #100;
A = 16'h00E9; B = 16'h00F4; #100;
A = 16'h00E9; B = 16'h00F5; #100;
A = 16'h00E9; B = 16'h00F6; #100;
A = 16'h00E9; B = 16'h00F7; #100;
A = 16'h00E9; B = 16'h00F8; #100;
A = 16'h00E9; B = 16'h00F9; #100;
A = 16'h00E9; B = 16'h00FA; #100;
A = 16'h00E9; B = 16'h00FB; #100;
A = 16'h00E9; B = 16'h00FC; #100;
A = 16'h00E9; B = 16'h00FD; #100;
A = 16'h00E9; B = 16'h00FE; #100;
A = 16'h00E9; B = 16'h00FF; #100;
A = 16'h00EA; B = 16'h000; #100;
A = 16'h00EA; B = 16'h001; #100;
A = 16'h00EA; B = 16'h002; #100;
A = 16'h00EA; B = 16'h003; #100;
A = 16'h00EA; B = 16'h004; #100;
A = 16'h00EA; B = 16'h005; #100;
A = 16'h00EA; B = 16'h006; #100;
A = 16'h00EA; B = 16'h007; #100;
A = 16'h00EA; B = 16'h008; #100;
A = 16'h00EA; B = 16'h009; #100;
A = 16'h00EA; B = 16'h00A; #100;
A = 16'h00EA; B = 16'h00B; #100;
A = 16'h00EA; B = 16'h00C; #100;
A = 16'h00EA; B = 16'h00D; #100;
A = 16'h00EA; B = 16'h00E; #100;
A = 16'h00EA; B = 16'h00F; #100;
A = 16'h00EA; B = 16'h0010; #100;
A = 16'h00EA; B = 16'h0011; #100;
A = 16'h00EA; B = 16'h0012; #100;
A = 16'h00EA; B = 16'h0013; #100;
A = 16'h00EA; B = 16'h0014; #100;
A = 16'h00EA; B = 16'h0015; #100;
A = 16'h00EA; B = 16'h0016; #100;
A = 16'h00EA; B = 16'h0017; #100;
A = 16'h00EA; B = 16'h0018; #100;
A = 16'h00EA; B = 16'h0019; #100;
A = 16'h00EA; B = 16'h001A; #100;
A = 16'h00EA; B = 16'h001B; #100;
A = 16'h00EA; B = 16'h001C; #100;
A = 16'h00EA; B = 16'h001D; #100;
A = 16'h00EA; B = 16'h001E; #100;
A = 16'h00EA; B = 16'h001F; #100;
A = 16'h00EA; B = 16'h0020; #100;
A = 16'h00EA; B = 16'h0021; #100;
A = 16'h00EA; B = 16'h0022; #100;
A = 16'h00EA; B = 16'h0023; #100;
A = 16'h00EA; B = 16'h0024; #100;
A = 16'h00EA; B = 16'h0025; #100;
A = 16'h00EA; B = 16'h0026; #100;
A = 16'h00EA; B = 16'h0027; #100;
A = 16'h00EA; B = 16'h0028; #100;
A = 16'h00EA; B = 16'h0029; #100;
A = 16'h00EA; B = 16'h002A; #100;
A = 16'h00EA; B = 16'h002B; #100;
A = 16'h00EA; B = 16'h002C; #100;
A = 16'h00EA; B = 16'h002D; #100;
A = 16'h00EA; B = 16'h002E; #100;
A = 16'h00EA; B = 16'h002F; #100;
A = 16'h00EA; B = 16'h0030; #100;
A = 16'h00EA; B = 16'h0031; #100;
A = 16'h00EA; B = 16'h0032; #100;
A = 16'h00EA; B = 16'h0033; #100;
A = 16'h00EA; B = 16'h0034; #100;
A = 16'h00EA; B = 16'h0035; #100;
A = 16'h00EA; B = 16'h0036; #100;
A = 16'h00EA; B = 16'h0037; #100;
A = 16'h00EA; B = 16'h0038; #100;
A = 16'h00EA; B = 16'h0039; #100;
A = 16'h00EA; B = 16'h003A; #100;
A = 16'h00EA; B = 16'h003B; #100;
A = 16'h00EA; B = 16'h003C; #100;
A = 16'h00EA; B = 16'h003D; #100;
A = 16'h00EA; B = 16'h003E; #100;
A = 16'h00EA; B = 16'h003F; #100;
A = 16'h00EA; B = 16'h0040; #100;
A = 16'h00EA; B = 16'h0041; #100;
A = 16'h00EA; B = 16'h0042; #100;
A = 16'h00EA; B = 16'h0043; #100;
A = 16'h00EA; B = 16'h0044; #100;
A = 16'h00EA; B = 16'h0045; #100;
A = 16'h00EA; B = 16'h0046; #100;
A = 16'h00EA; B = 16'h0047; #100;
A = 16'h00EA; B = 16'h0048; #100;
A = 16'h00EA; B = 16'h0049; #100;
A = 16'h00EA; B = 16'h004A; #100;
A = 16'h00EA; B = 16'h004B; #100;
A = 16'h00EA; B = 16'h004C; #100;
A = 16'h00EA; B = 16'h004D; #100;
A = 16'h00EA; B = 16'h004E; #100;
A = 16'h00EA; B = 16'h004F; #100;
A = 16'h00EA; B = 16'h0050; #100;
A = 16'h00EA; B = 16'h0051; #100;
A = 16'h00EA; B = 16'h0052; #100;
A = 16'h00EA; B = 16'h0053; #100;
A = 16'h00EA; B = 16'h0054; #100;
A = 16'h00EA; B = 16'h0055; #100;
A = 16'h00EA; B = 16'h0056; #100;
A = 16'h00EA; B = 16'h0057; #100;
A = 16'h00EA; B = 16'h0058; #100;
A = 16'h00EA; B = 16'h0059; #100;
A = 16'h00EA; B = 16'h005A; #100;
A = 16'h00EA; B = 16'h005B; #100;
A = 16'h00EA; B = 16'h005C; #100;
A = 16'h00EA; B = 16'h005D; #100;
A = 16'h00EA; B = 16'h005E; #100;
A = 16'h00EA; B = 16'h005F; #100;
A = 16'h00EA; B = 16'h0060; #100;
A = 16'h00EA; B = 16'h0061; #100;
A = 16'h00EA; B = 16'h0062; #100;
A = 16'h00EA; B = 16'h0063; #100;
A = 16'h00EA; B = 16'h0064; #100;
A = 16'h00EA; B = 16'h0065; #100;
A = 16'h00EA; B = 16'h0066; #100;
A = 16'h00EA; B = 16'h0067; #100;
A = 16'h00EA; B = 16'h0068; #100;
A = 16'h00EA; B = 16'h0069; #100;
A = 16'h00EA; B = 16'h006A; #100;
A = 16'h00EA; B = 16'h006B; #100;
A = 16'h00EA; B = 16'h006C; #100;
A = 16'h00EA; B = 16'h006D; #100;
A = 16'h00EA; B = 16'h006E; #100;
A = 16'h00EA; B = 16'h006F; #100;
A = 16'h00EA; B = 16'h0070; #100;
A = 16'h00EA; B = 16'h0071; #100;
A = 16'h00EA; B = 16'h0072; #100;
A = 16'h00EA; B = 16'h0073; #100;
A = 16'h00EA; B = 16'h0074; #100;
A = 16'h00EA; B = 16'h0075; #100;
A = 16'h00EA; B = 16'h0076; #100;
A = 16'h00EA; B = 16'h0077; #100;
A = 16'h00EA; B = 16'h0078; #100;
A = 16'h00EA; B = 16'h0079; #100;
A = 16'h00EA; B = 16'h007A; #100;
A = 16'h00EA; B = 16'h007B; #100;
A = 16'h00EA; B = 16'h007C; #100;
A = 16'h00EA; B = 16'h007D; #100;
A = 16'h00EA; B = 16'h007E; #100;
A = 16'h00EA; B = 16'h007F; #100;
A = 16'h00EA; B = 16'h0080; #100;
A = 16'h00EA; B = 16'h0081; #100;
A = 16'h00EA; B = 16'h0082; #100;
A = 16'h00EA; B = 16'h0083; #100;
A = 16'h00EA; B = 16'h0084; #100;
A = 16'h00EA; B = 16'h0085; #100;
A = 16'h00EA; B = 16'h0086; #100;
A = 16'h00EA; B = 16'h0087; #100;
A = 16'h00EA; B = 16'h0088; #100;
A = 16'h00EA; B = 16'h0089; #100;
A = 16'h00EA; B = 16'h008A; #100;
A = 16'h00EA; B = 16'h008B; #100;
A = 16'h00EA; B = 16'h008C; #100;
A = 16'h00EA; B = 16'h008D; #100;
A = 16'h00EA; B = 16'h008E; #100;
A = 16'h00EA; B = 16'h008F; #100;
A = 16'h00EA; B = 16'h0090; #100;
A = 16'h00EA; B = 16'h0091; #100;
A = 16'h00EA; B = 16'h0092; #100;
A = 16'h00EA; B = 16'h0093; #100;
A = 16'h00EA; B = 16'h0094; #100;
A = 16'h00EA; B = 16'h0095; #100;
A = 16'h00EA; B = 16'h0096; #100;
A = 16'h00EA; B = 16'h0097; #100;
A = 16'h00EA; B = 16'h0098; #100;
A = 16'h00EA; B = 16'h0099; #100;
A = 16'h00EA; B = 16'h009A; #100;
A = 16'h00EA; B = 16'h009B; #100;
A = 16'h00EA; B = 16'h009C; #100;
A = 16'h00EA; B = 16'h009D; #100;
A = 16'h00EA; B = 16'h009E; #100;
A = 16'h00EA; B = 16'h009F; #100;
A = 16'h00EA; B = 16'h00A0; #100;
A = 16'h00EA; B = 16'h00A1; #100;
A = 16'h00EA; B = 16'h00A2; #100;
A = 16'h00EA; B = 16'h00A3; #100;
A = 16'h00EA; B = 16'h00A4; #100;
A = 16'h00EA; B = 16'h00A5; #100;
A = 16'h00EA; B = 16'h00A6; #100;
A = 16'h00EA; B = 16'h00A7; #100;
A = 16'h00EA; B = 16'h00A8; #100;
A = 16'h00EA; B = 16'h00A9; #100;
A = 16'h00EA; B = 16'h00AA; #100;
A = 16'h00EA; B = 16'h00AB; #100;
A = 16'h00EA; B = 16'h00AC; #100;
A = 16'h00EA; B = 16'h00AD; #100;
A = 16'h00EA; B = 16'h00AE; #100;
A = 16'h00EA; B = 16'h00AF; #100;
A = 16'h00EA; B = 16'h00B0; #100;
A = 16'h00EA; B = 16'h00B1; #100;
A = 16'h00EA; B = 16'h00B2; #100;
A = 16'h00EA; B = 16'h00B3; #100;
A = 16'h00EA; B = 16'h00B4; #100;
A = 16'h00EA; B = 16'h00B5; #100;
A = 16'h00EA; B = 16'h00B6; #100;
A = 16'h00EA; B = 16'h00B7; #100;
A = 16'h00EA; B = 16'h00B8; #100;
A = 16'h00EA; B = 16'h00B9; #100;
A = 16'h00EA; B = 16'h00BA; #100;
A = 16'h00EA; B = 16'h00BB; #100;
A = 16'h00EA; B = 16'h00BC; #100;
A = 16'h00EA; B = 16'h00BD; #100;
A = 16'h00EA; B = 16'h00BE; #100;
A = 16'h00EA; B = 16'h00BF; #100;
A = 16'h00EA; B = 16'h00C0; #100;
A = 16'h00EA; B = 16'h00C1; #100;
A = 16'h00EA; B = 16'h00C2; #100;
A = 16'h00EA; B = 16'h00C3; #100;
A = 16'h00EA; B = 16'h00C4; #100;
A = 16'h00EA; B = 16'h00C5; #100;
A = 16'h00EA; B = 16'h00C6; #100;
A = 16'h00EA; B = 16'h00C7; #100;
A = 16'h00EA; B = 16'h00C8; #100;
A = 16'h00EA; B = 16'h00C9; #100;
A = 16'h00EA; B = 16'h00CA; #100;
A = 16'h00EA; B = 16'h00CB; #100;
A = 16'h00EA; B = 16'h00CC; #100;
A = 16'h00EA; B = 16'h00CD; #100;
A = 16'h00EA; B = 16'h00CE; #100;
A = 16'h00EA; B = 16'h00CF; #100;
A = 16'h00EA; B = 16'h00D0; #100;
A = 16'h00EA; B = 16'h00D1; #100;
A = 16'h00EA; B = 16'h00D2; #100;
A = 16'h00EA; B = 16'h00D3; #100;
A = 16'h00EA; B = 16'h00D4; #100;
A = 16'h00EA; B = 16'h00D5; #100;
A = 16'h00EA; B = 16'h00D6; #100;
A = 16'h00EA; B = 16'h00D7; #100;
A = 16'h00EA; B = 16'h00D8; #100;
A = 16'h00EA; B = 16'h00D9; #100;
A = 16'h00EA; B = 16'h00DA; #100;
A = 16'h00EA; B = 16'h00DB; #100;
A = 16'h00EA; B = 16'h00DC; #100;
A = 16'h00EA; B = 16'h00DD; #100;
A = 16'h00EA; B = 16'h00DE; #100;
A = 16'h00EA; B = 16'h00DF; #100;
A = 16'h00EA; B = 16'h00E0; #100;
A = 16'h00EA; B = 16'h00E1; #100;
A = 16'h00EA; B = 16'h00E2; #100;
A = 16'h00EA; B = 16'h00E3; #100;
A = 16'h00EA; B = 16'h00E4; #100;
A = 16'h00EA; B = 16'h00E5; #100;
A = 16'h00EA; B = 16'h00E6; #100;
A = 16'h00EA; B = 16'h00E7; #100;
A = 16'h00EA; B = 16'h00E8; #100;
A = 16'h00EA; B = 16'h00E9; #100;
A = 16'h00EA; B = 16'h00EA; #100;
A = 16'h00EA; B = 16'h00EB; #100;
A = 16'h00EA; B = 16'h00EC; #100;
A = 16'h00EA; B = 16'h00ED; #100;
A = 16'h00EA; B = 16'h00EE; #100;
A = 16'h00EA; B = 16'h00EF; #100;
A = 16'h00EA; B = 16'h00F0; #100;
A = 16'h00EA; B = 16'h00F1; #100;
A = 16'h00EA; B = 16'h00F2; #100;
A = 16'h00EA; B = 16'h00F3; #100;
A = 16'h00EA; B = 16'h00F4; #100;
A = 16'h00EA; B = 16'h00F5; #100;
A = 16'h00EA; B = 16'h00F6; #100;
A = 16'h00EA; B = 16'h00F7; #100;
A = 16'h00EA; B = 16'h00F8; #100;
A = 16'h00EA; B = 16'h00F9; #100;
A = 16'h00EA; B = 16'h00FA; #100;
A = 16'h00EA; B = 16'h00FB; #100;
A = 16'h00EA; B = 16'h00FC; #100;
A = 16'h00EA; B = 16'h00FD; #100;
A = 16'h00EA; B = 16'h00FE; #100;
A = 16'h00EA; B = 16'h00FF; #100;
A = 16'h00EB; B = 16'h000; #100;
A = 16'h00EB; B = 16'h001; #100;
A = 16'h00EB; B = 16'h002; #100;
A = 16'h00EB; B = 16'h003; #100;
A = 16'h00EB; B = 16'h004; #100;
A = 16'h00EB; B = 16'h005; #100;
A = 16'h00EB; B = 16'h006; #100;
A = 16'h00EB; B = 16'h007; #100;
A = 16'h00EB; B = 16'h008; #100;
A = 16'h00EB; B = 16'h009; #100;
A = 16'h00EB; B = 16'h00A; #100;
A = 16'h00EB; B = 16'h00B; #100;
A = 16'h00EB; B = 16'h00C; #100;
A = 16'h00EB; B = 16'h00D; #100;
A = 16'h00EB; B = 16'h00E; #100;
A = 16'h00EB; B = 16'h00F; #100;
A = 16'h00EB; B = 16'h0010; #100;
A = 16'h00EB; B = 16'h0011; #100;
A = 16'h00EB; B = 16'h0012; #100;
A = 16'h00EB; B = 16'h0013; #100;
A = 16'h00EB; B = 16'h0014; #100;
A = 16'h00EB; B = 16'h0015; #100;
A = 16'h00EB; B = 16'h0016; #100;
A = 16'h00EB; B = 16'h0017; #100;
A = 16'h00EB; B = 16'h0018; #100;
A = 16'h00EB; B = 16'h0019; #100;
A = 16'h00EB; B = 16'h001A; #100;
A = 16'h00EB; B = 16'h001B; #100;
A = 16'h00EB; B = 16'h001C; #100;
A = 16'h00EB; B = 16'h001D; #100;
A = 16'h00EB; B = 16'h001E; #100;
A = 16'h00EB; B = 16'h001F; #100;
A = 16'h00EB; B = 16'h0020; #100;
A = 16'h00EB; B = 16'h0021; #100;
A = 16'h00EB; B = 16'h0022; #100;
A = 16'h00EB; B = 16'h0023; #100;
A = 16'h00EB; B = 16'h0024; #100;
A = 16'h00EB; B = 16'h0025; #100;
A = 16'h00EB; B = 16'h0026; #100;
A = 16'h00EB; B = 16'h0027; #100;
A = 16'h00EB; B = 16'h0028; #100;
A = 16'h00EB; B = 16'h0029; #100;
A = 16'h00EB; B = 16'h002A; #100;
A = 16'h00EB; B = 16'h002B; #100;
A = 16'h00EB; B = 16'h002C; #100;
A = 16'h00EB; B = 16'h002D; #100;
A = 16'h00EB; B = 16'h002E; #100;
A = 16'h00EB; B = 16'h002F; #100;
A = 16'h00EB; B = 16'h0030; #100;
A = 16'h00EB; B = 16'h0031; #100;
A = 16'h00EB; B = 16'h0032; #100;
A = 16'h00EB; B = 16'h0033; #100;
A = 16'h00EB; B = 16'h0034; #100;
A = 16'h00EB; B = 16'h0035; #100;
A = 16'h00EB; B = 16'h0036; #100;
A = 16'h00EB; B = 16'h0037; #100;
A = 16'h00EB; B = 16'h0038; #100;
A = 16'h00EB; B = 16'h0039; #100;
A = 16'h00EB; B = 16'h003A; #100;
A = 16'h00EB; B = 16'h003B; #100;
A = 16'h00EB; B = 16'h003C; #100;
A = 16'h00EB; B = 16'h003D; #100;
A = 16'h00EB; B = 16'h003E; #100;
A = 16'h00EB; B = 16'h003F; #100;
A = 16'h00EB; B = 16'h0040; #100;
A = 16'h00EB; B = 16'h0041; #100;
A = 16'h00EB; B = 16'h0042; #100;
A = 16'h00EB; B = 16'h0043; #100;
A = 16'h00EB; B = 16'h0044; #100;
A = 16'h00EB; B = 16'h0045; #100;
A = 16'h00EB; B = 16'h0046; #100;
A = 16'h00EB; B = 16'h0047; #100;
A = 16'h00EB; B = 16'h0048; #100;
A = 16'h00EB; B = 16'h0049; #100;
A = 16'h00EB; B = 16'h004A; #100;
A = 16'h00EB; B = 16'h004B; #100;
A = 16'h00EB; B = 16'h004C; #100;
A = 16'h00EB; B = 16'h004D; #100;
A = 16'h00EB; B = 16'h004E; #100;
A = 16'h00EB; B = 16'h004F; #100;
A = 16'h00EB; B = 16'h0050; #100;
A = 16'h00EB; B = 16'h0051; #100;
A = 16'h00EB; B = 16'h0052; #100;
A = 16'h00EB; B = 16'h0053; #100;
A = 16'h00EB; B = 16'h0054; #100;
A = 16'h00EB; B = 16'h0055; #100;
A = 16'h00EB; B = 16'h0056; #100;
A = 16'h00EB; B = 16'h0057; #100;
A = 16'h00EB; B = 16'h0058; #100;
A = 16'h00EB; B = 16'h0059; #100;
A = 16'h00EB; B = 16'h005A; #100;
A = 16'h00EB; B = 16'h005B; #100;
A = 16'h00EB; B = 16'h005C; #100;
A = 16'h00EB; B = 16'h005D; #100;
A = 16'h00EB; B = 16'h005E; #100;
A = 16'h00EB; B = 16'h005F; #100;
A = 16'h00EB; B = 16'h0060; #100;
A = 16'h00EB; B = 16'h0061; #100;
A = 16'h00EB; B = 16'h0062; #100;
A = 16'h00EB; B = 16'h0063; #100;
A = 16'h00EB; B = 16'h0064; #100;
A = 16'h00EB; B = 16'h0065; #100;
A = 16'h00EB; B = 16'h0066; #100;
A = 16'h00EB; B = 16'h0067; #100;
A = 16'h00EB; B = 16'h0068; #100;
A = 16'h00EB; B = 16'h0069; #100;
A = 16'h00EB; B = 16'h006A; #100;
A = 16'h00EB; B = 16'h006B; #100;
A = 16'h00EB; B = 16'h006C; #100;
A = 16'h00EB; B = 16'h006D; #100;
A = 16'h00EB; B = 16'h006E; #100;
A = 16'h00EB; B = 16'h006F; #100;
A = 16'h00EB; B = 16'h0070; #100;
A = 16'h00EB; B = 16'h0071; #100;
A = 16'h00EB; B = 16'h0072; #100;
A = 16'h00EB; B = 16'h0073; #100;
A = 16'h00EB; B = 16'h0074; #100;
A = 16'h00EB; B = 16'h0075; #100;
A = 16'h00EB; B = 16'h0076; #100;
A = 16'h00EB; B = 16'h0077; #100;
A = 16'h00EB; B = 16'h0078; #100;
A = 16'h00EB; B = 16'h0079; #100;
A = 16'h00EB; B = 16'h007A; #100;
A = 16'h00EB; B = 16'h007B; #100;
A = 16'h00EB; B = 16'h007C; #100;
A = 16'h00EB; B = 16'h007D; #100;
A = 16'h00EB; B = 16'h007E; #100;
A = 16'h00EB; B = 16'h007F; #100;
A = 16'h00EB; B = 16'h0080; #100;
A = 16'h00EB; B = 16'h0081; #100;
A = 16'h00EB; B = 16'h0082; #100;
A = 16'h00EB; B = 16'h0083; #100;
A = 16'h00EB; B = 16'h0084; #100;
A = 16'h00EB; B = 16'h0085; #100;
A = 16'h00EB; B = 16'h0086; #100;
A = 16'h00EB; B = 16'h0087; #100;
A = 16'h00EB; B = 16'h0088; #100;
A = 16'h00EB; B = 16'h0089; #100;
A = 16'h00EB; B = 16'h008A; #100;
A = 16'h00EB; B = 16'h008B; #100;
A = 16'h00EB; B = 16'h008C; #100;
A = 16'h00EB; B = 16'h008D; #100;
A = 16'h00EB; B = 16'h008E; #100;
A = 16'h00EB; B = 16'h008F; #100;
A = 16'h00EB; B = 16'h0090; #100;
A = 16'h00EB; B = 16'h0091; #100;
A = 16'h00EB; B = 16'h0092; #100;
A = 16'h00EB; B = 16'h0093; #100;
A = 16'h00EB; B = 16'h0094; #100;
A = 16'h00EB; B = 16'h0095; #100;
A = 16'h00EB; B = 16'h0096; #100;
A = 16'h00EB; B = 16'h0097; #100;
A = 16'h00EB; B = 16'h0098; #100;
A = 16'h00EB; B = 16'h0099; #100;
A = 16'h00EB; B = 16'h009A; #100;
A = 16'h00EB; B = 16'h009B; #100;
A = 16'h00EB; B = 16'h009C; #100;
A = 16'h00EB; B = 16'h009D; #100;
A = 16'h00EB; B = 16'h009E; #100;
A = 16'h00EB; B = 16'h009F; #100;
A = 16'h00EB; B = 16'h00A0; #100;
A = 16'h00EB; B = 16'h00A1; #100;
A = 16'h00EB; B = 16'h00A2; #100;
A = 16'h00EB; B = 16'h00A3; #100;
A = 16'h00EB; B = 16'h00A4; #100;
A = 16'h00EB; B = 16'h00A5; #100;
A = 16'h00EB; B = 16'h00A6; #100;
A = 16'h00EB; B = 16'h00A7; #100;
A = 16'h00EB; B = 16'h00A8; #100;
A = 16'h00EB; B = 16'h00A9; #100;
A = 16'h00EB; B = 16'h00AA; #100;
A = 16'h00EB; B = 16'h00AB; #100;
A = 16'h00EB; B = 16'h00AC; #100;
A = 16'h00EB; B = 16'h00AD; #100;
A = 16'h00EB; B = 16'h00AE; #100;
A = 16'h00EB; B = 16'h00AF; #100;
A = 16'h00EB; B = 16'h00B0; #100;
A = 16'h00EB; B = 16'h00B1; #100;
A = 16'h00EB; B = 16'h00B2; #100;
A = 16'h00EB; B = 16'h00B3; #100;
A = 16'h00EB; B = 16'h00B4; #100;
A = 16'h00EB; B = 16'h00B5; #100;
A = 16'h00EB; B = 16'h00B6; #100;
A = 16'h00EB; B = 16'h00B7; #100;
A = 16'h00EB; B = 16'h00B8; #100;
A = 16'h00EB; B = 16'h00B9; #100;
A = 16'h00EB; B = 16'h00BA; #100;
A = 16'h00EB; B = 16'h00BB; #100;
A = 16'h00EB; B = 16'h00BC; #100;
A = 16'h00EB; B = 16'h00BD; #100;
A = 16'h00EB; B = 16'h00BE; #100;
A = 16'h00EB; B = 16'h00BF; #100;
A = 16'h00EB; B = 16'h00C0; #100;
A = 16'h00EB; B = 16'h00C1; #100;
A = 16'h00EB; B = 16'h00C2; #100;
A = 16'h00EB; B = 16'h00C3; #100;
A = 16'h00EB; B = 16'h00C4; #100;
A = 16'h00EB; B = 16'h00C5; #100;
A = 16'h00EB; B = 16'h00C6; #100;
A = 16'h00EB; B = 16'h00C7; #100;
A = 16'h00EB; B = 16'h00C8; #100;
A = 16'h00EB; B = 16'h00C9; #100;
A = 16'h00EB; B = 16'h00CA; #100;
A = 16'h00EB; B = 16'h00CB; #100;
A = 16'h00EB; B = 16'h00CC; #100;
A = 16'h00EB; B = 16'h00CD; #100;
A = 16'h00EB; B = 16'h00CE; #100;
A = 16'h00EB; B = 16'h00CF; #100;
A = 16'h00EB; B = 16'h00D0; #100;
A = 16'h00EB; B = 16'h00D1; #100;
A = 16'h00EB; B = 16'h00D2; #100;
A = 16'h00EB; B = 16'h00D3; #100;
A = 16'h00EB; B = 16'h00D4; #100;
A = 16'h00EB; B = 16'h00D5; #100;
A = 16'h00EB; B = 16'h00D6; #100;
A = 16'h00EB; B = 16'h00D7; #100;
A = 16'h00EB; B = 16'h00D8; #100;
A = 16'h00EB; B = 16'h00D9; #100;
A = 16'h00EB; B = 16'h00DA; #100;
A = 16'h00EB; B = 16'h00DB; #100;
A = 16'h00EB; B = 16'h00DC; #100;
A = 16'h00EB; B = 16'h00DD; #100;
A = 16'h00EB; B = 16'h00DE; #100;
A = 16'h00EB; B = 16'h00DF; #100;
A = 16'h00EB; B = 16'h00E0; #100;
A = 16'h00EB; B = 16'h00E1; #100;
A = 16'h00EB; B = 16'h00E2; #100;
A = 16'h00EB; B = 16'h00E3; #100;
A = 16'h00EB; B = 16'h00E4; #100;
A = 16'h00EB; B = 16'h00E5; #100;
A = 16'h00EB; B = 16'h00E6; #100;
A = 16'h00EB; B = 16'h00E7; #100;
A = 16'h00EB; B = 16'h00E8; #100;
A = 16'h00EB; B = 16'h00E9; #100;
A = 16'h00EB; B = 16'h00EA; #100;
A = 16'h00EB; B = 16'h00EB; #100;
A = 16'h00EB; B = 16'h00EC; #100;
A = 16'h00EB; B = 16'h00ED; #100;
A = 16'h00EB; B = 16'h00EE; #100;
A = 16'h00EB; B = 16'h00EF; #100;
A = 16'h00EB; B = 16'h00F0; #100;
A = 16'h00EB; B = 16'h00F1; #100;
A = 16'h00EB; B = 16'h00F2; #100;
A = 16'h00EB; B = 16'h00F3; #100;
A = 16'h00EB; B = 16'h00F4; #100;
A = 16'h00EB; B = 16'h00F5; #100;
A = 16'h00EB; B = 16'h00F6; #100;
A = 16'h00EB; B = 16'h00F7; #100;
A = 16'h00EB; B = 16'h00F8; #100;
A = 16'h00EB; B = 16'h00F9; #100;
A = 16'h00EB; B = 16'h00FA; #100;
A = 16'h00EB; B = 16'h00FB; #100;
A = 16'h00EB; B = 16'h00FC; #100;
A = 16'h00EB; B = 16'h00FD; #100;
A = 16'h00EB; B = 16'h00FE; #100;
A = 16'h00EB; B = 16'h00FF; #100;
A = 16'h00EC; B = 16'h000; #100;
A = 16'h00EC; B = 16'h001; #100;
A = 16'h00EC; B = 16'h002; #100;
A = 16'h00EC; B = 16'h003; #100;
A = 16'h00EC; B = 16'h004; #100;
A = 16'h00EC; B = 16'h005; #100;
A = 16'h00EC; B = 16'h006; #100;
A = 16'h00EC; B = 16'h007; #100;
A = 16'h00EC; B = 16'h008; #100;
A = 16'h00EC; B = 16'h009; #100;
A = 16'h00EC; B = 16'h00A; #100;
A = 16'h00EC; B = 16'h00B; #100;
A = 16'h00EC; B = 16'h00C; #100;
A = 16'h00EC; B = 16'h00D; #100;
A = 16'h00EC; B = 16'h00E; #100;
A = 16'h00EC; B = 16'h00F; #100;
A = 16'h00EC; B = 16'h0010; #100;
A = 16'h00EC; B = 16'h0011; #100;
A = 16'h00EC; B = 16'h0012; #100;
A = 16'h00EC; B = 16'h0013; #100;
A = 16'h00EC; B = 16'h0014; #100;
A = 16'h00EC; B = 16'h0015; #100;
A = 16'h00EC; B = 16'h0016; #100;
A = 16'h00EC; B = 16'h0017; #100;
A = 16'h00EC; B = 16'h0018; #100;
A = 16'h00EC; B = 16'h0019; #100;
A = 16'h00EC; B = 16'h001A; #100;
A = 16'h00EC; B = 16'h001B; #100;
A = 16'h00EC; B = 16'h001C; #100;
A = 16'h00EC; B = 16'h001D; #100;
A = 16'h00EC; B = 16'h001E; #100;
A = 16'h00EC; B = 16'h001F; #100;
A = 16'h00EC; B = 16'h0020; #100;
A = 16'h00EC; B = 16'h0021; #100;
A = 16'h00EC; B = 16'h0022; #100;
A = 16'h00EC; B = 16'h0023; #100;
A = 16'h00EC; B = 16'h0024; #100;
A = 16'h00EC; B = 16'h0025; #100;
A = 16'h00EC; B = 16'h0026; #100;
A = 16'h00EC; B = 16'h0027; #100;
A = 16'h00EC; B = 16'h0028; #100;
A = 16'h00EC; B = 16'h0029; #100;
A = 16'h00EC; B = 16'h002A; #100;
A = 16'h00EC; B = 16'h002B; #100;
A = 16'h00EC; B = 16'h002C; #100;
A = 16'h00EC; B = 16'h002D; #100;
A = 16'h00EC; B = 16'h002E; #100;
A = 16'h00EC; B = 16'h002F; #100;
A = 16'h00EC; B = 16'h0030; #100;
A = 16'h00EC; B = 16'h0031; #100;
A = 16'h00EC; B = 16'h0032; #100;
A = 16'h00EC; B = 16'h0033; #100;
A = 16'h00EC; B = 16'h0034; #100;
A = 16'h00EC; B = 16'h0035; #100;
A = 16'h00EC; B = 16'h0036; #100;
A = 16'h00EC; B = 16'h0037; #100;
A = 16'h00EC; B = 16'h0038; #100;
A = 16'h00EC; B = 16'h0039; #100;
A = 16'h00EC; B = 16'h003A; #100;
A = 16'h00EC; B = 16'h003B; #100;
A = 16'h00EC; B = 16'h003C; #100;
A = 16'h00EC; B = 16'h003D; #100;
A = 16'h00EC; B = 16'h003E; #100;
A = 16'h00EC; B = 16'h003F; #100;
A = 16'h00EC; B = 16'h0040; #100;
A = 16'h00EC; B = 16'h0041; #100;
A = 16'h00EC; B = 16'h0042; #100;
A = 16'h00EC; B = 16'h0043; #100;
A = 16'h00EC; B = 16'h0044; #100;
A = 16'h00EC; B = 16'h0045; #100;
A = 16'h00EC; B = 16'h0046; #100;
A = 16'h00EC; B = 16'h0047; #100;
A = 16'h00EC; B = 16'h0048; #100;
A = 16'h00EC; B = 16'h0049; #100;
A = 16'h00EC; B = 16'h004A; #100;
A = 16'h00EC; B = 16'h004B; #100;
A = 16'h00EC; B = 16'h004C; #100;
A = 16'h00EC; B = 16'h004D; #100;
A = 16'h00EC; B = 16'h004E; #100;
A = 16'h00EC; B = 16'h004F; #100;
A = 16'h00EC; B = 16'h0050; #100;
A = 16'h00EC; B = 16'h0051; #100;
A = 16'h00EC; B = 16'h0052; #100;
A = 16'h00EC; B = 16'h0053; #100;
A = 16'h00EC; B = 16'h0054; #100;
A = 16'h00EC; B = 16'h0055; #100;
A = 16'h00EC; B = 16'h0056; #100;
A = 16'h00EC; B = 16'h0057; #100;
A = 16'h00EC; B = 16'h0058; #100;
A = 16'h00EC; B = 16'h0059; #100;
A = 16'h00EC; B = 16'h005A; #100;
A = 16'h00EC; B = 16'h005B; #100;
A = 16'h00EC; B = 16'h005C; #100;
A = 16'h00EC; B = 16'h005D; #100;
A = 16'h00EC; B = 16'h005E; #100;
A = 16'h00EC; B = 16'h005F; #100;
A = 16'h00EC; B = 16'h0060; #100;
A = 16'h00EC; B = 16'h0061; #100;
A = 16'h00EC; B = 16'h0062; #100;
A = 16'h00EC; B = 16'h0063; #100;
A = 16'h00EC; B = 16'h0064; #100;
A = 16'h00EC; B = 16'h0065; #100;
A = 16'h00EC; B = 16'h0066; #100;
A = 16'h00EC; B = 16'h0067; #100;
A = 16'h00EC; B = 16'h0068; #100;
A = 16'h00EC; B = 16'h0069; #100;
A = 16'h00EC; B = 16'h006A; #100;
A = 16'h00EC; B = 16'h006B; #100;
A = 16'h00EC; B = 16'h006C; #100;
A = 16'h00EC; B = 16'h006D; #100;
A = 16'h00EC; B = 16'h006E; #100;
A = 16'h00EC; B = 16'h006F; #100;
A = 16'h00EC; B = 16'h0070; #100;
A = 16'h00EC; B = 16'h0071; #100;
A = 16'h00EC; B = 16'h0072; #100;
A = 16'h00EC; B = 16'h0073; #100;
A = 16'h00EC; B = 16'h0074; #100;
A = 16'h00EC; B = 16'h0075; #100;
A = 16'h00EC; B = 16'h0076; #100;
A = 16'h00EC; B = 16'h0077; #100;
A = 16'h00EC; B = 16'h0078; #100;
A = 16'h00EC; B = 16'h0079; #100;
A = 16'h00EC; B = 16'h007A; #100;
A = 16'h00EC; B = 16'h007B; #100;
A = 16'h00EC; B = 16'h007C; #100;
A = 16'h00EC; B = 16'h007D; #100;
A = 16'h00EC; B = 16'h007E; #100;
A = 16'h00EC; B = 16'h007F; #100;
A = 16'h00EC; B = 16'h0080; #100;
A = 16'h00EC; B = 16'h0081; #100;
A = 16'h00EC; B = 16'h0082; #100;
A = 16'h00EC; B = 16'h0083; #100;
A = 16'h00EC; B = 16'h0084; #100;
A = 16'h00EC; B = 16'h0085; #100;
A = 16'h00EC; B = 16'h0086; #100;
A = 16'h00EC; B = 16'h0087; #100;
A = 16'h00EC; B = 16'h0088; #100;
A = 16'h00EC; B = 16'h0089; #100;
A = 16'h00EC; B = 16'h008A; #100;
A = 16'h00EC; B = 16'h008B; #100;
A = 16'h00EC; B = 16'h008C; #100;
A = 16'h00EC; B = 16'h008D; #100;
A = 16'h00EC; B = 16'h008E; #100;
A = 16'h00EC; B = 16'h008F; #100;
A = 16'h00EC; B = 16'h0090; #100;
A = 16'h00EC; B = 16'h0091; #100;
A = 16'h00EC; B = 16'h0092; #100;
A = 16'h00EC; B = 16'h0093; #100;
A = 16'h00EC; B = 16'h0094; #100;
A = 16'h00EC; B = 16'h0095; #100;
A = 16'h00EC; B = 16'h0096; #100;
A = 16'h00EC; B = 16'h0097; #100;
A = 16'h00EC; B = 16'h0098; #100;
A = 16'h00EC; B = 16'h0099; #100;
A = 16'h00EC; B = 16'h009A; #100;
A = 16'h00EC; B = 16'h009B; #100;
A = 16'h00EC; B = 16'h009C; #100;
A = 16'h00EC; B = 16'h009D; #100;
A = 16'h00EC; B = 16'h009E; #100;
A = 16'h00EC; B = 16'h009F; #100;
A = 16'h00EC; B = 16'h00A0; #100;
A = 16'h00EC; B = 16'h00A1; #100;
A = 16'h00EC; B = 16'h00A2; #100;
A = 16'h00EC; B = 16'h00A3; #100;
A = 16'h00EC; B = 16'h00A4; #100;
A = 16'h00EC; B = 16'h00A5; #100;
A = 16'h00EC; B = 16'h00A6; #100;
A = 16'h00EC; B = 16'h00A7; #100;
A = 16'h00EC; B = 16'h00A8; #100;
A = 16'h00EC; B = 16'h00A9; #100;
A = 16'h00EC; B = 16'h00AA; #100;
A = 16'h00EC; B = 16'h00AB; #100;
A = 16'h00EC; B = 16'h00AC; #100;
A = 16'h00EC; B = 16'h00AD; #100;
A = 16'h00EC; B = 16'h00AE; #100;
A = 16'h00EC; B = 16'h00AF; #100;
A = 16'h00EC; B = 16'h00B0; #100;
A = 16'h00EC; B = 16'h00B1; #100;
A = 16'h00EC; B = 16'h00B2; #100;
A = 16'h00EC; B = 16'h00B3; #100;
A = 16'h00EC; B = 16'h00B4; #100;
A = 16'h00EC; B = 16'h00B5; #100;
A = 16'h00EC; B = 16'h00B6; #100;
A = 16'h00EC; B = 16'h00B7; #100;
A = 16'h00EC; B = 16'h00B8; #100;
A = 16'h00EC; B = 16'h00B9; #100;
A = 16'h00EC; B = 16'h00BA; #100;
A = 16'h00EC; B = 16'h00BB; #100;
A = 16'h00EC; B = 16'h00BC; #100;
A = 16'h00EC; B = 16'h00BD; #100;
A = 16'h00EC; B = 16'h00BE; #100;
A = 16'h00EC; B = 16'h00BF; #100;
A = 16'h00EC; B = 16'h00C0; #100;
A = 16'h00EC; B = 16'h00C1; #100;
A = 16'h00EC; B = 16'h00C2; #100;
A = 16'h00EC; B = 16'h00C3; #100;
A = 16'h00EC; B = 16'h00C4; #100;
A = 16'h00EC; B = 16'h00C5; #100;
A = 16'h00EC; B = 16'h00C6; #100;
A = 16'h00EC; B = 16'h00C7; #100;
A = 16'h00EC; B = 16'h00C8; #100;
A = 16'h00EC; B = 16'h00C9; #100;
A = 16'h00EC; B = 16'h00CA; #100;
A = 16'h00EC; B = 16'h00CB; #100;
A = 16'h00EC; B = 16'h00CC; #100;
A = 16'h00EC; B = 16'h00CD; #100;
A = 16'h00EC; B = 16'h00CE; #100;
A = 16'h00EC; B = 16'h00CF; #100;
A = 16'h00EC; B = 16'h00D0; #100;
A = 16'h00EC; B = 16'h00D1; #100;
A = 16'h00EC; B = 16'h00D2; #100;
A = 16'h00EC; B = 16'h00D3; #100;
A = 16'h00EC; B = 16'h00D4; #100;
A = 16'h00EC; B = 16'h00D5; #100;
A = 16'h00EC; B = 16'h00D6; #100;
A = 16'h00EC; B = 16'h00D7; #100;
A = 16'h00EC; B = 16'h00D8; #100;
A = 16'h00EC; B = 16'h00D9; #100;
A = 16'h00EC; B = 16'h00DA; #100;
A = 16'h00EC; B = 16'h00DB; #100;
A = 16'h00EC; B = 16'h00DC; #100;
A = 16'h00EC; B = 16'h00DD; #100;
A = 16'h00EC; B = 16'h00DE; #100;
A = 16'h00EC; B = 16'h00DF; #100;
A = 16'h00EC; B = 16'h00E0; #100;
A = 16'h00EC; B = 16'h00E1; #100;
A = 16'h00EC; B = 16'h00E2; #100;
A = 16'h00EC; B = 16'h00E3; #100;
A = 16'h00EC; B = 16'h00E4; #100;
A = 16'h00EC; B = 16'h00E5; #100;
A = 16'h00EC; B = 16'h00E6; #100;
A = 16'h00EC; B = 16'h00E7; #100;
A = 16'h00EC; B = 16'h00E8; #100;
A = 16'h00EC; B = 16'h00E9; #100;
A = 16'h00EC; B = 16'h00EA; #100;
A = 16'h00EC; B = 16'h00EB; #100;
A = 16'h00EC; B = 16'h00EC; #100;
A = 16'h00EC; B = 16'h00ED; #100;
A = 16'h00EC; B = 16'h00EE; #100;
A = 16'h00EC; B = 16'h00EF; #100;
A = 16'h00EC; B = 16'h00F0; #100;
A = 16'h00EC; B = 16'h00F1; #100;
A = 16'h00EC; B = 16'h00F2; #100;
A = 16'h00EC; B = 16'h00F3; #100;
A = 16'h00EC; B = 16'h00F4; #100;
A = 16'h00EC; B = 16'h00F5; #100;
A = 16'h00EC; B = 16'h00F6; #100;
A = 16'h00EC; B = 16'h00F7; #100;
A = 16'h00EC; B = 16'h00F8; #100;
A = 16'h00EC; B = 16'h00F9; #100;
A = 16'h00EC; B = 16'h00FA; #100;
A = 16'h00EC; B = 16'h00FB; #100;
A = 16'h00EC; B = 16'h00FC; #100;
A = 16'h00EC; B = 16'h00FD; #100;
A = 16'h00EC; B = 16'h00FE; #100;
A = 16'h00EC; B = 16'h00FF; #100;
A = 16'h00ED; B = 16'h000; #100;
A = 16'h00ED; B = 16'h001; #100;
A = 16'h00ED; B = 16'h002; #100;
A = 16'h00ED; B = 16'h003; #100;
A = 16'h00ED; B = 16'h004; #100;
A = 16'h00ED; B = 16'h005; #100;
A = 16'h00ED; B = 16'h006; #100;
A = 16'h00ED; B = 16'h007; #100;
A = 16'h00ED; B = 16'h008; #100;
A = 16'h00ED; B = 16'h009; #100;
A = 16'h00ED; B = 16'h00A; #100;
A = 16'h00ED; B = 16'h00B; #100;
A = 16'h00ED; B = 16'h00C; #100;
A = 16'h00ED; B = 16'h00D; #100;
A = 16'h00ED; B = 16'h00E; #100;
A = 16'h00ED; B = 16'h00F; #100;
A = 16'h00ED; B = 16'h0010; #100;
A = 16'h00ED; B = 16'h0011; #100;
A = 16'h00ED; B = 16'h0012; #100;
A = 16'h00ED; B = 16'h0013; #100;
A = 16'h00ED; B = 16'h0014; #100;
A = 16'h00ED; B = 16'h0015; #100;
A = 16'h00ED; B = 16'h0016; #100;
A = 16'h00ED; B = 16'h0017; #100;
A = 16'h00ED; B = 16'h0018; #100;
A = 16'h00ED; B = 16'h0019; #100;
A = 16'h00ED; B = 16'h001A; #100;
A = 16'h00ED; B = 16'h001B; #100;
A = 16'h00ED; B = 16'h001C; #100;
A = 16'h00ED; B = 16'h001D; #100;
A = 16'h00ED; B = 16'h001E; #100;
A = 16'h00ED; B = 16'h001F; #100;
A = 16'h00ED; B = 16'h0020; #100;
A = 16'h00ED; B = 16'h0021; #100;
A = 16'h00ED; B = 16'h0022; #100;
A = 16'h00ED; B = 16'h0023; #100;
A = 16'h00ED; B = 16'h0024; #100;
A = 16'h00ED; B = 16'h0025; #100;
A = 16'h00ED; B = 16'h0026; #100;
A = 16'h00ED; B = 16'h0027; #100;
A = 16'h00ED; B = 16'h0028; #100;
A = 16'h00ED; B = 16'h0029; #100;
A = 16'h00ED; B = 16'h002A; #100;
A = 16'h00ED; B = 16'h002B; #100;
A = 16'h00ED; B = 16'h002C; #100;
A = 16'h00ED; B = 16'h002D; #100;
A = 16'h00ED; B = 16'h002E; #100;
A = 16'h00ED; B = 16'h002F; #100;
A = 16'h00ED; B = 16'h0030; #100;
A = 16'h00ED; B = 16'h0031; #100;
A = 16'h00ED; B = 16'h0032; #100;
A = 16'h00ED; B = 16'h0033; #100;
A = 16'h00ED; B = 16'h0034; #100;
A = 16'h00ED; B = 16'h0035; #100;
A = 16'h00ED; B = 16'h0036; #100;
A = 16'h00ED; B = 16'h0037; #100;
A = 16'h00ED; B = 16'h0038; #100;
A = 16'h00ED; B = 16'h0039; #100;
A = 16'h00ED; B = 16'h003A; #100;
A = 16'h00ED; B = 16'h003B; #100;
A = 16'h00ED; B = 16'h003C; #100;
A = 16'h00ED; B = 16'h003D; #100;
A = 16'h00ED; B = 16'h003E; #100;
A = 16'h00ED; B = 16'h003F; #100;
A = 16'h00ED; B = 16'h0040; #100;
A = 16'h00ED; B = 16'h0041; #100;
A = 16'h00ED; B = 16'h0042; #100;
A = 16'h00ED; B = 16'h0043; #100;
A = 16'h00ED; B = 16'h0044; #100;
A = 16'h00ED; B = 16'h0045; #100;
A = 16'h00ED; B = 16'h0046; #100;
A = 16'h00ED; B = 16'h0047; #100;
A = 16'h00ED; B = 16'h0048; #100;
A = 16'h00ED; B = 16'h0049; #100;
A = 16'h00ED; B = 16'h004A; #100;
A = 16'h00ED; B = 16'h004B; #100;
A = 16'h00ED; B = 16'h004C; #100;
A = 16'h00ED; B = 16'h004D; #100;
A = 16'h00ED; B = 16'h004E; #100;
A = 16'h00ED; B = 16'h004F; #100;
A = 16'h00ED; B = 16'h0050; #100;
A = 16'h00ED; B = 16'h0051; #100;
A = 16'h00ED; B = 16'h0052; #100;
A = 16'h00ED; B = 16'h0053; #100;
A = 16'h00ED; B = 16'h0054; #100;
A = 16'h00ED; B = 16'h0055; #100;
A = 16'h00ED; B = 16'h0056; #100;
A = 16'h00ED; B = 16'h0057; #100;
A = 16'h00ED; B = 16'h0058; #100;
A = 16'h00ED; B = 16'h0059; #100;
A = 16'h00ED; B = 16'h005A; #100;
A = 16'h00ED; B = 16'h005B; #100;
A = 16'h00ED; B = 16'h005C; #100;
A = 16'h00ED; B = 16'h005D; #100;
A = 16'h00ED; B = 16'h005E; #100;
A = 16'h00ED; B = 16'h005F; #100;
A = 16'h00ED; B = 16'h0060; #100;
A = 16'h00ED; B = 16'h0061; #100;
A = 16'h00ED; B = 16'h0062; #100;
A = 16'h00ED; B = 16'h0063; #100;
A = 16'h00ED; B = 16'h0064; #100;
A = 16'h00ED; B = 16'h0065; #100;
A = 16'h00ED; B = 16'h0066; #100;
A = 16'h00ED; B = 16'h0067; #100;
A = 16'h00ED; B = 16'h0068; #100;
A = 16'h00ED; B = 16'h0069; #100;
A = 16'h00ED; B = 16'h006A; #100;
A = 16'h00ED; B = 16'h006B; #100;
A = 16'h00ED; B = 16'h006C; #100;
A = 16'h00ED; B = 16'h006D; #100;
A = 16'h00ED; B = 16'h006E; #100;
A = 16'h00ED; B = 16'h006F; #100;
A = 16'h00ED; B = 16'h0070; #100;
A = 16'h00ED; B = 16'h0071; #100;
A = 16'h00ED; B = 16'h0072; #100;
A = 16'h00ED; B = 16'h0073; #100;
A = 16'h00ED; B = 16'h0074; #100;
A = 16'h00ED; B = 16'h0075; #100;
A = 16'h00ED; B = 16'h0076; #100;
A = 16'h00ED; B = 16'h0077; #100;
A = 16'h00ED; B = 16'h0078; #100;
A = 16'h00ED; B = 16'h0079; #100;
A = 16'h00ED; B = 16'h007A; #100;
A = 16'h00ED; B = 16'h007B; #100;
A = 16'h00ED; B = 16'h007C; #100;
A = 16'h00ED; B = 16'h007D; #100;
A = 16'h00ED; B = 16'h007E; #100;
A = 16'h00ED; B = 16'h007F; #100;
A = 16'h00ED; B = 16'h0080; #100;
A = 16'h00ED; B = 16'h0081; #100;
A = 16'h00ED; B = 16'h0082; #100;
A = 16'h00ED; B = 16'h0083; #100;
A = 16'h00ED; B = 16'h0084; #100;
A = 16'h00ED; B = 16'h0085; #100;
A = 16'h00ED; B = 16'h0086; #100;
A = 16'h00ED; B = 16'h0087; #100;
A = 16'h00ED; B = 16'h0088; #100;
A = 16'h00ED; B = 16'h0089; #100;
A = 16'h00ED; B = 16'h008A; #100;
A = 16'h00ED; B = 16'h008B; #100;
A = 16'h00ED; B = 16'h008C; #100;
A = 16'h00ED; B = 16'h008D; #100;
A = 16'h00ED; B = 16'h008E; #100;
A = 16'h00ED; B = 16'h008F; #100;
A = 16'h00ED; B = 16'h0090; #100;
A = 16'h00ED; B = 16'h0091; #100;
A = 16'h00ED; B = 16'h0092; #100;
A = 16'h00ED; B = 16'h0093; #100;
A = 16'h00ED; B = 16'h0094; #100;
A = 16'h00ED; B = 16'h0095; #100;
A = 16'h00ED; B = 16'h0096; #100;
A = 16'h00ED; B = 16'h0097; #100;
A = 16'h00ED; B = 16'h0098; #100;
A = 16'h00ED; B = 16'h0099; #100;
A = 16'h00ED; B = 16'h009A; #100;
A = 16'h00ED; B = 16'h009B; #100;
A = 16'h00ED; B = 16'h009C; #100;
A = 16'h00ED; B = 16'h009D; #100;
A = 16'h00ED; B = 16'h009E; #100;
A = 16'h00ED; B = 16'h009F; #100;
A = 16'h00ED; B = 16'h00A0; #100;
A = 16'h00ED; B = 16'h00A1; #100;
A = 16'h00ED; B = 16'h00A2; #100;
A = 16'h00ED; B = 16'h00A3; #100;
A = 16'h00ED; B = 16'h00A4; #100;
A = 16'h00ED; B = 16'h00A5; #100;
A = 16'h00ED; B = 16'h00A6; #100;
A = 16'h00ED; B = 16'h00A7; #100;
A = 16'h00ED; B = 16'h00A8; #100;
A = 16'h00ED; B = 16'h00A9; #100;
A = 16'h00ED; B = 16'h00AA; #100;
A = 16'h00ED; B = 16'h00AB; #100;
A = 16'h00ED; B = 16'h00AC; #100;
A = 16'h00ED; B = 16'h00AD; #100;
A = 16'h00ED; B = 16'h00AE; #100;
A = 16'h00ED; B = 16'h00AF; #100;
A = 16'h00ED; B = 16'h00B0; #100;
A = 16'h00ED; B = 16'h00B1; #100;
A = 16'h00ED; B = 16'h00B2; #100;
A = 16'h00ED; B = 16'h00B3; #100;
A = 16'h00ED; B = 16'h00B4; #100;
A = 16'h00ED; B = 16'h00B5; #100;
A = 16'h00ED; B = 16'h00B6; #100;
A = 16'h00ED; B = 16'h00B7; #100;
A = 16'h00ED; B = 16'h00B8; #100;
A = 16'h00ED; B = 16'h00B9; #100;
A = 16'h00ED; B = 16'h00BA; #100;
A = 16'h00ED; B = 16'h00BB; #100;
A = 16'h00ED; B = 16'h00BC; #100;
A = 16'h00ED; B = 16'h00BD; #100;
A = 16'h00ED; B = 16'h00BE; #100;
A = 16'h00ED; B = 16'h00BF; #100;
A = 16'h00ED; B = 16'h00C0; #100;
A = 16'h00ED; B = 16'h00C1; #100;
A = 16'h00ED; B = 16'h00C2; #100;
A = 16'h00ED; B = 16'h00C3; #100;
A = 16'h00ED; B = 16'h00C4; #100;
A = 16'h00ED; B = 16'h00C5; #100;
A = 16'h00ED; B = 16'h00C6; #100;
A = 16'h00ED; B = 16'h00C7; #100;
A = 16'h00ED; B = 16'h00C8; #100;
A = 16'h00ED; B = 16'h00C9; #100;
A = 16'h00ED; B = 16'h00CA; #100;
A = 16'h00ED; B = 16'h00CB; #100;
A = 16'h00ED; B = 16'h00CC; #100;
A = 16'h00ED; B = 16'h00CD; #100;
A = 16'h00ED; B = 16'h00CE; #100;
A = 16'h00ED; B = 16'h00CF; #100;
A = 16'h00ED; B = 16'h00D0; #100;
A = 16'h00ED; B = 16'h00D1; #100;
A = 16'h00ED; B = 16'h00D2; #100;
A = 16'h00ED; B = 16'h00D3; #100;
A = 16'h00ED; B = 16'h00D4; #100;
A = 16'h00ED; B = 16'h00D5; #100;
A = 16'h00ED; B = 16'h00D6; #100;
A = 16'h00ED; B = 16'h00D7; #100;
A = 16'h00ED; B = 16'h00D8; #100;
A = 16'h00ED; B = 16'h00D9; #100;
A = 16'h00ED; B = 16'h00DA; #100;
A = 16'h00ED; B = 16'h00DB; #100;
A = 16'h00ED; B = 16'h00DC; #100;
A = 16'h00ED; B = 16'h00DD; #100;
A = 16'h00ED; B = 16'h00DE; #100;
A = 16'h00ED; B = 16'h00DF; #100;
A = 16'h00ED; B = 16'h00E0; #100;
A = 16'h00ED; B = 16'h00E1; #100;
A = 16'h00ED; B = 16'h00E2; #100;
A = 16'h00ED; B = 16'h00E3; #100;
A = 16'h00ED; B = 16'h00E4; #100;
A = 16'h00ED; B = 16'h00E5; #100;
A = 16'h00ED; B = 16'h00E6; #100;
A = 16'h00ED; B = 16'h00E7; #100;
A = 16'h00ED; B = 16'h00E8; #100;
A = 16'h00ED; B = 16'h00E9; #100;
A = 16'h00ED; B = 16'h00EA; #100;
A = 16'h00ED; B = 16'h00EB; #100;
A = 16'h00ED; B = 16'h00EC; #100;
A = 16'h00ED; B = 16'h00ED; #100;
A = 16'h00ED; B = 16'h00EE; #100;
A = 16'h00ED; B = 16'h00EF; #100;
A = 16'h00ED; B = 16'h00F0; #100;
A = 16'h00ED; B = 16'h00F1; #100;
A = 16'h00ED; B = 16'h00F2; #100;
A = 16'h00ED; B = 16'h00F3; #100;
A = 16'h00ED; B = 16'h00F4; #100;
A = 16'h00ED; B = 16'h00F5; #100;
A = 16'h00ED; B = 16'h00F6; #100;
A = 16'h00ED; B = 16'h00F7; #100;
A = 16'h00ED; B = 16'h00F8; #100;
A = 16'h00ED; B = 16'h00F9; #100;
A = 16'h00ED; B = 16'h00FA; #100;
A = 16'h00ED; B = 16'h00FB; #100;
A = 16'h00ED; B = 16'h00FC; #100;
A = 16'h00ED; B = 16'h00FD; #100;
A = 16'h00ED; B = 16'h00FE; #100;
A = 16'h00ED; B = 16'h00FF; #100;
A = 16'h00EE; B = 16'h000; #100;
A = 16'h00EE; B = 16'h001; #100;
A = 16'h00EE; B = 16'h002; #100;
A = 16'h00EE; B = 16'h003; #100;
A = 16'h00EE; B = 16'h004; #100;
A = 16'h00EE; B = 16'h005; #100;
A = 16'h00EE; B = 16'h006; #100;
A = 16'h00EE; B = 16'h007; #100;
A = 16'h00EE; B = 16'h008; #100;
A = 16'h00EE; B = 16'h009; #100;
A = 16'h00EE; B = 16'h00A; #100;
A = 16'h00EE; B = 16'h00B; #100;
A = 16'h00EE; B = 16'h00C; #100;
A = 16'h00EE; B = 16'h00D; #100;
A = 16'h00EE; B = 16'h00E; #100;
A = 16'h00EE; B = 16'h00F; #100;
A = 16'h00EE; B = 16'h0010; #100;
A = 16'h00EE; B = 16'h0011; #100;
A = 16'h00EE; B = 16'h0012; #100;
A = 16'h00EE; B = 16'h0013; #100;
A = 16'h00EE; B = 16'h0014; #100;
A = 16'h00EE; B = 16'h0015; #100;
A = 16'h00EE; B = 16'h0016; #100;
A = 16'h00EE; B = 16'h0017; #100;
A = 16'h00EE; B = 16'h0018; #100;
A = 16'h00EE; B = 16'h0019; #100;
A = 16'h00EE; B = 16'h001A; #100;
A = 16'h00EE; B = 16'h001B; #100;
A = 16'h00EE; B = 16'h001C; #100;
A = 16'h00EE; B = 16'h001D; #100;
A = 16'h00EE; B = 16'h001E; #100;
A = 16'h00EE; B = 16'h001F; #100;
A = 16'h00EE; B = 16'h0020; #100;
A = 16'h00EE; B = 16'h0021; #100;
A = 16'h00EE; B = 16'h0022; #100;
A = 16'h00EE; B = 16'h0023; #100;
A = 16'h00EE; B = 16'h0024; #100;
A = 16'h00EE; B = 16'h0025; #100;
A = 16'h00EE; B = 16'h0026; #100;
A = 16'h00EE; B = 16'h0027; #100;
A = 16'h00EE; B = 16'h0028; #100;
A = 16'h00EE; B = 16'h0029; #100;
A = 16'h00EE; B = 16'h002A; #100;
A = 16'h00EE; B = 16'h002B; #100;
A = 16'h00EE; B = 16'h002C; #100;
A = 16'h00EE; B = 16'h002D; #100;
A = 16'h00EE; B = 16'h002E; #100;
A = 16'h00EE; B = 16'h002F; #100;
A = 16'h00EE; B = 16'h0030; #100;
A = 16'h00EE; B = 16'h0031; #100;
A = 16'h00EE; B = 16'h0032; #100;
A = 16'h00EE; B = 16'h0033; #100;
A = 16'h00EE; B = 16'h0034; #100;
A = 16'h00EE; B = 16'h0035; #100;
A = 16'h00EE; B = 16'h0036; #100;
A = 16'h00EE; B = 16'h0037; #100;
A = 16'h00EE; B = 16'h0038; #100;
A = 16'h00EE; B = 16'h0039; #100;
A = 16'h00EE; B = 16'h003A; #100;
A = 16'h00EE; B = 16'h003B; #100;
A = 16'h00EE; B = 16'h003C; #100;
A = 16'h00EE; B = 16'h003D; #100;
A = 16'h00EE; B = 16'h003E; #100;
A = 16'h00EE; B = 16'h003F; #100;
A = 16'h00EE; B = 16'h0040; #100;
A = 16'h00EE; B = 16'h0041; #100;
A = 16'h00EE; B = 16'h0042; #100;
A = 16'h00EE; B = 16'h0043; #100;
A = 16'h00EE; B = 16'h0044; #100;
A = 16'h00EE; B = 16'h0045; #100;
A = 16'h00EE; B = 16'h0046; #100;
A = 16'h00EE; B = 16'h0047; #100;
A = 16'h00EE; B = 16'h0048; #100;
A = 16'h00EE; B = 16'h0049; #100;
A = 16'h00EE; B = 16'h004A; #100;
A = 16'h00EE; B = 16'h004B; #100;
A = 16'h00EE; B = 16'h004C; #100;
A = 16'h00EE; B = 16'h004D; #100;
A = 16'h00EE; B = 16'h004E; #100;
A = 16'h00EE; B = 16'h004F; #100;
A = 16'h00EE; B = 16'h0050; #100;
A = 16'h00EE; B = 16'h0051; #100;
A = 16'h00EE; B = 16'h0052; #100;
A = 16'h00EE; B = 16'h0053; #100;
A = 16'h00EE; B = 16'h0054; #100;
A = 16'h00EE; B = 16'h0055; #100;
A = 16'h00EE; B = 16'h0056; #100;
A = 16'h00EE; B = 16'h0057; #100;
A = 16'h00EE; B = 16'h0058; #100;
A = 16'h00EE; B = 16'h0059; #100;
A = 16'h00EE; B = 16'h005A; #100;
A = 16'h00EE; B = 16'h005B; #100;
A = 16'h00EE; B = 16'h005C; #100;
A = 16'h00EE; B = 16'h005D; #100;
A = 16'h00EE; B = 16'h005E; #100;
A = 16'h00EE; B = 16'h005F; #100;
A = 16'h00EE; B = 16'h0060; #100;
A = 16'h00EE; B = 16'h0061; #100;
A = 16'h00EE; B = 16'h0062; #100;
A = 16'h00EE; B = 16'h0063; #100;
A = 16'h00EE; B = 16'h0064; #100;
A = 16'h00EE; B = 16'h0065; #100;
A = 16'h00EE; B = 16'h0066; #100;
A = 16'h00EE; B = 16'h0067; #100;
A = 16'h00EE; B = 16'h0068; #100;
A = 16'h00EE; B = 16'h0069; #100;
A = 16'h00EE; B = 16'h006A; #100;
A = 16'h00EE; B = 16'h006B; #100;
A = 16'h00EE; B = 16'h006C; #100;
A = 16'h00EE; B = 16'h006D; #100;
A = 16'h00EE; B = 16'h006E; #100;
A = 16'h00EE; B = 16'h006F; #100;
A = 16'h00EE; B = 16'h0070; #100;
A = 16'h00EE; B = 16'h0071; #100;
A = 16'h00EE; B = 16'h0072; #100;
A = 16'h00EE; B = 16'h0073; #100;
A = 16'h00EE; B = 16'h0074; #100;
A = 16'h00EE; B = 16'h0075; #100;
A = 16'h00EE; B = 16'h0076; #100;
A = 16'h00EE; B = 16'h0077; #100;
A = 16'h00EE; B = 16'h0078; #100;
A = 16'h00EE; B = 16'h0079; #100;
A = 16'h00EE; B = 16'h007A; #100;
A = 16'h00EE; B = 16'h007B; #100;
A = 16'h00EE; B = 16'h007C; #100;
A = 16'h00EE; B = 16'h007D; #100;
A = 16'h00EE; B = 16'h007E; #100;
A = 16'h00EE; B = 16'h007F; #100;
A = 16'h00EE; B = 16'h0080; #100;
A = 16'h00EE; B = 16'h0081; #100;
A = 16'h00EE; B = 16'h0082; #100;
A = 16'h00EE; B = 16'h0083; #100;
A = 16'h00EE; B = 16'h0084; #100;
A = 16'h00EE; B = 16'h0085; #100;
A = 16'h00EE; B = 16'h0086; #100;
A = 16'h00EE; B = 16'h0087; #100;
A = 16'h00EE; B = 16'h0088; #100;
A = 16'h00EE; B = 16'h0089; #100;
A = 16'h00EE; B = 16'h008A; #100;
A = 16'h00EE; B = 16'h008B; #100;
A = 16'h00EE; B = 16'h008C; #100;
A = 16'h00EE; B = 16'h008D; #100;
A = 16'h00EE; B = 16'h008E; #100;
A = 16'h00EE; B = 16'h008F; #100;
A = 16'h00EE; B = 16'h0090; #100;
A = 16'h00EE; B = 16'h0091; #100;
A = 16'h00EE; B = 16'h0092; #100;
A = 16'h00EE; B = 16'h0093; #100;
A = 16'h00EE; B = 16'h0094; #100;
A = 16'h00EE; B = 16'h0095; #100;
A = 16'h00EE; B = 16'h0096; #100;
A = 16'h00EE; B = 16'h0097; #100;
A = 16'h00EE; B = 16'h0098; #100;
A = 16'h00EE; B = 16'h0099; #100;
A = 16'h00EE; B = 16'h009A; #100;
A = 16'h00EE; B = 16'h009B; #100;
A = 16'h00EE; B = 16'h009C; #100;
A = 16'h00EE; B = 16'h009D; #100;
A = 16'h00EE; B = 16'h009E; #100;
A = 16'h00EE; B = 16'h009F; #100;
A = 16'h00EE; B = 16'h00A0; #100;
A = 16'h00EE; B = 16'h00A1; #100;
A = 16'h00EE; B = 16'h00A2; #100;
A = 16'h00EE; B = 16'h00A3; #100;
A = 16'h00EE; B = 16'h00A4; #100;
A = 16'h00EE; B = 16'h00A5; #100;
A = 16'h00EE; B = 16'h00A6; #100;
A = 16'h00EE; B = 16'h00A7; #100;
A = 16'h00EE; B = 16'h00A8; #100;
A = 16'h00EE; B = 16'h00A9; #100;
A = 16'h00EE; B = 16'h00AA; #100;
A = 16'h00EE; B = 16'h00AB; #100;
A = 16'h00EE; B = 16'h00AC; #100;
A = 16'h00EE; B = 16'h00AD; #100;
A = 16'h00EE; B = 16'h00AE; #100;
A = 16'h00EE; B = 16'h00AF; #100;
A = 16'h00EE; B = 16'h00B0; #100;
A = 16'h00EE; B = 16'h00B1; #100;
A = 16'h00EE; B = 16'h00B2; #100;
A = 16'h00EE; B = 16'h00B3; #100;
A = 16'h00EE; B = 16'h00B4; #100;
A = 16'h00EE; B = 16'h00B5; #100;
A = 16'h00EE; B = 16'h00B6; #100;
A = 16'h00EE; B = 16'h00B7; #100;
A = 16'h00EE; B = 16'h00B8; #100;
A = 16'h00EE; B = 16'h00B9; #100;
A = 16'h00EE; B = 16'h00BA; #100;
A = 16'h00EE; B = 16'h00BB; #100;
A = 16'h00EE; B = 16'h00BC; #100;
A = 16'h00EE; B = 16'h00BD; #100;
A = 16'h00EE; B = 16'h00BE; #100;
A = 16'h00EE; B = 16'h00BF; #100;
A = 16'h00EE; B = 16'h00C0; #100;
A = 16'h00EE; B = 16'h00C1; #100;
A = 16'h00EE; B = 16'h00C2; #100;
A = 16'h00EE; B = 16'h00C3; #100;
A = 16'h00EE; B = 16'h00C4; #100;
A = 16'h00EE; B = 16'h00C5; #100;
A = 16'h00EE; B = 16'h00C6; #100;
A = 16'h00EE; B = 16'h00C7; #100;
A = 16'h00EE; B = 16'h00C8; #100;
A = 16'h00EE; B = 16'h00C9; #100;
A = 16'h00EE; B = 16'h00CA; #100;
A = 16'h00EE; B = 16'h00CB; #100;
A = 16'h00EE; B = 16'h00CC; #100;
A = 16'h00EE; B = 16'h00CD; #100;
A = 16'h00EE; B = 16'h00CE; #100;
A = 16'h00EE; B = 16'h00CF; #100;
A = 16'h00EE; B = 16'h00D0; #100;
A = 16'h00EE; B = 16'h00D1; #100;
A = 16'h00EE; B = 16'h00D2; #100;
A = 16'h00EE; B = 16'h00D3; #100;
A = 16'h00EE; B = 16'h00D4; #100;
A = 16'h00EE; B = 16'h00D5; #100;
A = 16'h00EE; B = 16'h00D6; #100;
A = 16'h00EE; B = 16'h00D7; #100;
A = 16'h00EE; B = 16'h00D8; #100;
A = 16'h00EE; B = 16'h00D9; #100;
A = 16'h00EE; B = 16'h00DA; #100;
A = 16'h00EE; B = 16'h00DB; #100;
A = 16'h00EE; B = 16'h00DC; #100;
A = 16'h00EE; B = 16'h00DD; #100;
A = 16'h00EE; B = 16'h00DE; #100;
A = 16'h00EE; B = 16'h00DF; #100;
A = 16'h00EE; B = 16'h00E0; #100;
A = 16'h00EE; B = 16'h00E1; #100;
A = 16'h00EE; B = 16'h00E2; #100;
A = 16'h00EE; B = 16'h00E3; #100;
A = 16'h00EE; B = 16'h00E4; #100;
A = 16'h00EE; B = 16'h00E5; #100;
A = 16'h00EE; B = 16'h00E6; #100;
A = 16'h00EE; B = 16'h00E7; #100;
A = 16'h00EE; B = 16'h00E8; #100;
A = 16'h00EE; B = 16'h00E9; #100;
A = 16'h00EE; B = 16'h00EA; #100;
A = 16'h00EE; B = 16'h00EB; #100;
A = 16'h00EE; B = 16'h00EC; #100;
A = 16'h00EE; B = 16'h00ED; #100;
A = 16'h00EE; B = 16'h00EE; #100;
A = 16'h00EE; B = 16'h00EF; #100;
A = 16'h00EE; B = 16'h00F0; #100;
A = 16'h00EE; B = 16'h00F1; #100;
A = 16'h00EE; B = 16'h00F2; #100;
A = 16'h00EE; B = 16'h00F3; #100;
A = 16'h00EE; B = 16'h00F4; #100;
A = 16'h00EE; B = 16'h00F5; #100;
A = 16'h00EE; B = 16'h00F6; #100;
A = 16'h00EE; B = 16'h00F7; #100;
A = 16'h00EE; B = 16'h00F8; #100;
A = 16'h00EE; B = 16'h00F9; #100;
A = 16'h00EE; B = 16'h00FA; #100;
A = 16'h00EE; B = 16'h00FB; #100;
A = 16'h00EE; B = 16'h00FC; #100;
A = 16'h00EE; B = 16'h00FD; #100;
A = 16'h00EE; B = 16'h00FE; #100;
A = 16'h00EE; B = 16'h00FF; #100;
A = 16'h00EF; B = 16'h000; #100;
A = 16'h00EF; B = 16'h001; #100;
A = 16'h00EF; B = 16'h002; #100;
A = 16'h00EF; B = 16'h003; #100;
A = 16'h00EF; B = 16'h004; #100;
A = 16'h00EF; B = 16'h005; #100;
A = 16'h00EF; B = 16'h006; #100;
A = 16'h00EF; B = 16'h007; #100;
A = 16'h00EF; B = 16'h008; #100;
A = 16'h00EF; B = 16'h009; #100;
A = 16'h00EF; B = 16'h00A; #100;
A = 16'h00EF; B = 16'h00B; #100;
A = 16'h00EF; B = 16'h00C; #100;
A = 16'h00EF; B = 16'h00D; #100;
A = 16'h00EF; B = 16'h00E; #100;
A = 16'h00EF; B = 16'h00F; #100;
A = 16'h00EF; B = 16'h0010; #100;
A = 16'h00EF; B = 16'h0011; #100;
A = 16'h00EF; B = 16'h0012; #100;
A = 16'h00EF; B = 16'h0013; #100;
A = 16'h00EF; B = 16'h0014; #100;
A = 16'h00EF; B = 16'h0015; #100;
A = 16'h00EF; B = 16'h0016; #100;
A = 16'h00EF; B = 16'h0017; #100;
A = 16'h00EF; B = 16'h0018; #100;
A = 16'h00EF; B = 16'h0019; #100;
A = 16'h00EF; B = 16'h001A; #100;
A = 16'h00EF; B = 16'h001B; #100;
A = 16'h00EF; B = 16'h001C; #100;
A = 16'h00EF; B = 16'h001D; #100;
A = 16'h00EF; B = 16'h001E; #100;
A = 16'h00EF; B = 16'h001F; #100;
A = 16'h00EF; B = 16'h0020; #100;
A = 16'h00EF; B = 16'h0021; #100;
A = 16'h00EF; B = 16'h0022; #100;
A = 16'h00EF; B = 16'h0023; #100;
A = 16'h00EF; B = 16'h0024; #100;
A = 16'h00EF; B = 16'h0025; #100;
A = 16'h00EF; B = 16'h0026; #100;
A = 16'h00EF; B = 16'h0027; #100;
A = 16'h00EF; B = 16'h0028; #100;
A = 16'h00EF; B = 16'h0029; #100;
A = 16'h00EF; B = 16'h002A; #100;
A = 16'h00EF; B = 16'h002B; #100;
A = 16'h00EF; B = 16'h002C; #100;
A = 16'h00EF; B = 16'h002D; #100;
A = 16'h00EF; B = 16'h002E; #100;
A = 16'h00EF; B = 16'h002F; #100;
A = 16'h00EF; B = 16'h0030; #100;
A = 16'h00EF; B = 16'h0031; #100;
A = 16'h00EF; B = 16'h0032; #100;
A = 16'h00EF; B = 16'h0033; #100;
A = 16'h00EF; B = 16'h0034; #100;
A = 16'h00EF; B = 16'h0035; #100;
A = 16'h00EF; B = 16'h0036; #100;
A = 16'h00EF; B = 16'h0037; #100;
A = 16'h00EF; B = 16'h0038; #100;
A = 16'h00EF; B = 16'h0039; #100;
A = 16'h00EF; B = 16'h003A; #100;
A = 16'h00EF; B = 16'h003B; #100;
A = 16'h00EF; B = 16'h003C; #100;
A = 16'h00EF; B = 16'h003D; #100;
A = 16'h00EF; B = 16'h003E; #100;
A = 16'h00EF; B = 16'h003F; #100;
A = 16'h00EF; B = 16'h0040; #100;
A = 16'h00EF; B = 16'h0041; #100;
A = 16'h00EF; B = 16'h0042; #100;
A = 16'h00EF; B = 16'h0043; #100;
A = 16'h00EF; B = 16'h0044; #100;
A = 16'h00EF; B = 16'h0045; #100;
A = 16'h00EF; B = 16'h0046; #100;
A = 16'h00EF; B = 16'h0047; #100;
A = 16'h00EF; B = 16'h0048; #100;
A = 16'h00EF; B = 16'h0049; #100;
A = 16'h00EF; B = 16'h004A; #100;
A = 16'h00EF; B = 16'h004B; #100;
A = 16'h00EF; B = 16'h004C; #100;
A = 16'h00EF; B = 16'h004D; #100;
A = 16'h00EF; B = 16'h004E; #100;
A = 16'h00EF; B = 16'h004F; #100;
A = 16'h00EF; B = 16'h0050; #100;
A = 16'h00EF; B = 16'h0051; #100;
A = 16'h00EF; B = 16'h0052; #100;
A = 16'h00EF; B = 16'h0053; #100;
A = 16'h00EF; B = 16'h0054; #100;
A = 16'h00EF; B = 16'h0055; #100;
A = 16'h00EF; B = 16'h0056; #100;
A = 16'h00EF; B = 16'h0057; #100;
A = 16'h00EF; B = 16'h0058; #100;
A = 16'h00EF; B = 16'h0059; #100;
A = 16'h00EF; B = 16'h005A; #100;
A = 16'h00EF; B = 16'h005B; #100;
A = 16'h00EF; B = 16'h005C; #100;
A = 16'h00EF; B = 16'h005D; #100;
A = 16'h00EF; B = 16'h005E; #100;
A = 16'h00EF; B = 16'h005F; #100;
A = 16'h00EF; B = 16'h0060; #100;
A = 16'h00EF; B = 16'h0061; #100;
A = 16'h00EF; B = 16'h0062; #100;
A = 16'h00EF; B = 16'h0063; #100;
A = 16'h00EF; B = 16'h0064; #100;
A = 16'h00EF; B = 16'h0065; #100;
A = 16'h00EF; B = 16'h0066; #100;
A = 16'h00EF; B = 16'h0067; #100;
A = 16'h00EF; B = 16'h0068; #100;
A = 16'h00EF; B = 16'h0069; #100;
A = 16'h00EF; B = 16'h006A; #100;
A = 16'h00EF; B = 16'h006B; #100;
A = 16'h00EF; B = 16'h006C; #100;
A = 16'h00EF; B = 16'h006D; #100;
A = 16'h00EF; B = 16'h006E; #100;
A = 16'h00EF; B = 16'h006F; #100;
A = 16'h00EF; B = 16'h0070; #100;
A = 16'h00EF; B = 16'h0071; #100;
A = 16'h00EF; B = 16'h0072; #100;
A = 16'h00EF; B = 16'h0073; #100;
A = 16'h00EF; B = 16'h0074; #100;
A = 16'h00EF; B = 16'h0075; #100;
A = 16'h00EF; B = 16'h0076; #100;
A = 16'h00EF; B = 16'h0077; #100;
A = 16'h00EF; B = 16'h0078; #100;
A = 16'h00EF; B = 16'h0079; #100;
A = 16'h00EF; B = 16'h007A; #100;
A = 16'h00EF; B = 16'h007B; #100;
A = 16'h00EF; B = 16'h007C; #100;
A = 16'h00EF; B = 16'h007D; #100;
A = 16'h00EF; B = 16'h007E; #100;
A = 16'h00EF; B = 16'h007F; #100;
A = 16'h00EF; B = 16'h0080; #100;
A = 16'h00EF; B = 16'h0081; #100;
A = 16'h00EF; B = 16'h0082; #100;
A = 16'h00EF; B = 16'h0083; #100;
A = 16'h00EF; B = 16'h0084; #100;
A = 16'h00EF; B = 16'h0085; #100;
A = 16'h00EF; B = 16'h0086; #100;
A = 16'h00EF; B = 16'h0087; #100;
A = 16'h00EF; B = 16'h0088; #100;
A = 16'h00EF; B = 16'h0089; #100;
A = 16'h00EF; B = 16'h008A; #100;
A = 16'h00EF; B = 16'h008B; #100;
A = 16'h00EF; B = 16'h008C; #100;
A = 16'h00EF; B = 16'h008D; #100;
A = 16'h00EF; B = 16'h008E; #100;
A = 16'h00EF; B = 16'h008F; #100;
A = 16'h00EF; B = 16'h0090; #100;
A = 16'h00EF; B = 16'h0091; #100;
A = 16'h00EF; B = 16'h0092; #100;
A = 16'h00EF; B = 16'h0093; #100;
A = 16'h00EF; B = 16'h0094; #100;
A = 16'h00EF; B = 16'h0095; #100;
A = 16'h00EF; B = 16'h0096; #100;
A = 16'h00EF; B = 16'h0097; #100;
A = 16'h00EF; B = 16'h0098; #100;
A = 16'h00EF; B = 16'h0099; #100;
A = 16'h00EF; B = 16'h009A; #100;
A = 16'h00EF; B = 16'h009B; #100;
A = 16'h00EF; B = 16'h009C; #100;
A = 16'h00EF; B = 16'h009D; #100;
A = 16'h00EF; B = 16'h009E; #100;
A = 16'h00EF; B = 16'h009F; #100;
A = 16'h00EF; B = 16'h00A0; #100;
A = 16'h00EF; B = 16'h00A1; #100;
A = 16'h00EF; B = 16'h00A2; #100;
A = 16'h00EF; B = 16'h00A3; #100;
A = 16'h00EF; B = 16'h00A4; #100;
A = 16'h00EF; B = 16'h00A5; #100;
A = 16'h00EF; B = 16'h00A6; #100;
A = 16'h00EF; B = 16'h00A7; #100;
A = 16'h00EF; B = 16'h00A8; #100;
A = 16'h00EF; B = 16'h00A9; #100;
A = 16'h00EF; B = 16'h00AA; #100;
A = 16'h00EF; B = 16'h00AB; #100;
A = 16'h00EF; B = 16'h00AC; #100;
A = 16'h00EF; B = 16'h00AD; #100;
A = 16'h00EF; B = 16'h00AE; #100;
A = 16'h00EF; B = 16'h00AF; #100;
A = 16'h00EF; B = 16'h00B0; #100;
A = 16'h00EF; B = 16'h00B1; #100;
A = 16'h00EF; B = 16'h00B2; #100;
A = 16'h00EF; B = 16'h00B3; #100;
A = 16'h00EF; B = 16'h00B4; #100;
A = 16'h00EF; B = 16'h00B5; #100;
A = 16'h00EF; B = 16'h00B6; #100;
A = 16'h00EF; B = 16'h00B7; #100;
A = 16'h00EF; B = 16'h00B8; #100;
A = 16'h00EF; B = 16'h00B9; #100;
A = 16'h00EF; B = 16'h00BA; #100;
A = 16'h00EF; B = 16'h00BB; #100;
A = 16'h00EF; B = 16'h00BC; #100;
A = 16'h00EF; B = 16'h00BD; #100;
A = 16'h00EF; B = 16'h00BE; #100;
A = 16'h00EF; B = 16'h00BF; #100;
A = 16'h00EF; B = 16'h00C0; #100;
A = 16'h00EF; B = 16'h00C1; #100;
A = 16'h00EF; B = 16'h00C2; #100;
A = 16'h00EF; B = 16'h00C3; #100;
A = 16'h00EF; B = 16'h00C4; #100;
A = 16'h00EF; B = 16'h00C5; #100;
A = 16'h00EF; B = 16'h00C6; #100;
A = 16'h00EF; B = 16'h00C7; #100;
A = 16'h00EF; B = 16'h00C8; #100;
A = 16'h00EF; B = 16'h00C9; #100;
A = 16'h00EF; B = 16'h00CA; #100;
A = 16'h00EF; B = 16'h00CB; #100;
A = 16'h00EF; B = 16'h00CC; #100;
A = 16'h00EF; B = 16'h00CD; #100;
A = 16'h00EF; B = 16'h00CE; #100;
A = 16'h00EF; B = 16'h00CF; #100;
A = 16'h00EF; B = 16'h00D0; #100;
A = 16'h00EF; B = 16'h00D1; #100;
A = 16'h00EF; B = 16'h00D2; #100;
A = 16'h00EF; B = 16'h00D3; #100;
A = 16'h00EF; B = 16'h00D4; #100;
A = 16'h00EF; B = 16'h00D5; #100;
A = 16'h00EF; B = 16'h00D6; #100;
A = 16'h00EF; B = 16'h00D7; #100;
A = 16'h00EF; B = 16'h00D8; #100;
A = 16'h00EF; B = 16'h00D9; #100;
A = 16'h00EF; B = 16'h00DA; #100;
A = 16'h00EF; B = 16'h00DB; #100;
A = 16'h00EF; B = 16'h00DC; #100;
A = 16'h00EF; B = 16'h00DD; #100;
A = 16'h00EF; B = 16'h00DE; #100;
A = 16'h00EF; B = 16'h00DF; #100;
A = 16'h00EF; B = 16'h00E0; #100;
A = 16'h00EF; B = 16'h00E1; #100;
A = 16'h00EF; B = 16'h00E2; #100;
A = 16'h00EF; B = 16'h00E3; #100;
A = 16'h00EF; B = 16'h00E4; #100;
A = 16'h00EF; B = 16'h00E5; #100;
A = 16'h00EF; B = 16'h00E6; #100;
A = 16'h00EF; B = 16'h00E7; #100;
A = 16'h00EF; B = 16'h00E8; #100;
A = 16'h00EF; B = 16'h00E9; #100;
A = 16'h00EF; B = 16'h00EA; #100;
A = 16'h00EF; B = 16'h00EB; #100;
A = 16'h00EF; B = 16'h00EC; #100;
A = 16'h00EF; B = 16'h00ED; #100;
A = 16'h00EF; B = 16'h00EE; #100;
A = 16'h00EF; B = 16'h00EF; #100;
A = 16'h00EF; B = 16'h00F0; #100;
A = 16'h00EF; B = 16'h00F1; #100;
A = 16'h00EF; B = 16'h00F2; #100;
A = 16'h00EF; B = 16'h00F3; #100;
A = 16'h00EF; B = 16'h00F4; #100;
A = 16'h00EF; B = 16'h00F5; #100;
A = 16'h00EF; B = 16'h00F6; #100;
A = 16'h00EF; B = 16'h00F7; #100;
A = 16'h00EF; B = 16'h00F8; #100;
A = 16'h00EF; B = 16'h00F9; #100;
A = 16'h00EF; B = 16'h00FA; #100;
A = 16'h00EF; B = 16'h00FB; #100;
A = 16'h00EF; B = 16'h00FC; #100;
A = 16'h00EF; B = 16'h00FD; #100;
A = 16'h00EF; B = 16'h00FE; #100;
A = 16'h00EF; B = 16'h00FF; #100;
A = 16'h00F0; B = 16'h000; #100;
A = 16'h00F0; B = 16'h001; #100;
A = 16'h00F0; B = 16'h002; #100;
A = 16'h00F0; B = 16'h003; #100;
A = 16'h00F0; B = 16'h004; #100;
A = 16'h00F0; B = 16'h005; #100;
A = 16'h00F0; B = 16'h006; #100;
A = 16'h00F0; B = 16'h007; #100;
A = 16'h00F0; B = 16'h008; #100;
A = 16'h00F0; B = 16'h009; #100;
A = 16'h00F0; B = 16'h00A; #100;
A = 16'h00F0; B = 16'h00B; #100;
A = 16'h00F0; B = 16'h00C; #100;
A = 16'h00F0; B = 16'h00D; #100;
A = 16'h00F0; B = 16'h00E; #100;
A = 16'h00F0; B = 16'h00F; #100;
A = 16'h00F0; B = 16'h0010; #100;
A = 16'h00F0; B = 16'h0011; #100;
A = 16'h00F0; B = 16'h0012; #100;
A = 16'h00F0; B = 16'h0013; #100;
A = 16'h00F0; B = 16'h0014; #100;
A = 16'h00F0; B = 16'h0015; #100;
A = 16'h00F0; B = 16'h0016; #100;
A = 16'h00F0; B = 16'h0017; #100;
A = 16'h00F0; B = 16'h0018; #100;
A = 16'h00F0; B = 16'h0019; #100;
A = 16'h00F0; B = 16'h001A; #100;
A = 16'h00F0; B = 16'h001B; #100;
A = 16'h00F0; B = 16'h001C; #100;
A = 16'h00F0; B = 16'h001D; #100;
A = 16'h00F0; B = 16'h001E; #100;
A = 16'h00F0; B = 16'h001F; #100;
A = 16'h00F0; B = 16'h0020; #100;
A = 16'h00F0; B = 16'h0021; #100;
A = 16'h00F0; B = 16'h0022; #100;
A = 16'h00F0; B = 16'h0023; #100;
A = 16'h00F0; B = 16'h0024; #100;
A = 16'h00F0; B = 16'h0025; #100;
A = 16'h00F0; B = 16'h0026; #100;
A = 16'h00F0; B = 16'h0027; #100;
A = 16'h00F0; B = 16'h0028; #100;
A = 16'h00F0; B = 16'h0029; #100;
A = 16'h00F0; B = 16'h002A; #100;
A = 16'h00F0; B = 16'h002B; #100;
A = 16'h00F0; B = 16'h002C; #100;
A = 16'h00F0; B = 16'h002D; #100;
A = 16'h00F0; B = 16'h002E; #100;
A = 16'h00F0; B = 16'h002F; #100;
A = 16'h00F0; B = 16'h0030; #100;
A = 16'h00F0; B = 16'h0031; #100;
A = 16'h00F0; B = 16'h0032; #100;
A = 16'h00F0; B = 16'h0033; #100;
A = 16'h00F0; B = 16'h0034; #100;
A = 16'h00F0; B = 16'h0035; #100;
A = 16'h00F0; B = 16'h0036; #100;
A = 16'h00F0; B = 16'h0037; #100;
A = 16'h00F0; B = 16'h0038; #100;
A = 16'h00F0; B = 16'h0039; #100;
A = 16'h00F0; B = 16'h003A; #100;
A = 16'h00F0; B = 16'h003B; #100;
A = 16'h00F0; B = 16'h003C; #100;
A = 16'h00F0; B = 16'h003D; #100;
A = 16'h00F0; B = 16'h003E; #100;
A = 16'h00F0; B = 16'h003F; #100;
A = 16'h00F0; B = 16'h0040; #100;
A = 16'h00F0; B = 16'h0041; #100;
A = 16'h00F0; B = 16'h0042; #100;
A = 16'h00F0; B = 16'h0043; #100;
A = 16'h00F0; B = 16'h0044; #100;
A = 16'h00F0; B = 16'h0045; #100;
A = 16'h00F0; B = 16'h0046; #100;
A = 16'h00F0; B = 16'h0047; #100;
A = 16'h00F0; B = 16'h0048; #100;
A = 16'h00F0; B = 16'h0049; #100;
A = 16'h00F0; B = 16'h004A; #100;
A = 16'h00F0; B = 16'h004B; #100;
A = 16'h00F0; B = 16'h004C; #100;
A = 16'h00F0; B = 16'h004D; #100;
A = 16'h00F0; B = 16'h004E; #100;
A = 16'h00F0; B = 16'h004F; #100;
A = 16'h00F0; B = 16'h0050; #100;
A = 16'h00F0; B = 16'h0051; #100;
A = 16'h00F0; B = 16'h0052; #100;
A = 16'h00F0; B = 16'h0053; #100;
A = 16'h00F0; B = 16'h0054; #100;
A = 16'h00F0; B = 16'h0055; #100;
A = 16'h00F0; B = 16'h0056; #100;
A = 16'h00F0; B = 16'h0057; #100;
A = 16'h00F0; B = 16'h0058; #100;
A = 16'h00F0; B = 16'h0059; #100;
A = 16'h00F0; B = 16'h005A; #100;
A = 16'h00F0; B = 16'h005B; #100;
A = 16'h00F0; B = 16'h005C; #100;
A = 16'h00F0; B = 16'h005D; #100;
A = 16'h00F0; B = 16'h005E; #100;
A = 16'h00F0; B = 16'h005F; #100;
A = 16'h00F0; B = 16'h0060; #100;
A = 16'h00F0; B = 16'h0061; #100;
A = 16'h00F0; B = 16'h0062; #100;
A = 16'h00F0; B = 16'h0063; #100;
A = 16'h00F0; B = 16'h0064; #100;
A = 16'h00F0; B = 16'h0065; #100;
A = 16'h00F0; B = 16'h0066; #100;
A = 16'h00F0; B = 16'h0067; #100;
A = 16'h00F0; B = 16'h0068; #100;
A = 16'h00F0; B = 16'h0069; #100;
A = 16'h00F0; B = 16'h006A; #100;
A = 16'h00F0; B = 16'h006B; #100;
A = 16'h00F0; B = 16'h006C; #100;
A = 16'h00F0; B = 16'h006D; #100;
A = 16'h00F0; B = 16'h006E; #100;
A = 16'h00F0; B = 16'h006F; #100;
A = 16'h00F0; B = 16'h0070; #100;
A = 16'h00F0; B = 16'h0071; #100;
A = 16'h00F0; B = 16'h0072; #100;
A = 16'h00F0; B = 16'h0073; #100;
A = 16'h00F0; B = 16'h0074; #100;
A = 16'h00F0; B = 16'h0075; #100;
A = 16'h00F0; B = 16'h0076; #100;
A = 16'h00F0; B = 16'h0077; #100;
A = 16'h00F0; B = 16'h0078; #100;
A = 16'h00F0; B = 16'h0079; #100;
A = 16'h00F0; B = 16'h007A; #100;
A = 16'h00F0; B = 16'h007B; #100;
A = 16'h00F0; B = 16'h007C; #100;
A = 16'h00F0; B = 16'h007D; #100;
A = 16'h00F0; B = 16'h007E; #100;
A = 16'h00F0; B = 16'h007F; #100;
A = 16'h00F0; B = 16'h0080; #100;
A = 16'h00F0; B = 16'h0081; #100;
A = 16'h00F0; B = 16'h0082; #100;
A = 16'h00F0; B = 16'h0083; #100;
A = 16'h00F0; B = 16'h0084; #100;
A = 16'h00F0; B = 16'h0085; #100;
A = 16'h00F0; B = 16'h0086; #100;
A = 16'h00F0; B = 16'h0087; #100;
A = 16'h00F0; B = 16'h0088; #100;
A = 16'h00F0; B = 16'h0089; #100;
A = 16'h00F0; B = 16'h008A; #100;
A = 16'h00F0; B = 16'h008B; #100;
A = 16'h00F0; B = 16'h008C; #100;
A = 16'h00F0; B = 16'h008D; #100;
A = 16'h00F0; B = 16'h008E; #100;
A = 16'h00F0; B = 16'h008F; #100;
A = 16'h00F0; B = 16'h0090; #100;
A = 16'h00F0; B = 16'h0091; #100;
A = 16'h00F0; B = 16'h0092; #100;
A = 16'h00F0; B = 16'h0093; #100;
A = 16'h00F0; B = 16'h0094; #100;
A = 16'h00F0; B = 16'h0095; #100;
A = 16'h00F0; B = 16'h0096; #100;
A = 16'h00F0; B = 16'h0097; #100;
A = 16'h00F0; B = 16'h0098; #100;
A = 16'h00F0; B = 16'h0099; #100;
A = 16'h00F0; B = 16'h009A; #100;
A = 16'h00F0; B = 16'h009B; #100;
A = 16'h00F0; B = 16'h009C; #100;
A = 16'h00F0; B = 16'h009D; #100;
A = 16'h00F0; B = 16'h009E; #100;
A = 16'h00F0; B = 16'h009F; #100;
A = 16'h00F0; B = 16'h00A0; #100;
A = 16'h00F0; B = 16'h00A1; #100;
A = 16'h00F0; B = 16'h00A2; #100;
A = 16'h00F0; B = 16'h00A3; #100;
A = 16'h00F0; B = 16'h00A4; #100;
A = 16'h00F0; B = 16'h00A5; #100;
A = 16'h00F0; B = 16'h00A6; #100;
A = 16'h00F0; B = 16'h00A7; #100;
A = 16'h00F0; B = 16'h00A8; #100;
A = 16'h00F0; B = 16'h00A9; #100;
A = 16'h00F0; B = 16'h00AA; #100;
A = 16'h00F0; B = 16'h00AB; #100;
A = 16'h00F0; B = 16'h00AC; #100;
A = 16'h00F0; B = 16'h00AD; #100;
A = 16'h00F0; B = 16'h00AE; #100;
A = 16'h00F0; B = 16'h00AF; #100;
A = 16'h00F0; B = 16'h00B0; #100;
A = 16'h00F0; B = 16'h00B1; #100;
A = 16'h00F0; B = 16'h00B2; #100;
A = 16'h00F0; B = 16'h00B3; #100;
A = 16'h00F0; B = 16'h00B4; #100;
A = 16'h00F0; B = 16'h00B5; #100;
A = 16'h00F0; B = 16'h00B6; #100;
A = 16'h00F0; B = 16'h00B7; #100;
A = 16'h00F0; B = 16'h00B8; #100;
A = 16'h00F0; B = 16'h00B9; #100;
A = 16'h00F0; B = 16'h00BA; #100;
A = 16'h00F0; B = 16'h00BB; #100;
A = 16'h00F0; B = 16'h00BC; #100;
A = 16'h00F0; B = 16'h00BD; #100;
A = 16'h00F0; B = 16'h00BE; #100;
A = 16'h00F0; B = 16'h00BF; #100;
A = 16'h00F0; B = 16'h00C0; #100;
A = 16'h00F0; B = 16'h00C1; #100;
A = 16'h00F0; B = 16'h00C2; #100;
A = 16'h00F0; B = 16'h00C3; #100;
A = 16'h00F0; B = 16'h00C4; #100;
A = 16'h00F0; B = 16'h00C5; #100;
A = 16'h00F0; B = 16'h00C6; #100;
A = 16'h00F0; B = 16'h00C7; #100;
A = 16'h00F0; B = 16'h00C8; #100;
A = 16'h00F0; B = 16'h00C9; #100;
A = 16'h00F0; B = 16'h00CA; #100;
A = 16'h00F0; B = 16'h00CB; #100;
A = 16'h00F0; B = 16'h00CC; #100;
A = 16'h00F0; B = 16'h00CD; #100;
A = 16'h00F0; B = 16'h00CE; #100;
A = 16'h00F0; B = 16'h00CF; #100;
A = 16'h00F0; B = 16'h00D0; #100;
A = 16'h00F0; B = 16'h00D1; #100;
A = 16'h00F0; B = 16'h00D2; #100;
A = 16'h00F0; B = 16'h00D3; #100;
A = 16'h00F0; B = 16'h00D4; #100;
A = 16'h00F0; B = 16'h00D5; #100;
A = 16'h00F0; B = 16'h00D6; #100;
A = 16'h00F0; B = 16'h00D7; #100;
A = 16'h00F0; B = 16'h00D8; #100;
A = 16'h00F0; B = 16'h00D9; #100;
A = 16'h00F0; B = 16'h00DA; #100;
A = 16'h00F0; B = 16'h00DB; #100;
A = 16'h00F0; B = 16'h00DC; #100;
A = 16'h00F0; B = 16'h00DD; #100;
A = 16'h00F0; B = 16'h00DE; #100;
A = 16'h00F0; B = 16'h00DF; #100;
A = 16'h00F0; B = 16'h00E0; #100;
A = 16'h00F0; B = 16'h00E1; #100;
A = 16'h00F0; B = 16'h00E2; #100;
A = 16'h00F0; B = 16'h00E3; #100;
A = 16'h00F0; B = 16'h00E4; #100;
A = 16'h00F0; B = 16'h00E5; #100;
A = 16'h00F0; B = 16'h00E6; #100;
A = 16'h00F0; B = 16'h00E7; #100;
A = 16'h00F0; B = 16'h00E8; #100;
A = 16'h00F0; B = 16'h00E9; #100;
A = 16'h00F0; B = 16'h00EA; #100;
A = 16'h00F0; B = 16'h00EB; #100;
A = 16'h00F0; B = 16'h00EC; #100;
A = 16'h00F0; B = 16'h00ED; #100;
A = 16'h00F0; B = 16'h00EE; #100;
A = 16'h00F0; B = 16'h00EF; #100;
A = 16'h00F0; B = 16'h00F0; #100;
A = 16'h00F0; B = 16'h00F1; #100;
A = 16'h00F0; B = 16'h00F2; #100;
A = 16'h00F0; B = 16'h00F3; #100;
A = 16'h00F0; B = 16'h00F4; #100;
A = 16'h00F0; B = 16'h00F5; #100;
A = 16'h00F0; B = 16'h00F6; #100;
A = 16'h00F0; B = 16'h00F7; #100;
A = 16'h00F0; B = 16'h00F8; #100;
A = 16'h00F0; B = 16'h00F9; #100;
A = 16'h00F0; B = 16'h00FA; #100;
A = 16'h00F0; B = 16'h00FB; #100;
A = 16'h00F0; B = 16'h00FC; #100;
A = 16'h00F0; B = 16'h00FD; #100;
A = 16'h00F0; B = 16'h00FE; #100;
A = 16'h00F0; B = 16'h00FF; #100;
A = 16'h00F1; B = 16'h000; #100;
A = 16'h00F1; B = 16'h001; #100;
A = 16'h00F1; B = 16'h002; #100;
A = 16'h00F1; B = 16'h003; #100;
A = 16'h00F1; B = 16'h004; #100;
A = 16'h00F1; B = 16'h005; #100;
A = 16'h00F1; B = 16'h006; #100;
A = 16'h00F1; B = 16'h007; #100;
A = 16'h00F1; B = 16'h008; #100;
A = 16'h00F1; B = 16'h009; #100;
A = 16'h00F1; B = 16'h00A; #100;
A = 16'h00F1; B = 16'h00B; #100;
A = 16'h00F1; B = 16'h00C; #100;
A = 16'h00F1; B = 16'h00D; #100;
A = 16'h00F1; B = 16'h00E; #100;
A = 16'h00F1; B = 16'h00F; #100;
A = 16'h00F1; B = 16'h0010; #100;
A = 16'h00F1; B = 16'h0011; #100;
A = 16'h00F1; B = 16'h0012; #100;
A = 16'h00F1; B = 16'h0013; #100;
A = 16'h00F1; B = 16'h0014; #100;
A = 16'h00F1; B = 16'h0015; #100;
A = 16'h00F1; B = 16'h0016; #100;
A = 16'h00F1; B = 16'h0017; #100;
A = 16'h00F1; B = 16'h0018; #100;
A = 16'h00F1; B = 16'h0019; #100;
A = 16'h00F1; B = 16'h001A; #100;
A = 16'h00F1; B = 16'h001B; #100;
A = 16'h00F1; B = 16'h001C; #100;
A = 16'h00F1; B = 16'h001D; #100;
A = 16'h00F1; B = 16'h001E; #100;
A = 16'h00F1; B = 16'h001F; #100;
A = 16'h00F1; B = 16'h0020; #100;
A = 16'h00F1; B = 16'h0021; #100;
A = 16'h00F1; B = 16'h0022; #100;
A = 16'h00F1; B = 16'h0023; #100;
A = 16'h00F1; B = 16'h0024; #100;
A = 16'h00F1; B = 16'h0025; #100;
A = 16'h00F1; B = 16'h0026; #100;
A = 16'h00F1; B = 16'h0027; #100;
A = 16'h00F1; B = 16'h0028; #100;
A = 16'h00F1; B = 16'h0029; #100;
A = 16'h00F1; B = 16'h002A; #100;
A = 16'h00F1; B = 16'h002B; #100;
A = 16'h00F1; B = 16'h002C; #100;
A = 16'h00F1; B = 16'h002D; #100;
A = 16'h00F1; B = 16'h002E; #100;
A = 16'h00F1; B = 16'h002F; #100;
A = 16'h00F1; B = 16'h0030; #100;
A = 16'h00F1; B = 16'h0031; #100;
A = 16'h00F1; B = 16'h0032; #100;
A = 16'h00F1; B = 16'h0033; #100;
A = 16'h00F1; B = 16'h0034; #100;
A = 16'h00F1; B = 16'h0035; #100;
A = 16'h00F1; B = 16'h0036; #100;
A = 16'h00F1; B = 16'h0037; #100;
A = 16'h00F1; B = 16'h0038; #100;
A = 16'h00F1; B = 16'h0039; #100;
A = 16'h00F1; B = 16'h003A; #100;
A = 16'h00F1; B = 16'h003B; #100;
A = 16'h00F1; B = 16'h003C; #100;
A = 16'h00F1; B = 16'h003D; #100;
A = 16'h00F1; B = 16'h003E; #100;
A = 16'h00F1; B = 16'h003F; #100;
A = 16'h00F1; B = 16'h0040; #100;
A = 16'h00F1; B = 16'h0041; #100;
A = 16'h00F1; B = 16'h0042; #100;
A = 16'h00F1; B = 16'h0043; #100;
A = 16'h00F1; B = 16'h0044; #100;
A = 16'h00F1; B = 16'h0045; #100;
A = 16'h00F1; B = 16'h0046; #100;
A = 16'h00F1; B = 16'h0047; #100;
A = 16'h00F1; B = 16'h0048; #100;
A = 16'h00F1; B = 16'h0049; #100;
A = 16'h00F1; B = 16'h004A; #100;
A = 16'h00F1; B = 16'h004B; #100;
A = 16'h00F1; B = 16'h004C; #100;
A = 16'h00F1; B = 16'h004D; #100;
A = 16'h00F1; B = 16'h004E; #100;
A = 16'h00F1; B = 16'h004F; #100;
A = 16'h00F1; B = 16'h0050; #100;
A = 16'h00F1; B = 16'h0051; #100;
A = 16'h00F1; B = 16'h0052; #100;
A = 16'h00F1; B = 16'h0053; #100;
A = 16'h00F1; B = 16'h0054; #100;
A = 16'h00F1; B = 16'h0055; #100;
A = 16'h00F1; B = 16'h0056; #100;
A = 16'h00F1; B = 16'h0057; #100;
A = 16'h00F1; B = 16'h0058; #100;
A = 16'h00F1; B = 16'h0059; #100;
A = 16'h00F1; B = 16'h005A; #100;
A = 16'h00F1; B = 16'h005B; #100;
A = 16'h00F1; B = 16'h005C; #100;
A = 16'h00F1; B = 16'h005D; #100;
A = 16'h00F1; B = 16'h005E; #100;
A = 16'h00F1; B = 16'h005F; #100;
A = 16'h00F1; B = 16'h0060; #100;
A = 16'h00F1; B = 16'h0061; #100;
A = 16'h00F1; B = 16'h0062; #100;
A = 16'h00F1; B = 16'h0063; #100;
A = 16'h00F1; B = 16'h0064; #100;
A = 16'h00F1; B = 16'h0065; #100;
A = 16'h00F1; B = 16'h0066; #100;
A = 16'h00F1; B = 16'h0067; #100;
A = 16'h00F1; B = 16'h0068; #100;
A = 16'h00F1; B = 16'h0069; #100;
A = 16'h00F1; B = 16'h006A; #100;
A = 16'h00F1; B = 16'h006B; #100;
A = 16'h00F1; B = 16'h006C; #100;
A = 16'h00F1; B = 16'h006D; #100;
A = 16'h00F1; B = 16'h006E; #100;
A = 16'h00F1; B = 16'h006F; #100;
A = 16'h00F1; B = 16'h0070; #100;
A = 16'h00F1; B = 16'h0071; #100;
A = 16'h00F1; B = 16'h0072; #100;
A = 16'h00F1; B = 16'h0073; #100;
A = 16'h00F1; B = 16'h0074; #100;
A = 16'h00F1; B = 16'h0075; #100;
A = 16'h00F1; B = 16'h0076; #100;
A = 16'h00F1; B = 16'h0077; #100;
A = 16'h00F1; B = 16'h0078; #100;
A = 16'h00F1; B = 16'h0079; #100;
A = 16'h00F1; B = 16'h007A; #100;
A = 16'h00F1; B = 16'h007B; #100;
A = 16'h00F1; B = 16'h007C; #100;
A = 16'h00F1; B = 16'h007D; #100;
A = 16'h00F1; B = 16'h007E; #100;
A = 16'h00F1; B = 16'h007F; #100;
A = 16'h00F1; B = 16'h0080; #100;
A = 16'h00F1; B = 16'h0081; #100;
A = 16'h00F1; B = 16'h0082; #100;
A = 16'h00F1; B = 16'h0083; #100;
A = 16'h00F1; B = 16'h0084; #100;
A = 16'h00F1; B = 16'h0085; #100;
A = 16'h00F1; B = 16'h0086; #100;
A = 16'h00F1; B = 16'h0087; #100;
A = 16'h00F1; B = 16'h0088; #100;
A = 16'h00F1; B = 16'h0089; #100;
A = 16'h00F1; B = 16'h008A; #100;
A = 16'h00F1; B = 16'h008B; #100;
A = 16'h00F1; B = 16'h008C; #100;
A = 16'h00F1; B = 16'h008D; #100;
A = 16'h00F1; B = 16'h008E; #100;
A = 16'h00F1; B = 16'h008F; #100;
A = 16'h00F1; B = 16'h0090; #100;
A = 16'h00F1; B = 16'h0091; #100;
A = 16'h00F1; B = 16'h0092; #100;
A = 16'h00F1; B = 16'h0093; #100;
A = 16'h00F1; B = 16'h0094; #100;
A = 16'h00F1; B = 16'h0095; #100;
A = 16'h00F1; B = 16'h0096; #100;
A = 16'h00F1; B = 16'h0097; #100;
A = 16'h00F1; B = 16'h0098; #100;
A = 16'h00F1; B = 16'h0099; #100;
A = 16'h00F1; B = 16'h009A; #100;
A = 16'h00F1; B = 16'h009B; #100;
A = 16'h00F1; B = 16'h009C; #100;
A = 16'h00F1; B = 16'h009D; #100;
A = 16'h00F1; B = 16'h009E; #100;
A = 16'h00F1; B = 16'h009F; #100;
A = 16'h00F1; B = 16'h00A0; #100;
A = 16'h00F1; B = 16'h00A1; #100;
A = 16'h00F1; B = 16'h00A2; #100;
A = 16'h00F1; B = 16'h00A3; #100;
A = 16'h00F1; B = 16'h00A4; #100;
A = 16'h00F1; B = 16'h00A5; #100;
A = 16'h00F1; B = 16'h00A6; #100;
A = 16'h00F1; B = 16'h00A7; #100;
A = 16'h00F1; B = 16'h00A8; #100;
A = 16'h00F1; B = 16'h00A9; #100;
A = 16'h00F1; B = 16'h00AA; #100;
A = 16'h00F1; B = 16'h00AB; #100;
A = 16'h00F1; B = 16'h00AC; #100;
A = 16'h00F1; B = 16'h00AD; #100;
A = 16'h00F1; B = 16'h00AE; #100;
A = 16'h00F1; B = 16'h00AF; #100;
A = 16'h00F1; B = 16'h00B0; #100;
A = 16'h00F1; B = 16'h00B1; #100;
A = 16'h00F1; B = 16'h00B2; #100;
A = 16'h00F1; B = 16'h00B3; #100;
A = 16'h00F1; B = 16'h00B4; #100;
A = 16'h00F1; B = 16'h00B5; #100;
A = 16'h00F1; B = 16'h00B6; #100;
A = 16'h00F1; B = 16'h00B7; #100;
A = 16'h00F1; B = 16'h00B8; #100;
A = 16'h00F1; B = 16'h00B9; #100;
A = 16'h00F1; B = 16'h00BA; #100;
A = 16'h00F1; B = 16'h00BB; #100;
A = 16'h00F1; B = 16'h00BC; #100;
A = 16'h00F1; B = 16'h00BD; #100;
A = 16'h00F1; B = 16'h00BE; #100;
A = 16'h00F1; B = 16'h00BF; #100;
A = 16'h00F1; B = 16'h00C0; #100;
A = 16'h00F1; B = 16'h00C1; #100;
A = 16'h00F1; B = 16'h00C2; #100;
A = 16'h00F1; B = 16'h00C3; #100;
A = 16'h00F1; B = 16'h00C4; #100;
A = 16'h00F1; B = 16'h00C5; #100;
A = 16'h00F1; B = 16'h00C6; #100;
A = 16'h00F1; B = 16'h00C7; #100;
A = 16'h00F1; B = 16'h00C8; #100;
A = 16'h00F1; B = 16'h00C9; #100;
A = 16'h00F1; B = 16'h00CA; #100;
A = 16'h00F1; B = 16'h00CB; #100;
A = 16'h00F1; B = 16'h00CC; #100;
A = 16'h00F1; B = 16'h00CD; #100;
A = 16'h00F1; B = 16'h00CE; #100;
A = 16'h00F1; B = 16'h00CF; #100;
A = 16'h00F1; B = 16'h00D0; #100;
A = 16'h00F1; B = 16'h00D1; #100;
A = 16'h00F1; B = 16'h00D2; #100;
A = 16'h00F1; B = 16'h00D3; #100;
A = 16'h00F1; B = 16'h00D4; #100;
A = 16'h00F1; B = 16'h00D5; #100;
A = 16'h00F1; B = 16'h00D6; #100;
A = 16'h00F1; B = 16'h00D7; #100;
A = 16'h00F1; B = 16'h00D8; #100;
A = 16'h00F1; B = 16'h00D9; #100;
A = 16'h00F1; B = 16'h00DA; #100;
A = 16'h00F1; B = 16'h00DB; #100;
A = 16'h00F1; B = 16'h00DC; #100;
A = 16'h00F1; B = 16'h00DD; #100;
A = 16'h00F1; B = 16'h00DE; #100;
A = 16'h00F1; B = 16'h00DF; #100;
A = 16'h00F1; B = 16'h00E0; #100;
A = 16'h00F1; B = 16'h00E1; #100;
A = 16'h00F1; B = 16'h00E2; #100;
A = 16'h00F1; B = 16'h00E3; #100;
A = 16'h00F1; B = 16'h00E4; #100;
A = 16'h00F1; B = 16'h00E5; #100;
A = 16'h00F1; B = 16'h00E6; #100;
A = 16'h00F1; B = 16'h00E7; #100;
A = 16'h00F1; B = 16'h00E8; #100;
A = 16'h00F1; B = 16'h00E9; #100;
A = 16'h00F1; B = 16'h00EA; #100;
A = 16'h00F1; B = 16'h00EB; #100;
A = 16'h00F1; B = 16'h00EC; #100;
A = 16'h00F1; B = 16'h00ED; #100;
A = 16'h00F1; B = 16'h00EE; #100;
A = 16'h00F1; B = 16'h00EF; #100;
A = 16'h00F1; B = 16'h00F0; #100;
A = 16'h00F1; B = 16'h00F1; #100;
A = 16'h00F1; B = 16'h00F2; #100;
A = 16'h00F1; B = 16'h00F3; #100;
A = 16'h00F1; B = 16'h00F4; #100;
A = 16'h00F1; B = 16'h00F5; #100;
A = 16'h00F1; B = 16'h00F6; #100;
A = 16'h00F1; B = 16'h00F7; #100;
A = 16'h00F1; B = 16'h00F8; #100;
A = 16'h00F1; B = 16'h00F9; #100;
A = 16'h00F1; B = 16'h00FA; #100;
A = 16'h00F1; B = 16'h00FB; #100;
A = 16'h00F1; B = 16'h00FC; #100;
A = 16'h00F1; B = 16'h00FD; #100;
A = 16'h00F1; B = 16'h00FE; #100;
A = 16'h00F1; B = 16'h00FF; #100;
A = 16'h00F2; B = 16'h000; #100;
A = 16'h00F2; B = 16'h001; #100;
A = 16'h00F2; B = 16'h002; #100;
A = 16'h00F2; B = 16'h003; #100;
A = 16'h00F2; B = 16'h004; #100;
A = 16'h00F2; B = 16'h005; #100;
A = 16'h00F2; B = 16'h006; #100;
A = 16'h00F2; B = 16'h007; #100;
A = 16'h00F2; B = 16'h008; #100;
A = 16'h00F2; B = 16'h009; #100;
A = 16'h00F2; B = 16'h00A; #100;
A = 16'h00F2; B = 16'h00B; #100;
A = 16'h00F2; B = 16'h00C; #100;
A = 16'h00F2; B = 16'h00D; #100;
A = 16'h00F2; B = 16'h00E; #100;
A = 16'h00F2; B = 16'h00F; #100;
A = 16'h00F2; B = 16'h0010; #100;
A = 16'h00F2; B = 16'h0011; #100;
A = 16'h00F2; B = 16'h0012; #100;
A = 16'h00F2; B = 16'h0013; #100;
A = 16'h00F2; B = 16'h0014; #100;
A = 16'h00F2; B = 16'h0015; #100;
A = 16'h00F2; B = 16'h0016; #100;
A = 16'h00F2; B = 16'h0017; #100;
A = 16'h00F2; B = 16'h0018; #100;
A = 16'h00F2; B = 16'h0019; #100;
A = 16'h00F2; B = 16'h001A; #100;
A = 16'h00F2; B = 16'h001B; #100;
A = 16'h00F2; B = 16'h001C; #100;
A = 16'h00F2; B = 16'h001D; #100;
A = 16'h00F2; B = 16'h001E; #100;
A = 16'h00F2; B = 16'h001F; #100;
A = 16'h00F2; B = 16'h0020; #100;
A = 16'h00F2; B = 16'h0021; #100;
A = 16'h00F2; B = 16'h0022; #100;
A = 16'h00F2; B = 16'h0023; #100;
A = 16'h00F2; B = 16'h0024; #100;
A = 16'h00F2; B = 16'h0025; #100;
A = 16'h00F2; B = 16'h0026; #100;
A = 16'h00F2; B = 16'h0027; #100;
A = 16'h00F2; B = 16'h0028; #100;
A = 16'h00F2; B = 16'h0029; #100;
A = 16'h00F2; B = 16'h002A; #100;
A = 16'h00F2; B = 16'h002B; #100;
A = 16'h00F2; B = 16'h002C; #100;
A = 16'h00F2; B = 16'h002D; #100;
A = 16'h00F2; B = 16'h002E; #100;
A = 16'h00F2; B = 16'h002F; #100;
A = 16'h00F2; B = 16'h0030; #100;
A = 16'h00F2; B = 16'h0031; #100;
A = 16'h00F2; B = 16'h0032; #100;
A = 16'h00F2; B = 16'h0033; #100;
A = 16'h00F2; B = 16'h0034; #100;
A = 16'h00F2; B = 16'h0035; #100;
A = 16'h00F2; B = 16'h0036; #100;
A = 16'h00F2; B = 16'h0037; #100;
A = 16'h00F2; B = 16'h0038; #100;
A = 16'h00F2; B = 16'h0039; #100;
A = 16'h00F2; B = 16'h003A; #100;
A = 16'h00F2; B = 16'h003B; #100;
A = 16'h00F2; B = 16'h003C; #100;
A = 16'h00F2; B = 16'h003D; #100;
A = 16'h00F2; B = 16'h003E; #100;
A = 16'h00F2; B = 16'h003F; #100;
A = 16'h00F2; B = 16'h0040; #100;
A = 16'h00F2; B = 16'h0041; #100;
A = 16'h00F2; B = 16'h0042; #100;
A = 16'h00F2; B = 16'h0043; #100;
A = 16'h00F2; B = 16'h0044; #100;
A = 16'h00F2; B = 16'h0045; #100;
A = 16'h00F2; B = 16'h0046; #100;
A = 16'h00F2; B = 16'h0047; #100;
A = 16'h00F2; B = 16'h0048; #100;
A = 16'h00F2; B = 16'h0049; #100;
A = 16'h00F2; B = 16'h004A; #100;
A = 16'h00F2; B = 16'h004B; #100;
A = 16'h00F2; B = 16'h004C; #100;
A = 16'h00F2; B = 16'h004D; #100;
A = 16'h00F2; B = 16'h004E; #100;
A = 16'h00F2; B = 16'h004F; #100;
A = 16'h00F2; B = 16'h0050; #100;
A = 16'h00F2; B = 16'h0051; #100;
A = 16'h00F2; B = 16'h0052; #100;
A = 16'h00F2; B = 16'h0053; #100;
A = 16'h00F2; B = 16'h0054; #100;
A = 16'h00F2; B = 16'h0055; #100;
A = 16'h00F2; B = 16'h0056; #100;
A = 16'h00F2; B = 16'h0057; #100;
A = 16'h00F2; B = 16'h0058; #100;
A = 16'h00F2; B = 16'h0059; #100;
A = 16'h00F2; B = 16'h005A; #100;
A = 16'h00F2; B = 16'h005B; #100;
A = 16'h00F2; B = 16'h005C; #100;
A = 16'h00F2; B = 16'h005D; #100;
A = 16'h00F2; B = 16'h005E; #100;
A = 16'h00F2; B = 16'h005F; #100;
A = 16'h00F2; B = 16'h0060; #100;
A = 16'h00F2; B = 16'h0061; #100;
A = 16'h00F2; B = 16'h0062; #100;
A = 16'h00F2; B = 16'h0063; #100;
A = 16'h00F2; B = 16'h0064; #100;
A = 16'h00F2; B = 16'h0065; #100;
A = 16'h00F2; B = 16'h0066; #100;
A = 16'h00F2; B = 16'h0067; #100;
A = 16'h00F2; B = 16'h0068; #100;
A = 16'h00F2; B = 16'h0069; #100;
A = 16'h00F2; B = 16'h006A; #100;
A = 16'h00F2; B = 16'h006B; #100;
A = 16'h00F2; B = 16'h006C; #100;
A = 16'h00F2; B = 16'h006D; #100;
A = 16'h00F2; B = 16'h006E; #100;
A = 16'h00F2; B = 16'h006F; #100;
A = 16'h00F2; B = 16'h0070; #100;
A = 16'h00F2; B = 16'h0071; #100;
A = 16'h00F2; B = 16'h0072; #100;
A = 16'h00F2; B = 16'h0073; #100;
A = 16'h00F2; B = 16'h0074; #100;
A = 16'h00F2; B = 16'h0075; #100;
A = 16'h00F2; B = 16'h0076; #100;
A = 16'h00F2; B = 16'h0077; #100;
A = 16'h00F2; B = 16'h0078; #100;
A = 16'h00F2; B = 16'h0079; #100;
A = 16'h00F2; B = 16'h007A; #100;
A = 16'h00F2; B = 16'h007B; #100;
A = 16'h00F2; B = 16'h007C; #100;
A = 16'h00F2; B = 16'h007D; #100;
A = 16'h00F2; B = 16'h007E; #100;
A = 16'h00F2; B = 16'h007F; #100;
A = 16'h00F2; B = 16'h0080; #100;
A = 16'h00F2; B = 16'h0081; #100;
A = 16'h00F2; B = 16'h0082; #100;
A = 16'h00F2; B = 16'h0083; #100;
A = 16'h00F2; B = 16'h0084; #100;
A = 16'h00F2; B = 16'h0085; #100;
A = 16'h00F2; B = 16'h0086; #100;
A = 16'h00F2; B = 16'h0087; #100;
A = 16'h00F2; B = 16'h0088; #100;
A = 16'h00F2; B = 16'h0089; #100;
A = 16'h00F2; B = 16'h008A; #100;
A = 16'h00F2; B = 16'h008B; #100;
A = 16'h00F2; B = 16'h008C; #100;
A = 16'h00F2; B = 16'h008D; #100;
A = 16'h00F2; B = 16'h008E; #100;
A = 16'h00F2; B = 16'h008F; #100;
A = 16'h00F2; B = 16'h0090; #100;
A = 16'h00F2; B = 16'h0091; #100;
A = 16'h00F2; B = 16'h0092; #100;
A = 16'h00F2; B = 16'h0093; #100;
A = 16'h00F2; B = 16'h0094; #100;
A = 16'h00F2; B = 16'h0095; #100;
A = 16'h00F2; B = 16'h0096; #100;
A = 16'h00F2; B = 16'h0097; #100;
A = 16'h00F2; B = 16'h0098; #100;
A = 16'h00F2; B = 16'h0099; #100;
A = 16'h00F2; B = 16'h009A; #100;
A = 16'h00F2; B = 16'h009B; #100;
A = 16'h00F2; B = 16'h009C; #100;
A = 16'h00F2; B = 16'h009D; #100;
A = 16'h00F2; B = 16'h009E; #100;
A = 16'h00F2; B = 16'h009F; #100;
A = 16'h00F2; B = 16'h00A0; #100;
A = 16'h00F2; B = 16'h00A1; #100;
A = 16'h00F2; B = 16'h00A2; #100;
A = 16'h00F2; B = 16'h00A3; #100;
A = 16'h00F2; B = 16'h00A4; #100;
A = 16'h00F2; B = 16'h00A5; #100;
A = 16'h00F2; B = 16'h00A6; #100;
A = 16'h00F2; B = 16'h00A7; #100;
A = 16'h00F2; B = 16'h00A8; #100;
A = 16'h00F2; B = 16'h00A9; #100;
A = 16'h00F2; B = 16'h00AA; #100;
A = 16'h00F2; B = 16'h00AB; #100;
A = 16'h00F2; B = 16'h00AC; #100;
A = 16'h00F2; B = 16'h00AD; #100;
A = 16'h00F2; B = 16'h00AE; #100;
A = 16'h00F2; B = 16'h00AF; #100;
A = 16'h00F2; B = 16'h00B0; #100;
A = 16'h00F2; B = 16'h00B1; #100;
A = 16'h00F2; B = 16'h00B2; #100;
A = 16'h00F2; B = 16'h00B3; #100;
A = 16'h00F2; B = 16'h00B4; #100;
A = 16'h00F2; B = 16'h00B5; #100;
A = 16'h00F2; B = 16'h00B6; #100;
A = 16'h00F2; B = 16'h00B7; #100;
A = 16'h00F2; B = 16'h00B8; #100;
A = 16'h00F2; B = 16'h00B9; #100;
A = 16'h00F2; B = 16'h00BA; #100;
A = 16'h00F2; B = 16'h00BB; #100;
A = 16'h00F2; B = 16'h00BC; #100;
A = 16'h00F2; B = 16'h00BD; #100;
A = 16'h00F2; B = 16'h00BE; #100;
A = 16'h00F2; B = 16'h00BF; #100;
A = 16'h00F2; B = 16'h00C0; #100;
A = 16'h00F2; B = 16'h00C1; #100;
A = 16'h00F2; B = 16'h00C2; #100;
A = 16'h00F2; B = 16'h00C3; #100;
A = 16'h00F2; B = 16'h00C4; #100;
A = 16'h00F2; B = 16'h00C5; #100;
A = 16'h00F2; B = 16'h00C6; #100;
A = 16'h00F2; B = 16'h00C7; #100;
A = 16'h00F2; B = 16'h00C8; #100;
A = 16'h00F2; B = 16'h00C9; #100;
A = 16'h00F2; B = 16'h00CA; #100;
A = 16'h00F2; B = 16'h00CB; #100;
A = 16'h00F2; B = 16'h00CC; #100;
A = 16'h00F2; B = 16'h00CD; #100;
A = 16'h00F2; B = 16'h00CE; #100;
A = 16'h00F2; B = 16'h00CF; #100;
A = 16'h00F2; B = 16'h00D0; #100;
A = 16'h00F2; B = 16'h00D1; #100;
A = 16'h00F2; B = 16'h00D2; #100;
A = 16'h00F2; B = 16'h00D3; #100;
A = 16'h00F2; B = 16'h00D4; #100;
A = 16'h00F2; B = 16'h00D5; #100;
A = 16'h00F2; B = 16'h00D6; #100;
A = 16'h00F2; B = 16'h00D7; #100;
A = 16'h00F2; B = 16'h00D8; #100;
A = 16'h00F2; B = 16'h00D9; #100;
A = 16'h00F2; B = 16'h00DA; #100;
A = 16'h00F2; B = 16'h00DB; #100;
A = 16'h00F2; B = 16'h00DC; #100;
A = 16'h00F2; B = 16'h00DD; #100;
A = 16'h00F2; B = 16'h00DE; #100;
A = 16'h00F2; B = 16'h00DF; #100;
A = 16'h00F2; B = 16'h00E0; #100;
A = 16'h00F2; B = 16'h00E1; #100;
A = 16'h00F2; B = 16'h00E2; #100;
A = 16'h00F2; B = 16'h00E3; #100;
A = 16'h00F2; B = 16'h00E4; #100;
A = 16'h00F2; B = 16'h00E5; #100;
A = 16'h00F2; B = 16'h00E6; #100;
A = 16'h00F2; B = 16'h00E7; #100;
A = 16'h00F2; B = 16'h00E8; #100;
A = 16'h00F2; B = 16'h00E9; #100;
A = 16'h00F2; B = 16'h00EA; #100;
A = 16'h00F2; B = 16'h00EB; #100;
A = 16'h00F2; B = 16'h00EC; #100;
A = 16'h00F2; B = 16'h00ED; #100;
A = 16'h00F2; B = 16'h00EE; #100;
A = 16'h00F2; B = 16'h00EF; #100;
A = 16'h00F2; B = 16'h00F0; #100;
A = 16'h00F2; B = 16'h00F1; #100;
A = 16'h00F2; B = 16'h00F2; #100;
A = 16'h00F2; B = 16'h00F3; #100;
A = 16'h00F2; B = 16'h00F4; #100;
A = 16'h00F2; B = 16'h00F5; #100;
A = 16'h00F2; B = 16'h00F6; #100;
A = 16'h00F2; B = 16'h00F7; #100;
A = 16'h00F2; B = 16'h00F8; #100;
A = 16'h00F2; B = 16'h00F9; #100;
A = 16'h00F2; B = 16'h00FA; #100;
A = 16'h00F2; B = 16'h00FB; #100;
A = 16'h00F2; B = 16'h00FC; #100;
A = 16'h00F2; B = 16'h00FD; #100;
A = 16'h00F2; B = 16'h00FE; #100;
A = 16'h00F2; B = 16'h00FF; #100;
A = 16'h00F3; B = 16'h000; #100;
A = 16'h00F3; B = 16'h001; #100;
A = 16'h00F3; B = 16'h002; #100;
A = 16'h00F3; B = 16'h003; #100;
A = 16'h00F3; B = 16'h004; #100;
A = 16'h00F3; B = 16'h005; #100;
A = 16'h00F3; B = 16'h006; #100;
A = 16'h00F3; B = 16'h007; #100;
A = 16'h00F3; B = 16'h008; #100;
A = 16'h00F3; B = 16'h009; #100;
A = 16'h00F3; B = 16'h00A; #100;
A = 16'h00F3; B = 16'h00B; #100;
A = 16'h00F3; B = 16'h00C; #100;
A = 16'h00F3; B = 16'h00D; #100;
A = 16'h00F3; B = 16'h00E; #100;
A = 16'h00F3; B = 16'h00F; #100;
A = 16'h00F3; B = 16'h0010; #100;
A = 16'h00F3; B = 16'h0011; #100;
A = 16'h00F3; B = 16'h0012; #100;
A = 16'h00F3; B = 16'h0013; #100;
A = 16'h00F3; B = 16'h0014; #100;
A = 16'h00F3; B = 16'h0015; #100;
A = 16'h00F3; B = 16'h0016; #100;
A = 16'h00F3; B = 16'h0017; #100;
A = 16'h00F3; B = 16'h0018; #100;
A = 16'h00F3; B = 16'h0019; #100;
A = 16'h00F3; B = 16'h001A; #100;
A = 16'h00F3; B = 16'h001B; #100;
A = 16'h00F3; B = 16'h001C; #100;
A = 16'h00F3; B = 16'h001D; #100;
A = 16'h00F3; B = 16'h001E; #100;
A = 16'h00F3; B = 16'h001F; #100;
A = 16'h00F3; B = 16'h0020; #100;
A = 16'h00F3; B = 16'h0021; #100;
A = 16'h00F3; B = 16'h0022; #100;
A = 16'h00F3; B = 16'h0023; #100;
A = 16'h00F3; B = 16'h0024; #100;
A = 16'h00F3; B = 16'h0025; #100;
A = 16'h00F3; B = 16'h0026; #100;
A = 16'h00F3; B = 16'h0027; #100;
A = 16'h00F3; B = 16'h0028; #100;
A = 16'h00F3; B = 16'h0029; #100;
A = 16'h00F3; B = 16'h002A; #100;
A = 16'h00F3; B = 16'h002B; #100;
A = 16'h00F3; B = 16'h002C; #100;
A = 16'h00F3; B = 16'h002D; #100;
A = 16'h00F3; B = 16'h002E; #100;
A = 16'h00F3; B = 16'h002F; #100;
A = 16'h00F3; B = 16'h0030; #100;
A = 16'h00F3; B = 16'h0031; #100;
A = 16'h00F3; B = 16'h0032; #100;
A = 16'h00F3; B = 16'h0033; #100;
A = 16'h00F3; B = 16'h0034; #100;
A = 16'h00F3; B = 16'h0035; #100;
A = 16'h00F3; B = 16'h0036; #100;
A = 16'h00F3; B = 16'h0037; #100;
A = 16'h00F3; B = 16'h0038; #100;
A = 16'h00F3; B = 16'h0039; #100;
A = 16'h00F3; B = 16'h003A; #100;
A = 16'h00F3; B = 16'h003B; #100;
A = 16'h00F3; B = 16'h003C; #100;
A = 16'h00F3; B = 16'h003D; #100;
A = 16'h00F3; B = 16'h003E; #100;
A = 16'h00F3; B = 16'h003F; #100;
A = 16'h00F3; B = 16'h0040; #100;
A = 16'h00F3; B = 16'h0041; #100;
A = 16'h00F3; B = 16'h0042; #100;
A = 16'h00F3; B = 16'h0043; #100;
A = 16'h00F3; B = 16'h0044; #100;
A = 16'h00F3; B = 16'h0045; #100;
A = 16'h00F3; B = 16'h0046; #100;
A = 16'h00F3; B = 16'h0047; #100;
A = 16'h00F3; B = 16'h0048; #100;
A = 16'h00F3; B = 16'h0049; #100;
A = 16'h00F3; B = 16'h004A; #100;
A = 16'h00F3; B = 16'h004B; #100;
A = 16'h00F3; B = 16'h004C; #100;
A = 16'h00F3; B = 16'h004D; #100;
A = 16'h00F3; B = 16'h004E; #100;
A = 16'h00F3; B = 16'h004F; #100;
A = 16'h00F3; B = 16'h0050; #100;
A = 16'h00F3; B = 16'h0051; #100;
A = 16'h00F3; B = 16'h0052; #100;
A = 16'h00F3; B = 16'h0053; #100;
A = 16'h00F3; B = 16'h0054; #100;
A = 16'h00F3; B = 16'h0055; #100;
A = 16'h00F3; B = 16'h0056; #100;
A = 16'h00F3; B = 16'h0057; #100;
A = 16'h00F3; B = 16'h0058; #100;
A = 16'h00F3; B = 16'h0059; #100;
A = 16'h00F3; B = 16'h005A; #100;
A = 16'h00F3; B = 16'h005B; #100;
A = 16'h00F3; B = 16'h005C; #100;
A = 16'h00F3; B = 16'h005D; #100;
A = 16'h00F3; B = 16'h005E; #100;
A = 16'h00F3; B = 16'h005F; #100;
A = 16'h00F3; B = 16'h0060; #100;
A = 16'h00F3; B = 16'h0061; #100;
A = 16'h00F3; B = 16'h0062; #100;
A = 16'h00F3; B = 16'h0063; #100;
A = 16'h00F3; B = 16'h0064; #100;
A = 16'h00F3; B = 16'h0065; #100;
A = 16'h00F3; B = 16'h0066; #100;
A = 16'h00F3; B = 16'h0067; #100;
A = 16'h00F3; B = 16'h0068; #100;
A = 16'h00F3; B = 16'h0069; #100;
A = 16'h00F3; B = 16'h006A; #100;
A = 16'h00F3; B = 16'h006B; #100;
A = 16'h00F3; B = 16'h006C; #100;
A = 16'h00F3; B = 16'h006D; #100;
A = 16'h00F3; B = 16'h006E; #100;
A = 16'h00F3; B = 16'h006F; #100;
A = 16'h00F3; B = 16'h0070; #100;
A = 16'h00F3; B = 16'h0071; #100;
A = 16'h00F3; B = 16'h0072; #100;
A = 16'h00F3; B = 16'h0073; #100;
A = 16'h00F3; B = 16'h0074; #100;
A = 16'h00F3; B = 16'h0075; #100;
A = 16'h00F3; B = 16'h0076; #100;
A = 16'h00F3; B = 16'h0077; #100;
A = 16'h00F3; B = 16'h0078; #100;
A = 16'h00F3; B = 16'h0079; #100;
A = 16'h00F3; B = 16'h007A; #100;
A = 16'h00F3; B = 16'h007B; #100;
A = 16'h00F3; B = 16'h007C; #100;
A = 16'h00F3; B = 16'h007D; #100;
A = 16'h00F3; B = 16'h007E; #100;
A = 16'h00F3; B = 16'h007F; #100;
A = 16'h00F3; B = 16'h0080; #100;
A = 16'h00F3; B = 16'h0081; #100;
A = 16'h00F3; B = 16'h0082; #100;
A = 16'h00F3; B = 16'h0083; #100;
A = 16'h00F3; B = 16'h0084; #100;
A = 16'h00F3; B = 16'h0085; #100;
A = 16'h00F3; B = 16'h0086; #100;
A = 16'h00F3; B = 16'h0087; #100;
A = 16'h00F3; B = 16'h0088; #100;
A = 16'h00F3; B = 16'h0089; #100;
A = 16'h00F3; B = 16'h008A; #100;
A = 16'h00F3; B = 16'h008B; #100;
A = 16'h00F3; B = 16'h008C; #100;
A = 16'h00F3; B = 16'h008D; #100;
A = 16'h00F3; B = 16'h008E; #100;
A = 16'h00F3; B = 16'h008F; #100;
A = 16'h00F3; B = 16'h0090; #100;
A = 16'h00F3; B = 16'h0091; #100;
A = 16'h00F3; B = 16'h0092; #100;
A = 16'h00F3; B = 16'h0093; #100;
A = 16'h00F3; B = 16'h0094; #100;
A = 16'h00F3; B = 16'h0095; #100;
A = 16'h00F3; B = 16'h0096; #100;
A = 16'h00F3; B = 16'h0097; #100;
A = 16'h00F3; B = 16'h0098; #100;
A = 16'h00F3; B = 16'h0099; #100;
A = 16'h00F3; B = 16'h009A; #100;
A = 16'h00F3; B = 16'h009B; #100;
A = 16'h00F3; B = 16'h009C; #100;
A = 16'h00F3; B = 16'h009D; #100;
A = 16'h00F3; B = 16'h009E; #100;
A = 16'h00F3; B = 16'h009F; #100;
A = 16'h00F3; B = 16'h00A0; #100;
A = 16'h00F3; B = 16'h00A1; #100;
A = 16'h00F3; B = 16'h00A2; #100;
A = 16'h00F3; B = 16'h00A3; #100;
A = 16'h00F3; B = 16'h00A4; #100;
A = 16'h00F3; B = 16'h00A5; #100;
A = 16'h00F3; B = 16'h00A6; #100;
A = 16'h00F3; B = 16'h00A7; #100;
A = 16'h00F3; B = 16'h00A8; #100;
A = 16'h00F3; B = 16'h00A9; #100;
A = 16'h00F3; B = 16'h00AA; #100;
A = 16'h00F3; B = 16'h00AB; #100;
A = 16'h00F3; B = 16'h00AC; #100;
A = 16'h00F3; B = 16'h00AD; #100;
A = 16'h00F3; B = 16'h00AE; #100;
A = 16'h00F3; B = 16'h00AF; #100;
A = 16'h00F3; B = 16'h00B0; #100;
A = 16'h00F3; B = 16'h00B1; #100;
A = 16'h00F3; B = 16'h00B2; #100;
A = 16'h00F3; B = 16'h00B3; #100;
A = 16'h00F3; B = 16'h00B4; #100;
A = 16'h00F3; B = 16'h00B5; #100;
A = 16'h00F3; B = 16'h00B6; #100;
A = 16'h00F3; B = 16'h00B7; #100;
A = 16'h00F3; B = 16'h00B8; #100;
A = 16'h00F3; B = 16'h00B9; #100;
A = 16'h00F3; B = 16'h00BA; #100;
A = 16'h00F3; B = 16'h00BB; #100;
A = 16'h00F3; B = 16'h00BC; #100;
A = 16'h00F3; B = 16'h00BD; #100;
A = 16'h00F3; B = 16'h00BE; #100;
A = 16'h00F3; B = 16'h00BF; #100;
A = 16'h00F3; B = 16'h00C0; #100;
A = 16'h00F3; B = 16'h00C1; #100;
A = 16'h00F3; B = 16'h00C2; #100;
A = 16'h00F3; B = 16'h00C3; #100;
A = 16'h00F3; B = 16'h00C4; #100;
A = 16'h00F3; B = 16'h00C5; #100;
A = 16'h00F3; B = 16'h00C6; #100;
A = 16'h00F3; B = 16'h00C7; #100;
A = 16'h00F3; B = 16'h00C8; #100;
A = 16'h00F3; B = 16'h00C9; #100;
A = 16'h00F3; B = 16'h00CA; #100;
A = 16'h00F3; B = 16'h00CB; #100;
A = 16'h00F3; B = 16'h00CC; #100;
A = 16'h00F3; B = 16'h00CD; #100;
A = 16'h00F3; B = 16'h00CE; #100;
A = 16'h00F3; B = 16'h00CF; #100;
A = 16'h00F3; B = 16'h00D0; #100;
A = 16'h00F3; B = 16'h00D1; #100;
A = 16'h00F3; B = 16'h00D2; #100;
A = 16'h00F3; B = 16'h00D3; #100;
A = 16'h00F3; B = 16'h00D4; #100;
A = 16'h00F3; B = 16'h00D5; #100;
A = 16'h00F3; B = 16'h00D6; #100;
A = 16'h00F3; B = 16'h00D7; #100;
A = 16'h00F3; B = 16'h00D8; #100;
A = 16'h00F3; B = 16'h00D9; #100;
A = 16'h00F3; B = 16'h00DA; #100;
A = 16'h00F3; B = 16'h00DB; #100;
A = 16'h00F3; B = 16'h00DC; #100;
A = 16'h00F3; B = 16'h00DD; #100;
A = 16'h00F3; B = 16'h00DE; #100;
A = 16'h00F3; B = 16'h00DF; #100;
A = 16'h00F3; B = 16'h00E0; #100;
A = 16'h00F3; B = 16'h00E1; #100;
A = 16'h00F3; B = 16'h00E2; #100;
A = 16'h00F3; B = 16'h00E3; #100;
A = 16'h00F3; B = 16'h00E4; #100;
A = 16'h00F3; B = 16'h00E5; #100;
A = 16'h00F3; B = 16'h00E6; #100;
A = 16'h00F3; B = 16'h00E7; #100;
A = 16'h00F3; B = 16'h00E8; #100;
A = 16'h00F3; B = 16'h00E9; #100;
A = 16'h00F3; B = 16'h00EA; #100;
A = 16'h00F3; B = 16'h00EB; #100;
A = 16'h00F3; B = 16'h00EC; #100;
A = 16'h00F3; B = 16'h00ED; #100;
A = 16'h00F3; B = 16'h00EE; #100;
A = 16'h00F3; B = 16'h00EF; #100;
A = 16'h00F3; B = 16'h00F0; #100;
A = 16'h00F3; B = 16'h00F1; #100;
A = 16'h00F3; B = 16'h00F2; #100;
A = 16'h00F3; B = 16'h00F3; #100;
A = 16'h00F3; B = 16'h00F4; #100;
A = 16'h00F3; B = 16'h00F5; #100;
A = 16'h00F3; B = 16'h00F6; #100;
A = 16'h00F3; B = 16'h00F7; #100;
A = 16'h00F3; B = 16'h00F8; #100;
A = 16'h00F3; B = 16'h00F9; #100;
A = 16'h00F3; B = 16'h00FA; #100;
A = 16'h00F3; B = 16'h00FB; #100;
A = 16'h00F3; B = 16'h00FC; #100;
A = 16'h00F3; B = 16'h00FD; #100;
A = 16'h00F3; B = 16'h00FE; #100;
A = 16'h00F3; B = 16'h00FF; #100;
A = 16'h00F4; B = 16'h000; #100;
A = 16'h00F4; B = 16'h001; #100;
A = 16'h00F4; B = 16'h002; #100;
A = 16'h00F4; B = 16'h003; #100;
A = 16'h00F4; B = 16'h004; #100;
A = 16'h00F4; B = 16'h005; #100;
A = 16'h00F4; B = 16'h006; #100;
A = 16'h00F4; B = 16'h007; #100;
A = 16'h00F4; B = 16'h008; #100;
A = 16'h00F4; B = 16'h009; #100;
A = 16'h00F4; B = 16'h00A; #100;
A = 16'h00F4; B = 16'h00B; #100;
A = 16'h00F4; B = 16'h00C; #100;
A = 16'h00F4; B = 16'h00D; #100;
A = 16'h00F4; B = 16'h00E; #100;
A = 16'h00F4; B = 16'h00F; #100;
A = 16'h00F4; B = 16'h0010; #100;
A = 16'h00F4; B = 16'h0011; #100;
A = 16'h00F4; B = 16'h0012; #100;
A = 16'h00F4; B = 16'h0013; #100;
A = 16'h00F4; B = 16'h0014; #100;
A = 16'h00F4; B = 16'h0015; #100;
A = 16'h00F4; B = 16'h0016; #100;
A = 16'h00F4; B = 16'h0017; #100;
A = 16'h00F4; B = 16'h0018; #100;
A = 16'h00F4; B = 16'h0019; #100;
A = 16'h00F4; B = 16'h001A; #100;
A = 16'h00F4; B = 16'h001B; #100;
A = 16'h00F4; B = 16'h001C; #100;
A = 16'h00F4; B = 16'h001D; #100;
A = 16'h00F4; B = 16'h001E; #100;
A = 16'h00F4; B = 16'h001F; #100;
A = 16'h00F4; B = 16'h0020; #100;
A = 16'h00F4; B = 16'h0021; #100;
A = 16'h00F4; B = 16'h0022; #100;
A = 16'h00F4; B = 16'h0023; #100;
A = 16'h00F4; B = 16'h0024; #100;
A = 16'h00F4; B = 16'h0025; #100;
A = 16'h00F4; B = 16'h0026; #100;
A = 16'h00F4; B = 16'h0027; #100;
A = 16'h00F4; B = 16'h0028; #100;
A = 16'h00F4; B = 16'h0029; #100;
A = 16'h00F4; B = 16'h002A; #100;
A = 16'h00F4; B = 16'h002B; #100;
A = 16'h00F4; B = 16'h002C; #100;
A = 16'h00F4; B = 16'h002D; #100;
A = 16'h00F4; B = 16'h002E; #100;
A = 16'h00F4; B = 16'h002F; #100;
A = 16'h00F4; B = 16'h0030; #100;
A = 16'h00F4; B = 16'h0031; #100;
A = 16'h00F4; B = 16'h0032; #100;
A = 16'h00F4; B = 16'h0033; #100;
A = 16'h00F4; B = 16'h0034; #100;
A = 16'h00F4; B = 16'h0035; #100;
A = 16'h00F4; B = 16'h0036; #100;
A = 16'h00F4; B = 16'h0037; #100;
A = 16'h00F4; B = 16'h0038; #100;
A = 16'h00F4; B = 16'h0039; #100;
A = 16'h00F4; B = 16'h003A; #100;
A = 16'h00F4; B = 16'h003B; #100;
A = 16'h00F4; B = 16'h003C; #100;
A = 16'h00F4; B = 16'h003D; #100;
A = 16'h00F4; B = 16'h003E; #100;
A = 16'h00F4; B = 16'h003F; #100;
A = 16'h00F4; B = 16'h0040; #100;
A = 16'h00F4; B = 16'h0041; #100;
A = 16'h00F4; B = 16'h0042; #100;
A = 16'h00F4; B = 16'h0043; #100;
A = 16'h00F4; B = 16'h0044; #100;
A = 16'h00F4; B = 16'h0045; #100;
A = 16'h00F4; B = 16'h0046; #100;
A = 16'h00F4; B = 16'h0047; #100;
A = 16'h00F4; B = 16'h0048; #100;
A = 16'h00F4; B = 16'h0049; #100;
A = 16'h00F4; B = 16'h004A; #100;
A = 16'h00F4; B = 16'h004B; #100;
A = 16'h00F4; B = 16'h004C; #100;
A = 16'h00F4; B = 16'h004D; #100;
A = 16'h00F4; B = 16'h004E; #100;
A = 16'h00F4; B = 16'h004F; #100;
A = 16'h00F4; B = 16'h0050; #100;
A = 16'h00F4; B = 16'h0051; #100;
A = 16'h00F4; B = 16'h0052; #100;
A = 16'h00F4; B = 16'h0053; #100;
A = 16'h00F4; B = 16'h0054; #100;
A = 16'h00F4; B = 16'h0055; #100;
A = 16'h00F4; B = 16'h0056; #100;
A = 16'h00F4; B = 16'h0057; #100;
A = 16'h00F4; B = 16'h0058; #100;
A = 16'h00F4; B = 16'h0059; #100;
A = 16'h00F4; B = 16'h005A; #100;
A = 16'h00F4; B = 16'h005B; #100;
A = 16'h00F4; B = 16'h005C; #100;
A = 16'h00F4; B = 16'h005D; #100;
A = 16'h00F4; B = 16'h005E; #100;
A = 16'h00F4; B = 16'h005F; #100;
A = 16'h00F4; B = 16'h0060; #100;
A = 16'h00F4; B = 16'h0061; #100;
A = 16'h00F4; B = 16'h0062; #100;
A = 16'h00F4; B = 16'h0063; #100;
A = 16'h00F4; B = 16'h0064; #100;
A = 16'h00F4; B = 16'h0065; #100;
A = 16'h00F4; B = 16'h0066; #100;
A = 16'h00F4; B = 16'h0067; #100;
A = 16'h00F4; B = 16'h0068; #100;
A = 16'h00F4; B = 16'h0069; #100;
A = 16'h00F4; B = 16'h006A; #100;
A = 16'h00F4; B = 16'h006B; #100;
A = 16'h00F4; B = 16'h006C; #100;
A = 16'h00F4; B = 16'h006D; #100;
A = 16'h00F4; B = 16'h006E; #100;
A = 16'h00F4; B = 16'h006F; #100;
A = 16'h00F4; B = 16'h0070; #100;
A = 16'h00F4; B = 16'h0071; #100;
A = 16'h00F4; B = 16'h0072; #100;
A = 16'h00F4; B = 16'h0073; #100;
A = 16'h00F4; B = 16'h0074; #100;
A = 16'h00F4; B = 16'h0075; #100;
A = 16'h00F4; B = 16'h0076; #100;
A = 16'h00F4; B = 16'h0077; #100;
A = 16'h00F4; B = 16'h0078; #100;
A = 16'h00F4; B = 16'h0079; #100;
A = 16'h00F4; B = 16'h007A; #100;
A = 16'h00F4; B = 16'h007B; #100;
A = 16'h00F4; B = 16'h007C; #100;
A = 16'h00F4; B = 16'h007D; #100;
A = 16'h00F4; B = 16'h007E; #100;
A = 16'h00F4; B = 16'h007F; #100;
A = 16'h00F4; B = 16'h0080; #100;
A = 16'h00F4; B = 16'h0081; #100;
A = 16'h00F4; B = 16'h0082; #100;
A = 16'h00F4; B = 16'h0083; #100;
A = 16'h00F4; B = 16'h0084; #100;
A = 16'h00F4; B = 16'h0085; #100;
A = 16'h00F4; B = 16'h0086; #100;
A = 16'h00F4; B = 16'h0087; #100;
A = 16'h00F4; B = 16'h0088; #100;
A = 16'h00F4; B = 16'h0089; #100;
A = 16'h00F4; B = 16'h008A; #100;
A = 16'h00F4; B = 16'h008B; #100;
A = 16'h00F4; B = 16'h008C; #100;
A = 16'h00F4; B = 16'h008D; #100;
A = 16'h00F4; B = 16'h008E; #100;
A = 16'h00F4; B = 16'h008F; #100;
A = 16'h00F4; B = 16'h0090; #100;
A = 16'h00F4; B = 16'h0091; #100;
A = 16'h00F4; B = 16'h0092; #100;
A = 16'h00F4; B = 16'h0093; #100;
A = 16'h00F4; B = 16'h0094; #100;
A = 16'h00F4; B = 16'h0095; #100;
A = 16'h00F4; B = 16'h0096; #100;
A = 16'h00F4; B = 16'h0097; #100;
A = 16'h00F4; B = 16'h0098; #100;
A = 16'h00F4; B = 16'h0099; #100;
A = 16'h00F4; B = 16'h009A; #100;
A = 16'h00F4; B = 16'h009B; #100;
A = 16'h00F4; B = 16'h009C; #100;
A = 16'h00F4; B = 16'h009D; #100;
A = 16'h00F4; B = 16'h009E; #100;
A = 16'h00F4; B = 16'h009F; #100;
A = 16'h00F4; B = 16'h00A0; #100;
A = 16'h00F4; B = 16'h00A1; #100;
A = 16'h00F4; B = 16'h00A2; #100;
A = 16'h00F4; B = 16'h00A3; #100;
A = 16'h00F4; B = 16'h00A4; #100;
A = 16'h00F4; B = 16'h00A5; #100;
A = 16'h00F4; B = 16'h00A6; #100;
A = 16'h00F4; B = 16'h00A7; #100;
A = 16'h00F4; B = 16'h00A8; #100;
A = 16'h00F4; B = 16'h00A9; #100;
A = 16'h00F4; B = 16'h00AA; #100;
A = 16'h00F4; B = 16'h00AB; #100;
A = 16'h00F4; B = 16'h00AC; #100;
A = 16'h00F4; B = 16'h00AD; #100;
A = 16'h00F4; B = 16'h00AE; #100;
A = 16'h00F4; B = 16'h00AF; #100;
A = 16'h00F4; B = 16'h00B0; #100;
A = 16'h00F4; B = 16'h00B1; #100;
A = 16'h00F4; B = 16'h00B2; #100;
A = 16'h00F4; B = 16'h00B3; #100;
A = 16'h00F4; B = 16'h00B4; #100;
A = 16'h00F4; B = 16'h00B5; #100;
A = 16'h00F4; B = 16'h00B6; #100;
A = 16'h00F4; B = 16'h00B7; #100;
A = 16'h00F4; B = 16'h00B8; #100;
A = 16'h00F4; B = 16'h00B9; #100;
A = 16'h00F4; B = 16'h00BA; #100;
A = 16'h00F4; B = 16'h00BB; #100;
A = 16'h00F4; B = 16'h00BC; #100;
A = 16'h00F4; B = 16'h00BD; #100;
A = 16'h00F4; B = 16'h00BE; #100;
A = 16'h00F4; B = 16'h00BF; #100;
A = 16'h00F4; B = 16'h00C0; #100;
A = 16'h00F4; B = 16'h00C1; #100;
A = 16'h00F4; B = 16'h00C2; #100;
A = 16'h00F4; B = 16'h00C3; #100;
A = 16'h00F4; B = 16'h00C4; #100;
A = 16'h00F4; B = 16'h00C5; #100;
A = 16'h00F4; B = 16'h00C6; #100;
A = 16'h00F4; B = 16'h00C7; #100;
A = 16'h00F4; B = 16'h00C8; #100;
A = 16'h00F4; B = 16'h00C9; #100;
A = 16'h00F4; B = 16'h00CA; #100;
A = 16'h00F4; B = 16'h00CB; #100;
A = 16'h00F4; B = 16'h00CC; #100;
A = 16'h00F4; B = 16'h00CD; #100;
A = 16'h00F4; B = 16'h00CE; #100;
A = 16'h00F4; B = 16'h00CF; #100;
A = 16'h00F4; B = 16'h00D0; #100;
A = 16'h00F4; B = 16'h00D1; #100;
A = 16'h00F4; B = 16'h00D2; #100;
A = 16'h00F4; B = 16'h00D3; #100;
A = 16'h00F4; B = 16'h00D4; #100;
A = 16'h00F4; B = 16'h00D5; #100;
A = 16'h00F4; B = 16'h00D6; #100;
A = 16'h00F4; B = 16'h00D7; #100;
A = 16'h00F4; B = 16'h00D8; #100;
A = 16'h00F4; B = 16'h00D9; #100;
A = 16'h00F4; B = 16'h00DA; #100;
A = 16'h00F4; B = 16'h00DB; #100;
A = 16'h00F4; B = 16'h00DC; #100;
A = 16'h00F4; B = 16'h00DD; #100;
A = 16'h00F4; B = 16'h00DE; #100;
A = 16'h00F4; B = 16'h00DF; #100;
A = 16'h00F4; B = 16'h00E0; #100;
A = 16'h00F4; B = 16'h00E1; #100;
A = 16'h00F4; B = 16'h00E2; #100;
A = 16'h00F4; B = 16'h00E3; #100;
A = 16'h00F4; B = 16'h00E4; #100;
A = 16'h00F4; B = 16'h00E5; #100;
A = 16'h00F4; B = 16'h00E6; #100;
A = 16'h00F4; B = 16'h00E7; #100;
A = 16'h00F4; B = 16'h00E8; #100;
A = 16'h00F4; B = 16'h00E9; #100;
A = 16'h00F4; B = 16'h00EA; #100;
A = 16'h00F4; B = 16'h00EB; #100;
A = 16'h00F4; B = 16'h00EC; #100;
A = 16'h00F4; B = 16'h00ED; #100;
A = 16'h00F4; B = 16'h00EE; #100;
A = 16'h00F4; B = 16'h00EF; #100;
A = 16'h00F4; B = 16'h00F0; #100;
A = 16'h00F4; B = 16'h00F1; #100;
A = 16'h00F4; B = 16'h00F2; #100;
A = 16'h00F4; B = 16'h00F3; #100;
A = 16'h00F4; B = 16'h00F4; #100;
A = 16'h00F4; B = 16'h00F5; #100;
A = 16'h00F4; B = 16'h00F6; #100;
A = 16'h00F4; B = 16'h00F7; #100;
A = 16'h00F4; B = 16'h00F8; #100;
A = 16'h00F4; B = 16'h00F9; #100;
A = 16'h00F4; B = 16'h00FA; #100;
A = 16'h00F4; B = 16'h00FB; #100;
A = 16'h00F4; B = 16'h00FC; #100;
A = 16'h00F4; B = 16'h00FD; #100;
A = 16'h00F4; B = 16'h00FE; #100;
A = 16'h00F4; B = 16'h00FF; #100;
A = 16'h00F5; B = 16'h000; #100;
A = 16'h00F5; B = 16'h001; #100;
A = 16'h00F5; B = 16'h002; #100;
A = 16'h00F5; B = 16'h003; #100;
A = 16'h00F5; B = 16'h004; #100;
A = 16'h00F5; B = 16'h005; #100;
A = 16'h00F5; B = 16'h006; #100;
A = 16'h00F5; B = 16'h007; #100;
A = 16'h00F5; B = 16'h008; #100;
A = 16'h00F5; B = 16'h009; #100;
A = 16'h00F5; B = 16'h00A; #100;
A = 16'h00F5; B = 16'h00B; #100;
A = 16'h00F5; B = 16'h00C; #100;
A = 16'h00F5; B = 16'h00D; #100;
A = 16'h00F5; B = 16'h00E; #100;
A = 16'h00F5; B = 16'h00F; #100;
A = 16'h00F5; B = 16'h0010; #100;
A = 16'h00F5; B = 16'h0011; #100;
A = 16'h00F5; B = 16'h0012; #100;
A = 16'h00F5; B = 16'h0013; #100;
A = 16'h00F5; B = 16'h0014; #100;
A = 16'h00F5; B = 16'h0015; #100;
A = 16'h00F5; B = 16'h0016; #100;
A = 16'h00F5; B = 16'h0017; #100;
A = 16'h00F5; B = 16'h0018; #100;
A = 16'h00F5; B = 16'h0019; #100;
A = 16'h00F5; B = 16'h001A; #100;
A = 16'h00F5; B = 16'h001B; #100;
A = 16'h00F5; B = 16'h001C; #100;
A = 16'h00F5; B = 16'h001D; #100;
A = 16'h00F5; B = 16'h001E; #100;
A = 16'h00F5; B = 16'h001F; #100;
A = 16'h00F5; B = 16'h0020; #100;
A = 16'h00F5; B = 16'h0021; #100;
A = 16'h00F5; B = 16'h0022; #100;
A = 16'h00F5; B = 16'h0023; #100;
A = 16'h00F5; B = 16'h0024; #100;
A = 16'h00F5; B = 16'h0025; #100;
A = 16'h00F5; B = 16'h0026; #100;
A = 16'h00F5; B = 16'h0027; #100;
A = 16'h00F5; B = 16'h0028; #100;
A = 16'h00F5; B = 16'h0029; #100;
A = 16'h00F5; B = 16'h002A; #100;
A = 16'h00F5; B = 16'h002B; #100;
A = 16'h00F5; B = 16'h002C; #100;
A = 16'h00F5; B = 16'h002D; #100;
A = 16'h00F5; B = 16'h002E; #100;
A = 16'h00F5; B = 16'h002F; #100;
A = 16'h00F5; B = 16'h0030; #100;
A = 16'h00F5; B = 16'h0031; #100;
A = 16'h00F5; B = 16'h0032; #100;
A = 16'h00F5; B = 16'h0033; #100;
A = 16'h00F5; B = 16'h0034; #100;
A = 16'h00F5; B = 16'h0035; #100;
A = 16'h00F5; B = 16'h0036; #100;
A = 16'h00F5; B = 16'h0037; #100;
A = 16'h00F5; B = 16'h0038; #100;
A = 16'h00F5; B = 16'h0039; #100;
A = 16'h00F5; B = 16'h003A; #100;
A = 16'h00F5; B = 16'h003B; #100;
A = 16'h00F5; B = 16'h003C; #100;
A = 16'h00F5; B = 16'h003D; #100;
A = 16'h00F5; B = 16'h003E; #100;
A = 16'h00F5; B = 16'h003F; #100;
A = 16'h00F5; B = 16'h0040; #100;
A = 16'h00F5; B = 16'h0041; #100;
A = 16'h00F5; B = 16'h0042; #100;
A = 16'h00F5; B = 16'h0043; #100;
A = 16'h00F5; B = 16'h0044; #100;
A = 16'h00F5; B = 16'h0045; #100;
A = 16'h00F5; B = 16'h0046; #100;
A = 16'h00F5; B = 16'h0047; #100;
A = 16'h00F5; B = 16'h0048; #100;
A = 16'h00F5; B = 16'h0049; #100;
A = 16'h00F5; B = 16'h004A; #100;
A = 16'h00F5; B = 16'h004B; #100;
A = 16'h00F5; B = 16'h004C; #100;
A = 16'h00F5; B = 16'h004D; #100;
A = 16'h00F5; B = 16'h004E; #100;
A = 16'h00F5; B = 16'h004F; #100;
A = 16'h00F5; B = 16'h0050; #100;
A = 16'h00F5; B = 16'h0051; #100;
A = 16'h00F5; B = 16'h0052; #100;
A = 16'h00F5; B = 16'h0053; #100;
A = 16'h00F5; B = 16'h0054; #100;
A = 16'h00F5; B = 16'h0055; #100;
A = 16'h00F5; B = 16'h0056; #100;
A = 16'h00F5; B = 16'h0057; #100;
A = 16'h00F5; B = 16'h0058; #100;
A = 16'h00F5; B = 16'h0059; #100;
A = 16'h00F5; B = 16'h005A; #100;
A = 16'h00F5; B = 16'h005B; #100;
A = 16'h00F5; B = 16'h005C; #100;
A = 16'h00F5; B = 16'h005D; #100;
A = 16'h00F5; B = 16'h005E; #100;
A = 16'h00F5; B = 16'h005F; #100;
A = 16'h00F5; B = 16'h0060; #100;
A = 16'h00F5; B = 16'h0061; #100;
A = 16'h00F5; B = 16'h0062; #100;
A = 16'h00F5; B = 16'h0063; #100;
A = 16'h00F5; B = 16'h0064; #100;
A = 16'h00F5; B = 16'h0065; #100;
A = 16'h00F5; B = 16'h0066; #100;
A = 16'h00F5; B = 16'h0067; #100;
A = 16'h00F5; B = 16'h0068; #100;
A = 16'h00F5; B = 16'h0069; #100;
A = 16'h00F5; B = 16'h006A; #100;
A = 16'h00F5; B = 16'h006B; #100;
A = 16'h00F5; B = 16'h006C; #100;
A = 16'h00F5; B = 16'h006D; #100;
A = 16'h00F5; B = 16'h006E; #100;
A = 16'h00F5; B = 16'h006F; #100;
A = 16'h00F5; B = 16'h0070; #100;
A = 16'h00F5; B = 16'h0071; #100;
A = 16'h00F5; B = 16'h0072; #100;
A = 16'h00F5; B = 16'h0073; #100;
A = 16'h00F5; B = 16'h0074; #100;
A = 16'h00F5; B = 16'h0075; #100;
A = 16'h00F5; B = 16'h0076; #100;
A = 16'h00F5; B = 16'h0077; #100;
A = 16'h00F5; B = 16'h0078; #100;
A = 16'h00F5; B = 16'h0079; #100;
A = 16'h00F5; B = 16'h007A; #100;
A = 16'h00F5; B = 16'h007B; #100;
A = 16'h00F5; B = 16'h007C; #100;
A = 16'h00F5; B = 16'h007D; #100;
A = 16'h00F5; B = 16'h007E; #100;
A = 16'h00F5; B = 16'h007F; #100;
A = 16'h00F5; B = 16'h0080; #100;
A = 16'h00F5; B = 16'h0081; #100;
A = 16'h00F5; B = 16'h0082; #100;
A = 16'h00F5; B = 16'h0083; #100;
A = 16'h00F5; B = 16'h0084; #100;
A = 16'h00F5; B = 16'h0085; #100;
A = 16'h00F5; B = 16'h0086; #100;
A = 16'h00F5; B = 16'h0087; #100;
A = 16'h00F5; B = 16'h0088; #100;
A = 16'h00F5; B = 16'h0089; #100;
A = 16'h00F5; B = 16'h008A; #100;
A = 16'h00F5; B = 16'h008B; #100;
A = 16'h00F5; B = 16'h008C; #100;
A = 16'h00F5; B = 16'h008D; #100;
A = 16'h00F5; B = 16'h008E; #100;
A = 16'h00F5; B = 16'h008F; #100;
A = 16'h00F5; B = 16'h0090; #100;
A = 16'h00F5; B = 16'h0091; #100;
A = 16'h00F5; B = 16'h0092; #100;
A = 16'h00F5; B = 16'h0093; #100;
A = 16'h00F5; B = 16'h0094; #100;
A = 16'h00F5; B = 16'h0095; #100;
A = 16'h00F5; B = 16'h0096; #100;
A = 16'h00F5; B = 16'h0097; #100;
A = 16'h00F5; B = 16'h0098; #100;
A = 16'h00F5; B = 16'h0099; #100;
A = 16'h00F5; B = 16'h009A; #100;
A = 16'h00F5; B = 16'h009B; #100;
A = 16'h00F5; B = 16'h009C; #100;
A = 16'h00F5; B = 16'h009D; #100;
A = 16'h00F5; B = 16'h009E; #100;
A = 16'h00F5; B = 16'h009F; #100;
A = 16'h00F5; B = 16'h00A0; #100;
A = 16'h00F5; B = 16'h00A1; #100;
A = 16'h00F5; B = 16'h00A2; #100;
A = 16'h00F5; B = 16'h00A3; #100;
A = 16'h00F5; B = 16'h00A4; #100;
A = 16'h00F5; B = 16'h00A5; #100;
A = 16'h00F5; B = 16'h00A6; #100;
A = 16'h00F5; B = 16'h00A7; #100;
A = 16'h00F5; B = 16'h00A8; #100;
A = 16'h00F5; B = 16'h00A9; #100;
A = 16'h00F5; B = 16'h00AA; #100;
A = 16'h00F5; B = 16'h00AB; #100;
A = 16'h00F5; B = 16'h00AC; #100;
A = 16'h00F5; B = 16'h00AD; #100;
A = 16'h00F5; B = 16'h00AE; #100;
A = 16'h00F5; B = 16'h00AF; #100;
A = 16'h00F5; B = 16'h00B0; #100;
A = 16'h00F5; B = 16'h00B1; #100;
A = 16'h00F5; B = 16'h00B2; #100;
A = 16'h00F5; B = 16'h00B3; #100;
A = 16'h00F5; B = 16'h00B4; #100;
A = 16'h00F5; B = 16'h00B5; #100;
A = 16'h00F5; B = 16'h00B6; #100;
A = 16'h00F5; B = 16'h00B7; #100;
A = 16'h00F5; B = 16'h00B8; #100;
A = 16'h00F5; B = 16'h00B9; #100;
A = 16'h00F5; B = 16'h00BA; #100;
A = 16'h00F5; B = 16'h00BB; #100;
A = 16'h00F5; B = 16'h00BC; #100;
A = 16'h00F5; B = 16'h00BD; #100;
A = 16'h00F5; B = 16'h00BE; #100;
A = 16'h00F5; B = 16'h00BF; #100;
A = 16'h00F5; B = 16'h00C0; #100;
A = 16'h00F5; B = 16'h00C1; #100;
A = 16'h00F5; B = 16'h00C2; #100;
A = 16'h00F5; B = 16'h00C3; #100;
A = 16'h00F5; B = 16'h00C4; #100;
A = 16'h00F5; B = 16'h00C5; #100;
A = 16'h00F5; B = 16'h00C6; #100;
A = 16'h00F5; B = 16'h00C7; #100;
A = 16'h00F5; B = 16'h00C8; #100;
A = 16'h00F5; B = 16'h00C9; #100;
A = 16'h00F5; B = 16'h00CA; #100;
A = 16'h00F5; B = 16'h00CB; #100;
A = 16'h00F5; B = 16'h00CC; #100;
A = 16'h00F5; B = 16'h00CD; #100;
A = 16'h00F5; B = 16'h00CE; #100;
A = 16'h00F5; B = 16'h00CF; #100;
A = 16'h00F5; B = 16'h00D0; #100;
A = 16'h00F5; B = 16'h00D1; #100;
A = 16'h00F5; B = 16'h00D2; #100;
A = 16'h00F5; B = 16'h00D3; #100;
A = 16'h00F5; B = 16'h00D4; #100;
A = 16'h00F5; B = 16'h00D5; #100;
A = 16'h00F5; B = 16'h00D6; #100;
A = 16'h00F5; B = 16'h00D7; #100;
A = 16'h00F5; B = 16'h00D8; #100;
A = 16'h00F5; B = 16'h00D9; #100;
A = 16'h00F5; B = 16'h00DA; #100;
A = 16'h00F5; B = 16'h00DB; #100;
A = 16'h00F5; B = 16'h00DC; #100;
A = 16'h00F5; B = 16'h00DD; #100;
A = 16'h00F5; B = 16'h00DE; #100;
A = 16'h00F5; B = 16'h00DF; #100;
A = 16'h00F5; B = 16'h00E0; #100;
A = 16'h00F5; B = 16'h00E1; #100;
A = 16'h00F5; B = 16'h00E2; #100;
A = 16'h00F5; B = 16'h00E3; #100;
A = 16'h00F5; B = 16'h00E4; #100;
A = 16'h00F5; B = 16'h00E5; #100;
A = 16'h00F5; B = 16'h00E6; #100;
A = 16'h00F5; B = 16'h00E7; #100;
A = 16'h00F5; B = 16'h00E8; #100;
A = 16'h00F5; B = 16'h00E9; #100;
A = 16'h00F5; B = 16'h00EA; #100;
A = 16'h00F5; B = 16'h00EB; #100;
A = 16'h00F5; B = 16'h00EC; #100;
A = 16'h00F5; B = 16'h00ED; #100;
A = 16'h00F5; B = 16'h00EE; #100;
A = 16'h00F5; B = 16'h00EF; #100;
A = 16'h00F5; B = 16'h00F0; #100;
A = 16'h00F5; B = 16'h00F1; #100;
A = 16'h00F5; B = 16'h00F2; #100;
A = 16'h00F5; B = 16'h00F3; #100;
A = 16'h00F5; B = 16'h00F4; #100;
A = 16'h00F5; B = 16'h00F5; #100;
A = 16'h00F5; B = 16'h00F6; #100;
A = 16'h00F5; B = 16'h00F7; #100;
A = 16'h00F5; B = 16'h00F8; #100;
A = 16'h00F5; B = 16'h00F9; #100;
A = 16'h00F5; B = 16'h00FA; #100;
A = 16'h00F5; B = 16'h00FB; #100;
A = 16'h00F5; B = 16'h00FC; #100;
A = 16'h00F5; B = 16'h00FD; #100;
A = 16'h00F5; B = 16'h00FE; #100;
A = 16'h00F5; B = 16'h00FF; #100;
A = 16'h00F6; B = 16'h000; #100;
A = 16'h00F6; B = 16'h001; #100;
A = 16'h00F6; B = 16'h002; #100;
A = 16'h00F6; B = 16'h003; #100;
A = 16'h00F6; B = 16'h004; #100;
A = 16'h00F6; B = 16'h005; #100;
A = 16'h00F6; B = 16'h006; #100;
A = 16'h00F6; B = 16'h007; #100;
A = 16'h00F6; B = 16'h008; #100;
A = 16'h00F6; B = 16'h009; #100;
A = 16'h00F6; B = 16'h00A; #100;
A = 16'h00F6; B = 16'h00B; #100;
A = 16'h00F6; B = 16'h00C; #100;
A = 16'h00F6; B = 16'h00D; #100;
A = 16'h00F6; B = 16'h00E; #100;
A = 16'h00F6; B = 16'h00F; #100;
A = 16'h00F6; B = 16'h0010; #100;
A = 16'h00F6; B = 16'h0011; #100;
A = 16'h00F6; B = 16'h0012; #100;
A = 16'h00F6; B = 16'h0013; #100;
A = 16'h00F6; B = 16'h0014; #100;
A = 16'h00F6; B = 16'h0015; #100;
A = 16'h00F6; B = 16'h0016; #100;
A = 16'h00F6; B = 16'h0017; #100;
A = 16'h00F6; B = 16'h0018; #100;
A = 16'h00F6; B = 16'h0019; #100;
A = 16'h00F6; B = 16'h001A; #100;
A = 16'h00F6; B = 16'h001B; #100;
A = 16'h00F6; B = 16'h001C; #100;
A = 16'h00F6; B = 16'h001D; #100;
A = 16'h00F6; B = 16'h001E; #100;
A = 16'h00F6; B = 16'h001F; #100;
A = 16'h00F6; B = 16'h0020; #100;
A = 16'h00F6; B = 16'h0021; #100;
A = 16'h00F6; B = 16'h0022; #100;
A = 16'h00F6; B = 16'h0023; #100;
A = 16'h00F6; B = 16'h0024; #100;
A = 16'h00F6; B = 16'h0025; #100;
A = 16'h00F6; B = 16'h0026; #100;
A = 16'h00F6; B = 16'h0027; #100;
A = 16'h00F6; B = 16'h0028; #100;
A = 16'h00F6; B = 16'h0029; #100;
A = 16'h00F6; B = 16'h002A; #100;
A = 16'h00F6; B = 16'h002B; #100;
A = 16'h00F6; B = 16'h002C; #100;
A = 16'h00F6; B = 16'h002D; #100;
A = 16'h00F6; B = 16'h002E; #100;
A = 16'h00F6; B = 16'h002F; #100;
A = 16'h00F6; B = 16'h0030; #100;
A = 16'h00F6; B = 16'h0031; #100;
A = 16'h00F6; B = 16'h0032; #100;
A = 16'h00F6; B = 16'h0033; #100;
A = 16'h00F6; B = 16'h0034; #100;
A = 16'h00F6; B = 16'h0035; #100;
A = 16'h00F6; B = 16'h0036; #100;
A = 16'h00F6; B = 16'h0037; #100;
A = 16'h00F6; B = 16'h0038; #100;
A = 16'h00F6; B = 16'h0039; #100;
A = 16'h00F6; B = 16'h003A; #100;
A = 16'h00F6; B = 16'h003B; #100;
A = 16'h00F6; B = 16'h003C; #100;
A = 16'h00F6; B = 16'h003D; #100;
A = 16'h00F6; B = 16'h003E; #100;
A = 16'h00F6; B = 16'h003F; #100;
A = 16'h00F6; B = 16'h0040; #100;
A = 16'h00F6; B = 16'h0041; #100;
A = 16'h00F6; B = 16'h0042; #100;
A = 16'h00F6; B = 16'h0043; #100;
A = 16'h00F6; B = 16'h0044; #100;
A = 16'h00F6; B = 16'h0045; #100;
A = 16'h00F6; B = 16'h0046; #100;
A = 16'h00F6; B = 16'h0047; #100;
A = 16'h00F6; B = 16'h0048; #100;
A = 16'h00F6; B = 16'h0049; #100;
A = 16'h00F6; B = 16'h004A; #100;
A = 16'h00F6; B = 16'h004B; #100;
A = 16'h00F6; B = 16'h004C; #100;
A = 16'h00F6; B = 16'h004D; #100;
A = 16'h00F6; B = 16'h004E; #100;
A = 16'h00F6; B = 16'h004F; #100;
A = 16'h00F6; B = 16'h0050; #100;
A = 16'h00F6; B = 16'h0051; #100;
A = 16'h00F6; B = 16'h0052; #100;
A = 16'h00F6; B = 16'h0053; #100;
A = 16'h00F6; B = 16'h0054; #100;
A = 16'h00F6; B = 16'h0055; #100;
A = 16'h00F6; B = 16'h0056; #100;
A = 16'h00F6; B = 16'h0057; #100;
A = 16'h00F6; B = 16'h0058; #100;
A = 16'h00F6; B = 16'h0059; #100;
A = 16'h00F6; B = 16'h005A; #100;
A = 16'h00F6; B = 16'h005B; #100;
A = 16'h00F6; B = 16'h005C; #100;
A = 16'h00F6; B = 16'h005D; #100;
A = 16'h00F6; B = 16'h005E; #100;
A = 16'h00F6; B = 16'h005F; #100;
A = 16'h00F6; B = 16'h0060; #100;
A = 16'h00F6; B = 16'h0061; #100;
A = 16'h00F6; B = 16'h0062; #100;
A = 16'h00F6; B = 16'h0063; #100;
A = 16'h00F6; B = 16'h0064; #100;
A = 16'h00F6; B = 16'h0065; #100;
A = 16'h00F6; B = 16'h0066; #100;
A = 16'h00F6; B = 16'h0067; #100;
A = 16'h00F6; B = 16'h0068; #100;
A = 16'h00F6; B = 16'h0069; #100;
A = 16'h00F6; B = 16'h006A; #100;
A = 16'h00F6; B = 16'h006B; #100;
A = 16'h00F6; B = 16'h006C; #100;
A = 16'h00F6; B = 16'h006D; #100;
A = 16'h00F6; B = 16'h006E; #100;
A = 16'h00F6; B = 16'h006F; #100;
A = 16'h00F6; B = 16'h0070; #100;
A = 16'h00F6; B = 16'h0071; #100;
A = 16'h00F6; B = 16'h0072; #100;
A = 16'h00F6; B = 16'h0073; #100;
A = 16'h00F6; B = 16'h0074; #100;
A = 16'h00F6; B = 16'h0075; #100;
A = 16'h00F6; B = 16'h0076; #100;
A = 16'h00F6; B = 16'h0077; #100;
A = 16'h00F6; B = 16'h0078; #100;
A = 16'h00F6; B = 16'h0079; #100;
A = 16'h00F6; B = 16'h007A; #100;
A = 16'h00F6; B = 16'h007B; #100;
A = 16'h00F6; B = 16'h007C; #100;
A = 16'h00F6; B = 16'h007D; #100;
A = 16'h00F6; B = 16'h007E; #100;
A = 16'h00F6; B = 16'h007F; #100;
A = 16'h00F6; B = 16'h0080; #100;
A = 16'h00F6; B = 16'h0081; #100;
A = 16'h00F6; B = 16'h0082; #100;
A = 16'h00F6; B = 16'h0083; #100;
A = 16'h00F6; B = 16'h0084; #100;
A = 16'h00F6; B = 16'h0085; #100;
A = 16'h00F6; B = 16'h0086; #100;
A = 16'h00F6; B = 16'h0087; #100;
A = 16'h00F6; B = 16'h0088; #100;
A = 16'h00F6; B = 16'h0089; #100;
A = 16'h00F6; B = 16'h008A; #100;
A = 16'h00F6; B = 16'h008B; #100;
A = 16'h00F6; B = 16'h008C; #100;
A = 16'h00F6; B = 16'h008D; #100;
A = 16'h00F6; B = 16'h008E; #100;
A = 16'h00F6; B = 16'h008F; #100;
A = 16'h00F6; B = 16'h0090; #100;
A = 16'h00F6; B = 16'h0091; #100;
A = 16'h00F6; B = 16'h0092; #100;
A = 16'h00F6; B = 16'h0093; #100;
A = 16'h00F6; B = 16'h0094; #100;
A = 16'h00F6; B = 16'h0095; #100;
A = 16'h00F6; B = 16'h0096; #100;
A = 16'h00F6; B = 16'h0097; #100;
A = 16'h00F6; B = 16'h0098; #100;
A = 16'h00F6; B = 16'h0099; #100;
A = 16'h00F6; B = 16'h009A; #100;
A = 16'h00F6; B = 16'h009B; #100;
A = 16'h00F6; B = 16'h009C; #100;
A = 16'h00F6; B = 16'h009D; #100;
A = 16'h00F6; B = 16'h009E; #100;
A = 16'h00F6; B = 16'h009F; #100;
A = 16'h00F6; B = 16'h00A0; #100;
A = 16'h00F6; B = 16'h00A1; #100;
A = 16'h00F6; B = 16'h00A2; #100;
A = 16'h00F6; B = 16'h00A3; #100;
A = 16'h00F6; B = 16'h00A4; #100;
A = 16'h00F6; B = 16'h00A5; #100;
A = 16'h00F6; B = 16'h00A6; #100;
A = 16'h00F6; B = 16'h00A7; #100;
A = 16'h00F6; B = 16'h00A8; #100;
A = 16'h00F6; B = 16'h00A9; #100;
A = 16'h00F6; B = 16'h00AA; #100;
A = 16'h00F6; B = 16'h00AB; #100;
A = 16'h00F6; B = 16'h00AC; #100;
A = 16'h00F6; B = 16'h00AD; #100;
A = 16'h00F6; B = 16'h00AE; #100;
A = 16'h00F6; B = 16'h00AF; #100;
A = 16'h00F6; B = 16'h00B0; #100;
A = 16'h00F6; B = 16'h00B1; #100;
A = 16'h00F6; B = 16'h00B2; #100;
A = 16'h00F6; B = 16'h00B3; #100;
A = 16'h00F6; B = 16'h00B4; #100;
A = 16'h00F6; B = 16'h00B5; #100;
A = 16'h00F6; B = 16'h00B6; #100;
A = 16'h00F6; B = 16'h00B7; #100;
A = 16'h00F6; B = 16'h00B8; #100;
A = 16'h00F6; B = 16'h00B9; #100;
A = 16'h00F6; B = 16'h00BA; #100;
A = 16'h00F6; B = 16'h00BB; #100;
A = 16'h00F6; B = 16'h00BC; #100;
A = 16'h00F6; B = 16'h00BD; #100;
A = 16'h00F6; B = 16'h00BE; #100;
A = 16'h00F6; B = 16'h00BF; #100;
A = 16'h00F6; B = 16'h00C0; #100;
A = 16'h00F6; B = 16'h00C1; #100;
A = 16'h00F6; B = 16'h00C2; #100;
A = 16'h00F6; B = 16'h00C3; #100;
A = 16'h00F6; B = 16'h00C4; #100;
A = 16'h00F6; B = 16'h00C5; #100;
A = 16'h00F6; B = 16'h00C6; #100;
A = 16'h00F6; B = 16'h00C7; #100;
A = 16'h00F6; B = 16'h00C8; #100;
A = 16'h00F6; B = 16'h00C9; #100;
A = 16'h00F6; B = 16'h00CA; #100;
A = 16'h00F6; B = 16'h00CB; #100;
A = 16'h00F6; B = 16'h00CC; #100;
A = 16'h00F6; B = 16'h00CD; #100;
A = 16'h00F6; B = 16'h00CE; #100;
A = 16'h00F6; B = 16'h00CF; #100;
A = 16'h00F6; B = 16'h00D0; #100;
A = 16'h00F6; B = 16'h00D1; #100;
A = 16'h00F6; B = 16'h00D2; #100;
A = 16'h00F6; B = 16'h00D3; #100;
A = 16'h00F6; B = 16'h00D4; #100;
A = 16'h00F6; B = 16'h00D5; #100;
A = 16'h00F6; B = 16'h00D6; #100;
A = 16'h00F6; B = 16'h00D7; #100;
A = 16'h00F6; B = 16'h00D8; #100;
A = 16'h00F6; B = 16'h00D9; #100;
A = 16'h00F6; B = 16'h00DA; #100;
A = 16'h00F6; B = 16'h00DB; #100;
A = 16'h00F6; B = 16'h00DC; #100;
A = 16'h00F6; B = 16'h00DD; #100;
A = 16'h00F6; B = 16'h00DE; #100;
A = 16'h00F6; B = 16'h00DF; #100;
A = 16'h00F6; B = 16'h00E0; #100;
A = 16'h00F6; B = 16'h00E1; #100;
A = 16'h00F6; B = 16'h00E2; #100;
A = 16'h00F6; B = 16'h00E3; #100;
A = 16'h00F6; B = 16'h00E4; #100;
A = 16'h00F6; B = 16'h00E5; #100;
A = 16'h00F6; B = 16'h00E6; #100;
A = 16'h00F6; B = 16'h00E7; #100;
A = 16'h00F6; B = 16'h00E8; #100;
A = 16'h00F6; B = 16'h00E9; #100;
A = 16'h00F6; B = 16'h00EA; #100;
A = 16'h00F6; B = 16'h00EB; #100;
A = 16'h00F6; B = 16'h00EC; #100;
A = 16'h00F6; B = 16'h00ED; #100;
A = 16'h00F6; B = 16'h00EE; #100;
A = 16'h00F6; B = 16'h00EF; #100;
A = 16'h00F6; B = 16'h00F0; #100;
A = 16'h00F6; B = 16'h00F1; #100;
A = 16'h00F6; B = 16'h00F2; #100;
A = 16'h00F6; B = 16'h00F3; #100;
A = 16'h00F6; B = 16'h00F4; #100;
A = 16'h00F6; B = 16'h00F5; #100;
A = 16'h00F6; B = 16'h00F6; #100;
A = 16'h00F6; B = 16'h00F7; #100;
A = 16'h00F6; B = 16'h00F8; #100;
A = 16'h00F6; B = 16'h00F9; #100;
A = 16'h00F6; B = 16'h00FA; #100;
A = 16'h00F6; B = 16'h00FB; #100;
A = 16'h00F6; B = 16'h00FC; #100;
A = 16'h00F6; B = 16'h00FD; #100;
A = 16'h00F6; B = 16'h00FE; #100;
A = 16'h00F6; B = 16'h00FF; #100;
A = 16'h00F7; B = 16'h000; #100;
A = 16'h00F7; B = 16'h001; #100;
A = 16'h00F7; B = 16'h002; #100;
A = 16'h00F7; B = 16'h003; #100;
A = 16'h00F7; B = 16'h004; #100;
A = 16'h00F7; B = 16'h005; #100;
A = 16'h00F7; B = 16'h006; #100;
A = 16'h00F7; B = 16'h007; #100;
A = 16'h00F7; B = 16'h008; #100;
A = 16'h00F7; B = 16'h009; #100;
A = 16'h00F7; B = 16'h00A; #100;
A = 16'h00F7; B = 16'h00B; #100;
A = 16'h00F7; B = 16'h00C; #100;
A = 16'h00F7; B = 16'h00D; #100;
A = 16'h00F7; B = 16'h00E; #100;
A = 16'h00F7; B = 16'h00F; #100;
A = 16'h00F7; B = 16'h0010; #100;
A = 16'h00F7; B = 16'h0011; #100;
A = 16'h00F7; B = 16'h0012; #100;
A = 16'h00F7; B = 16'h0013; #100;
A = 16'h00F7; B = 16'h0014; #100;
A = 16'h00F7; B = 16'h0015; #100;
A = 16'h00F7; B = 16'h0016; #100;
A = 16'h00F7; B = 16'h0017; #100;
A = 16'h00F7; B = 16'h0018; #100;
A = 16'h00F7; B = 16'h0019; #100;
A = 16'h00F7; B = 16'h001A; #100;
A = 16'h00F7; B = 16'h001B; #100;
A = 16'h00F7; B = 16'h001C; #100;
A = 16'h00F7; B = 16'h001D; #100;
A = 16'h00F7; B = 16'h001E; #100;
A = 16'h00F7; B = 16'h001F; #100;
A = 16'h00F7; B = 16'h0020; #100;
A = 16'h00F7; B = 16'h0021; #100;
A = 16'h00F7; B = 16'h0022; #100;
A = 16'h00F7; B = 16'h0023; #100;
A = 16'h00F7; B = 16'h0024; #100;
A = 16'h00F7; B = 16'h0025; #100;
A = 16'h00F7; B = 16'h0026; #100;
A = 16'h00F7; B = 16'h0027; #100;
A = 16'h00F7; B = 16'h0028; #100;
A = 16'h00F7; B = 16'h0029; #100;
A = 16'h00F7; B = 16'h002A; #100;
A = 16'h00F7; B = 16'h002B; #100;
A = 16'h00F7; B = 16'h002C; #100;
A = 16'h00F7; B = 16'h002D; #100;
A = 16'h00F7; B = 16'h002E; #100;
A = 16'h00F7; B = 16'h002F; #100;
A = 16'h00F7; B = 16'h0030; #100;
A = 16'h00F7; B = 16'h0031; #100;
A = 16'h00F7; B = 16'h0032; #100;
A = 16'h00F7; B = 16'h0033; #100;
A = 16'h00F7; B = 16'h0034; #100;
A = 16'h00F7; B = 16'h0035; #100;
A = 16'h00F7; B = 16'h0036; #100;
A = 16'h00F7; B = 16'h0037; #100;
A = 16'h00F7; B = 16'h0038; #100;
A = 16'h00F7; B = 16'h0039; #100;
A = 16'h00F7; B = 16'h003A; #100;
A = 16'h00F7; B = 16'h003B; #100;
A = 16'h00F7; B = 16'h003C; #100;
A = 16'h00F7; B = 16'h003D; #100;
A = 16'h00F7; B = 16'h003E; #100;
A = 16'h00F7; B = 16'h003F; #100;
A = 16'h00F7; B = 16'h0040; #100;
A = 16'h00F7; B = 16'h0041; #100;
A = 16'h00F7; B = 16'h0042; #100;
A = 16'h00F7; B = 16'h0043; #100;
A = 16'h00F7; B = 16'h0044; #100;
A = 16'h00F7; B = 16'h0045; #100;
A = 16'h00F7; B = 16'h0046; #100;
A = 16'h00F7; B = 16'h0047; #100;
A = 16'h00F7; B = 16'h0048; #100;
A = 16'h00F7; B = 16'h0049; #100;
A = 16'h00F7; B = 16'h004A; #100;
A = 16'h00F7; B = 16'h004B; #100;
A = 16'h00F7; B = 16'h004C; #100;
A = 16'h00F7; B = 16'h004D; #100;
A = 16'h00F7; B = 16'h004E; #100;
A = 16'h00F7; B = 16'h004F; #100;
A = 16'h00F7; B = 16'h0050; #100;
A = 16'h00F7; B = 16'h0051; #100;
A = 16'h00F7; B = 16'h0052; #100;
A = 16'h00F7; B = 16'h0053; #100;
A = 16'h00F7; B = 16'h0054; #100;
A = 16'h00F7; B = 16'h0055; #100;
A = 16'h00F7; B = 16'h0056; #100;
A = 16'h00F7; B = 16'h0057; #100;
A = 16'h00F7; B = 16'h0058; #100;
A = 16'h00F7; B = 16'h0059; #100;
A = 16'h00F7; B = 16'h005A; #100;
A = 16'h00F7; B = 16'h005B; #100;
A = 16'h00F7; B = 16'h005C; #100;
A = 16'h00F7; B = 16'h005D; #100;
A = 16'h00F7; B = 16'h005E; #100;
A = 16'h00F7; B = 16'h005F; #100;
A = 16'h00F7; B = 16'h0060; #100;
A = 16'h00F7; B = 16'h0061; #100;
A = 16'h00F7; B = 16'h0062; #100;
A = 16'h00F7; B = 16'h0063; #100;
A = 16'h00F7; B = 16'h0064; #100;
A = 16'h00F7; B = 16'h0065; #100;
A = 16'h00F7; B = 16'h0066; #100;
A = 16'h00F7; B = 16'h0067; #100;
A = 16'h00F7; B = 16'h0068; #100;
A = 16'h00F7; B = 16'h0069; #100;
A = 16'h00F7; B = 16'h006A; #100;
A = 16'h00F7; B = 16'h006B; #100;
A = 16'h00F7; B = 16'h006C; #100;
A = 16'h00F7; B = 16'h006D; #100;
A = 16'h00F7; B = 16'h006E; #100;
A = 16'h00F7; B = 16'h006F; #100;
A = 16'h00F7; B = 16'h0070; #100;
A = 16'h00F7; B = 16'h0071; #100;
A = 16'h00F7; B = 16'h0072; #100;
A = 16'h00F7; B = 16'h0073; #100;
A = 16'h00F7; B = 16'h0074; #100;
A = 16'h00F7; B = 16'h0075; #100;
A = 16'h00F7; B = 16'h0076; #100;
A = 16'h00F7; B = 16'h0077; #100;
A = 16'h00F7; B = 16'h0078; #100;
A = 16'h00F7; B = 16'h0079; #100;
A = 16'h00F7; B = 16'h007A; #100;
A = 16'h00F7; B = 16'h007B; #100;
A = 16'h00F7; B = 16'h007C; #100;
A = 16'h00F7; B = 16'h007D; #100;
A = 16'h00F7; B = 16'h007E; #100;
A = 16'h00F7; B = 16'h007F; #100;
A = 16'h00F7; B = 16'h0080; #100;
A = 16'h00F7; B = 16'h0081; #100;
A = 16'h00F7; B = 16'h0082; #100;
A = 16'h00F7; B = 16'h0083; #100;
A = 16'h00F7; B = 16'h0084; #100;
A = 16'h00F7; B = 16'h0085; #100;
A = 16'h00F7; B = 16'h0086; #100;
A = 16'h00F7; B = 16'h0087; #100;
A = 16'h00F7; B = 16'h0088; #100;
A = 16'h00F7; B = 16'h0089; #100;
A = 16'h00F7; B = 16'h008A; #100;
A = 16'h00F7; B = 16'h008B; #100;
A = 16'h00F7; B = 16'h008C; #100;
A = 16'h00F7; B = 16'h008D; #100;
A = 16'h00F7; B = 16'h008E; #100;
A = 16'h00F7; B = 16'h008F; #100;
A = 16'h00F7; B = 16'h0090; #100;
A = 16'h00F7; B = 16'h0091; #100;
A = 16'h00F7; B = 16'h0092; #100;
A = 16'h00F7; B = 16'h0093; #100;
A = 16'h00F7; B = 16'h0094; #100;
A = 16'h00F7; B = 16'h0095; #100;
A = 16'h00F7; B = 16'h0096; #100;
A = 16'h00F7; B = 16'h0097; #100;
A = 16'h00F7; B = 16'h0098; #100;
A = 16'h00F7; B = 16'h0099; #100;
A = 16'h00F7; B = 16'h009A; #100;
A = 16'h00F7; B = 16'h009B; #100;
A = 16'h00F7; B = 16'h009C; #100;
A = 16'h00F7; B = 16'h009D; #100;
A = 16'h00F7; B = 16'h009E; #100;
A = 16'h00F7; B = 16'h009F; #100;
A = 16'h00F7; B = 16'h00A0; #100;
A = 16'h00F7; B = 16'h00A1; #100;
A = 16'h00F7; B = 16'h00A2; #100;
A = 16'h00F7; B = 16'h00A3; #100;
A = 16'h00F7; B = 16'h00A4; #100;
A = 16'h00F7; B = 16'h00A5; #100;
A = 16'h00F7; B = 16'h00A6; #100;
A = 16'h00F7; B = 16'h00A7; #100;
A = 16'h00F7; B = 16'h00A8; #100;
A = 16'h00F7; B = 16'h00A9; #100;
A = 16'h00F7; B = 16'h00AA; #100;
A = 16'h00F7; B = 16'h00AB; #100;
A = 16'h00F7; B = 16'h00AC; #100;
A = 16'h00F7; B = 16'h00AD; #100;
A = 16'h00F7; B = 16'h00AE; #100;
A = 16'h00F7; B = 16'h00AF; #100;
A = 16'h00F7; B = 16'h00B0; #100;
A = 16'h00F7; B = 16'h00B1; #100;
A = 16'h00F7; B = 16'h00B2; #100;
A = 16'h00F7; B = 16'h00B3; #100;
A = 16'h00F7; B = 16'h00B4; #100;
A = 16'h00F7; B = 16'h00B5; #100;
A = 16'h00F7; B = 16'h00B6; #100;
A = 16'h00F7; B = 16'h00B7; #100;
A = 16'h00F7; B = 16'h00B8; #100;
A = 16'h00F7; B = 16'h00B9; #100;
A = 16'h00F7; B = 16'h00BA; #100;
A = 16'h00F7; B = 16'h00BB; #100;
A = 16'h00F7; B = 16'h00BC; #100;
A = 16'h00F7; B = 16'h00BD; #100;
A = 16'h00F7; B = 16'h00BE; #100;
A = 16'h00F7; B = 16'h00BF; #100;
A = 16'h00F7; B = 16'h00C0; #100;
A = 16'h00F7; B = 16'h00C1; #100;
A = 16'h00F7; B = 16'h00C2; #100;
A = 16'h00F7; B = 16'h00C3; #100;
A = 16'h00F7; B = 16'h00C4; #100;
A = 16'h00F7; B = 16'h00C5; #100;
A = 16'h00F7; B = 16'h00C6; #100;
A = 16'h00F7; B = 16'h00C7; #100;
A = 16'h00F7; B = 16'h00C8; #100;
A = 16'h00F7; B = 16'h00C9; #100;
A = 16'h00F7; B = 16'h00CA; #100;
A = 16'h00F7; B = 16'h00CB; #100;
A = 16'h00F7; B = 16'h00CC; #100;
A = 16'h00F7; B = 16'h00CD; #100;
A = 16'h00F7; B = 16'h00CE; #100;
A = 16'h00F7; B = 16'h00CF; #100;
A = 16'h00F7; B = 16'h00D0; #100;
A = 16'h00F7; B = 16'h00D1; #100;
A = 16'h00F7; B = 16'h00D2; #100;
A = 16'h00F7; B = 16'h00D3; #100;
A = 16'h00F7; B = 16'h00D4; #100;
A = 16'h00F7; B = 16'h00D5; #100;
A = 16'h00F7; B = 16'h00D6; #100;
A = 16'h00F7; B = 16'h00D7; #100;
A = 16'h00F7; B = 16'h00D8; #100;
A = 16'h00F7; B = 16'h00D9; #100;
A = 16'h00F7; B = 16'h00DA; #100;
A = 16'h00F7; B = 16'h00DB; #100;
A = 16'h00F7; B = 16'h00DC; #100;
A = 16'h00F7; B = 16'h00DD; #100;
A = 16'h00F7; B = 16'h00DE; #100;
A = 16'h00F7; B = 16'h00DF; #100;
A = 16'h00F7; B = 16'h00E0; #100;
A = 16'h00F7; B = 16'h00E1; #100;
A = 16'h00F7; B = 16'h00E2; #100;
A = 16'h00F7; B = 16'h00E3; #100;
A = 16'h00F7; B = 16'h00E4; #100;
A = 16'h00F7; B = 16'h00E5; #100;
A = 16'h00F7; B = 16'h00E6; #100;
A = 16'h00F7; B = 16'h00E7; #100;
A = 16'h00F7; B = 16'h00E8; #100;
A = 16'h00F7; B = 16'h00E9; #100;
A = 16'h00F7; B = 16'h00EA; #100;
A = 16'h00F7; B = 16'h00EB; #100;
A = 16'h00F7; B = 16'h00EC; #100;
A = 16'h00F7; B = 16'h00ED; #100;
A = 16'h00F7; B = 16'h00EE; #100;
A = 16'h00F7; B = 16'h00EF; #100;
A = 16'h00F7; B = 16'h00F0; #100;
A = 16'h00F7; B = 16'h00F1; #100;
A = 16'h00F7; B = 16'h00F2; #100;
A = 16'h00F7; B = 16'h00F3; #100;
A = 16'h00F7; B = 16'h00F4; #100;
A = 16'h00F7; B = 16'h00F5; #100;
A = 16'h00F7; B = 16'h00F6; #100;
A = 16'h00F7; B = 16'h00F7; #100;
A = 16'h00F7; B = 16'h00F8; #100;
A = 16'h00F7; B = 16'h00F9; #100;
A = 16'h00F7; B = 16'h00FA; #100;
A = 16'h00F7; B = 16'h00FB; #100;
A = 16'h00F7; B = 16'h00FC; #100;
A = 16'h00F7; B = 16'h00FD; #100;
A = 16'h00F7; B = 16'h00FE; #100;
A = 16'h00F7; B = 16'h00FF; #100;
A = 16'h00F8; B = 16'h000; #100;
A = 16'h00F8; B = 16'h001; #100;
A = 16'h00F8; B = 16'h002; #100;
A = 16'h00F8; B = 16'h003; #100;
A = 16'h00F8; B = 16'h004; #100;
A = 16'h00F8; B = 16'h005; #100;
A = 16'h00F8; B = 16'h006; #100;
A = 16'h00F8; B = 16'h007; #100;
A = 16'h00F8; B = 16'h008; #100;
A = 16'h00F8; B = 16'h009; #100;
A = 16'h00F8; B = 16'h00A; #100;
A = 16'h00F8; B = 16'h00B; #100;
A = 16'h00F8; B = 16'h00C; #100;
A = 16'h00F8; B = 16'h00D; #100;
A = 16'h00F8; B = 16'h00E; #100;
A = 16'h00F8; B = 16'h00F; #100;
A = 16'h00F8; B = 16'h0010; #100;
A = 16'h00F8; B = 16'h0011; #100;
A = 16'h00F8; B = 16'h0012; #100;
A = 16'h00F8; B = 16'h0013; #100;
A = 16'h00F8; B = 16'h0014; #100;
A = 16'h00F8; B = 16'h0015; #100;
A = 16'h00F8; B = 16'h0016; #100;
A = 16'h00F8; B = 16'h0017; #100;
A = 16'h00F8; B = 16'h0018; #100;
A = 16'h00F8; B = 16'h0019; #100;
A = 16'h00F8; B = 16'h001A; #100;
A = 16'h00F8; B = 16'h001B; #100;
A = 16'h00F8; B = 16'h001C; #100;
A = 16'h00F8; B = 16'h001D; #100;
A = 16'h00F8; B = 16'h001E; #100;
A = 16'h00F8; B = 16'h001F; #100;
A = 16'h00F8; B = 16'h0020; #100;
A = 16'h00F8; B = 16'h0021; #100;
A = 16'h00F8; B = 16'h0022; #100;
A = 16'h00F8; B = 16'h0023; #100;
A = 16'h00F8; B = 16'h0024; #100;
A = 16'h00F8; B = 16'h0025; #100;
A = 16'h00F8; B = 16'h0026; #100;
A = 16'h00F8; B = 16'h0027; #100;
A = 16'h00F8; B = 16'h0028; #100;
A = 16'h00F8; B = 16'h0029; #100;
A = 16'h00F8; B = 16'h002A; #100;
A = 16'h00F8; B = 16'h002B; #100;
A = 16'h00F8; B = 16'h002C; #100;
A = 16'h00F8; B = 16'h002D; #100;
A = 16'h00F8; B = 16'h002E; #100;
A = 16'h00F8; B = 16'h002F; #100;
A = 16'h00F8; B = 16'h0030; #100;
A = 16'h00F8; B = 16'h0031; #100;
A = 16'h00F8; B = 16'h0032; #100;
A = 16'h00F8; B = 16'h0033; #100;
A = 16'h00F8; B = 16'h0034; #100;
A = 16'h00F8; B = 16'h0035; #100;
A = 16'h00F8; B = 16'h0036; #100;
A = 16'h00F8; B = 16'h0037; #100;
A = 16'h00F8; B = 16'h0038; #100;
A = 16'h00F8; B = 16'h0039; #100;
A = 16'h00F8; B = 16'h003A; #100;
A = 16'h00F8; B = 16'h003B; #100;
A = 16'h00F8; B = 16'h003C; #100;
A = 16'h00F8; B = 16'h003D; #100;
A = 16'h00F8; B = 16'h003E; #100;
A = 16'h00F8; B = 16'h003F; #100;
A = 16'h00F8; B = 16'h0040; #100;
A = 16'h00F8; B = 16'h0041; #100;
A = 16'h00F8; B = 16'h0042; #100;
A = 16'h00F8; B = 16'h0043; #100;
A = 16'h00F8; B = 16'h0044; #100;
A = 16'h00F8; B = 16'h0045; #100;
A = 16'h00F8; B = 16'h0046; #100;
A = 16'h00F8; B = 16'h0047; #100;
A = 16'h00F8; B = 16'h0048; #100;
A = 16'h00F8; B = 16'h0049; #100;
A = 16'h00F8; B = 16'h004A; #100;
A = 16'h00F8; B = 16'h004B; #100;
A = 16'h00F8; B = 16'h004C; #100;
A = 16'h00F8; B = 16'h004D; #100;
A = 16'h00F8; B = 16'h004E; #100;
A = 16'h00F8; B = 16'h004F; #100;
A = 16'h00F8; B = 16'h0050; #100;
A = 16'h00F8; B = 16'h0051; #100;
A = 16'h00F8; B = 16'h0052; #100;
A = 16'h00F8; B = 16'h0053; #100;
A = 16'h00F8; B = 16'h0054; #100;
A = 16'h00F8; B = 16'h0055; #100;
A = 16'h00F8; B = 16'h0056; #100;
A = 16'h00F8; B = 16'h0057; #100;
A = 16'h00F8; B = 16'h0058; #100;
A = 16'h00F8; B = 16'h0059; #100;
A = 16'h00F8; B = 16'h005A; #100;
A = 16'h00F8; B = 16'h005B; #100;
A = 16'h00F8; B = 16'h005C; #100;
A = 16'h00F8; B = 16'h005D; #100;
A = 16'h00F8; B = 16'h005E; #100;
A = 16'h00F8; B = 16'h005F; #100;
A = 16'h00F8; B = 16'h0060; #100;
A = 16'h00F8; B = 16'h0061; #100;
A = 16'h00F8; B = 16'h0062; #100;
A = 16'h00F8; B = 16'h0063; #100;
A = 16'h00F8; B = 16'h0064; #100;
A = 16'h00F8; B = 16'h0065; #100;
A = 16'h00F8; B = 16'h0066; #100;
A = 16'h00F8; B = 16'h0067; #100;
A = 16'h00F8; B = 16'h0068; #100;
A = 16'h00F8; B = 16'h0069; #100;
A = 16'h00F8; B = 16'h006A; #100;
A = 16'h00F8; B = 16'h006B; #100;
A = 16'h00F8; B = 16'h006C; #100;
A = 16'h00F8; B = 16'h006D; #100;
A = 16'h00F8; B = 16'h006E; #100;
A = 16'h00F8; B = 16'h006F; #100;
A = 16'h00F8; B = 16'h0070; #100;
A = 16'h00F8; B = 16'h0071; #100;
A = 16'h00F8; B = 16'h0072; #100;
A = 16'h00F8; B = 16'h0073; #100;
A = 16'h00F8; B = 16'h0074; #100;
A = 16'h00F8; B = 16'h0075; #100;
A = 16'h00F8; B = 16'h0076; #100;
A = 16'h00F8; B = 16'h0077; #100;
A = 16'h00F8; B = 16'h0078; #100;
A = 16'h00F8; B = 16'h0079; #100;
A = 16'h00F8; B = 16'h007A; #100;
A = 16'h00F8; B = 16'h007B; #100;
A = 16'h00F8; B = 16'h007C; #100;
A = 16'h00F8; B = 16'h007D; #100;
A = 16'h00F8; B = 16'h007E; #100;
A = 16'h00F8; B = 16'h007F; #100;
A = 16'h00F8; B = 16'h0080; #100;
A = 16'h00F8; B = 16'h0081; #100;
A = 16'h00F8; B = 16'h0082; #100;
A = 16'h00F8; B = 16'h0083; #100;
A = 16'h00F8; B = 16'h0084; #100;
A = 16'h00F8; B = 16'h0085; #100;
A = 16'h00F8; B = 16'h0086; #100;
A = 16'h00F8; B = 16'h0087; #100;
A = 16'h00F8; B = 16'h0088; #100;
A = 16'h00F8; B = 16'h0089; #100;
A = 16'h00F8; B = 16'h008A; #100;
A = 16'h00F8; B = 16'h008B; #100;
A = 16'h00F8; B = 16'h008C; #100;
A = 16'h00F8; B = 16'h008D; #100;
A = 16'h00F8; B = 16'h008E; #100;
A = 16'h00F8; B = 16'h008F; #100;
A = 16'h00F8; B = 16'h0090; #100;
A = 16'h00F8; B = 16'h0091; #100;
A = 16'h00F8; B = 16'h0092; #100;
A = 16'h00F8; B = 16'h0093; #100;
A = 16'h00F8; B = 16'h0094; #100;
A = 16'h00F8; B = 16'h0095; #100;
A = 16'h00F8; B = 16'h0096; #100;
A = 16'h00F8; B = 16'h0097; #100;
A = 16'h00F8; B = 16'h0098; #100;
A = 16'h00F8; B = 16'h0099; #100;
A = 16'h00F8; B = 16'h009A; #100;
A = 16'h00F8; B = 16'h009B; #100;
A = 16'h00F8; B = 16'h009C; #100;
A = 16'h00F8; B = 16'h009D; #100;
A = 16'h00F8; B = 16'h009E; #100;
A = 16'h00F8; B = 16'h009F; #100;
A = 16'h00F8; B = 16'h00A0; #100;
A = 16'h00F8; B = 16'h00A1; #100;
A = 16'h00F8; B = 16'h00A2; #100;
A = 16'h00F8; B = 16'h00A3; #100;
A = 16'h00F8; B = 16'h00A4; #100;
A = 16'h00F8; B = 16'h00A5; #100;
A = 16'h00F8; B = 16'h00A6; #100;
A = 16'h00F8; B = 16'h00A7; #100;
A = 16'h00F8; B = 16'h00A8; #100;
A = 16'h00F8; B = 16'h00A9; #100;
A = 16'h00F8; B = 16'h00AA; #100;
A = 16'h00F8; B = 16'h00AB; #100;
A = 16'h00F8; B = 16'h00AC; #100;
A = 16'h00F8; B = 16'h00AD; #100;
A = 16'h00F8; B = 16'h00AE; #100;
A = 16'h00F8; B = 16'h00AF; #100;
A = 16'h00F8; B = 16'h00B0; #100;
A = 16'h00F8; B = 16'h00B1; #100;
A = 16'h00F8; B = 16'h00B2; #100;
A = 16'h00F8; B = 16'h00B3; #100;
A = 16'h00F8; B = 16'h00B4; #100;
A = 16'h00F8; B = 16'h00B5; #100;
A = 16'h00F8; B = 16'h00B6; #100;
A = 16'h00F8; B = 16'h00B7; #100;
A = 16'h00F8; B = 16'h00B8; #100;
A = 16'h00F8; B = 16'h00B9; #100;
A = 16'h00F8; B = 16'h00BA; #100;
A = 16'h00F8; B = 16'h00BB; #100;
A = 16'h00F8; B = 16'h00BC; #100;
A = 16'h00F8; B = 16'h00BD; #100;
A = 16'h00F8; B = 16'h00BE; #100;
A = 16'h00F8; B = 16'h00BF; #100;
A = 16'h00F8; B = 16'h00C0; #100;
A = 16'h00F8; B = 16'h00C1; #100;
A = 16'h00F8; B = 16'h00C2; #100;
A = 16'h00F8; B = 16'h00C3; #100;
A = 16'h00F8; B = 16'h00C4; #100;
A = 16'h00F8; B = 16'h00C5; #100;
A = 16'h00F8; B = 16'h00C6; #100;
A = 16'h00F8; B = 16'h00C7; #100;
A = 16'h00F8; B = 16'h00C8; #100;
A = 16'h00F8; B = 16'h00C9; #100;
A = 16'h00F8; B = 16'h00CA; #100;
A = 16'h00F8; B = 16'h00CB; #100;
A = 16'h00F8; B = 16'h00CC; #100;
A = 16'h00F8; B = 16'h00CD; #100;
A = 16'h00F8; B = 16'h00CE; #100;
A = 16'h00F8; B = 16'h00CF; #100;
A = 16'h00F8; B = 16'h00D0; #100;
A = 16'h00F8; B = 16'h00D1; #100;
A = 16'h00F8; B = 16'h00D2; #100;
A = 16'h00F8; B = 16'h00D3; #100;
A = 16'h00F8; B = 16'h00D4; #100;
A = 16'h00F8; B = 16'h00D5; #100;
A = 16'h00F8; B = 16'h00D6; #100;
A = 16'h00F8; B = 16'h00D7; #100;
A = 16'h00F8; B = 16'h00D8; #100;
A = 16'h00F8; B = 16'h00D9; #100;
A = 16'h00F8; B = 16'h00DA; #100;
A = 16'h00F8; B = 16'h00DB; #100;
A = 16'h00F8; B = 16'h00DC; #100;
A = 16'h00F8; B = 16'h00DD; #100;
A = 16'h00F8; B = 16'h00DE; #100;
A = 16'h00F8; B = 16'h00DF; #100;
A = 16'h00F8; B = 16'h00E0; #100;
A = 16'h00F8; B = 16'h00E1; #100;
A = 16'h00F8; B = 16'h00E2; #100;
A = 16'h00F8; B = 16'h00E3; #100;
A = 16'h00F8; B = 16'h00E4; #100;
A = 16'h00F8; B = 16'h00E5; #100;
A = 16'h00F8; B = 16'h00E6; #100;
A = 16'h00F8; B = 16'h00E7; #100;
A = 16'h00F8; B = 16'h00E8; #100;
A = 16'h00F8; B = 16'h00E9; #100;
A = 16'h00F8; B = 16'h00EA; #100;
A = 16'h00F8; B = 16'h00EB; #100;
A = 16'h00F8; B = 16'h00EC; #100;
A = 16'h00F8; B = 16'h00ED; #100;
A = 16'h00F8; B = 16'h00EE; #100;
A = 16'h00F8; B = 16'h00EF; #100;
A = 16'h00F8; B = 16'h00F0; #100;
A = 16'h00F8; B = 16'h00F1; #100;
A = 16'h00F8; B = 16'h00F2; #100;
A = 16'h00F8; B = 16'h00F3; #100;
A = 16'h00F8; B = 16'h00F4; #100;
A = 16'h00F8; B = 16'h00F5; #100;
A = 16'h00F8; B = 16'h00F6; #100;
A = 16'h00F8; B = 16'h00F7; #100;
A = 16'h00F8; B = 16'h00F8; #100;
A = 16'h00F8; B = 16'h00F9; #100;
A = 16'h00F8; B = 16'h00FA; #100;
A = 16'h00F8; B = 16'h00FB; #100;
A = 16'h00F8; B = 16'h00FC; #100;
A = 16'h00F8; B = 16'h00FD; #100;
A = 16'h00F8; B = 16'h00FE; #100;
A = 16'h00F8; B = 16'h00FF; #100;
A = 16'h00F9; B = 16'h000; #100;
A = 16'h00F9; B = 16'h001; #100;
A = 16'h00F9; B = 16'h002; #100;
A = 16'h00F9; B = 16'h003; #100;
A = 16'h00F9; B = 16'h004; #100;
A = 16'h00F9; B = 16'h005; #100;
A = 16'h00F9; B = 16'h006; #100;
A = 16'h00F9; B = 16'h007; #100;
A = 16'h00F9; B = 16'h008; #100;
A = 16'h00F9; B = 16'h009; #100;
A = 16'h00F9; B = 16'h00A; #100;
A = 16'h00F9; B = 16'h00B; #100;
A = 16'h00F9; B = 16'h00C; #100;
A = 16'h00F9; B = 16'h00D; #100;
A = 16'h00F9; B = 16'h00E; #100;
A = 16'h00F9; B = 16'h00F; #100;
A = 16'h00F9; B = 16'h0010; #100;
A = 16'h00F9; B = 16'h0011; #100;
A = 16'h00F9; B = 16'h0012; #100;
A = 16'h00F9; B = 16'h0013; #100;
A = 16'h00F9; B = 16'h0014; #100;
A = 16'h00F9; B = 16'h0015; #100;
A = 16'h00F9; B = 16'h0016; #100;
A = 16'h00F9; B = 16'h0017; #100;
A = 16'h00F9; B = 16'h0018; #100;
A = 16'h00F9; B = 16'h0019; #100;
A = 16'h00F9; B = 16'h001A; #100;
A = 16'h00F9; B = 16'h001B; #100;
A = 16'h00F9; B = 16'h001C; #100;
A = 16'h00F9; B = 16'h001D; #100;
A = 16'h00F9; B = 16'h001E; #100;
A = 16'h00F9; B = 16'h001F; #100;
A = 16'h00F9; B = 16'h0020; #100;
A = 16'h00F9; B = 16'h0021; #100;
A = 16'h00F9; B = 16'h0022; #100;
A = 16'h00F9; B = 16'h0023; #100;
A = 16'h00F9; B = 16'h0024; #100;
A = 16'h00F9; B = 16'h0025; #100;
A = 16'h00F9; B = 16'h0026; #100;
A = 16'h00F9; B = 16'h0027; #100;
A = 16'h00F9; B = 16'h0028; #100;
A = 16'h00F9; B = 16'h0029; #100;
A = 16'h00F9; B = 16'h002A; #100;
A = 16'h00F9; B = 16'h002B; #100;
A = 16'h00F9; B = 16'h002C; #100;
A = 16'h00F9; B = 16'h002D; #100;
A = 16'h00F9; B = 16'h002E; #100;
A = 16'h00F9; B = 16'h002F; #100;
A = 16'h00F9; B = 16'h0030; #100;
A = 16'h00F9; B = 16'h0031; #100;
A = 16'h00F9; B = 16'h0032; #100;
A = 16'h00F9; B = 16'h0033; #100;
A = 16'h00F9; B = 16'h0034; #100;
A = 16'h00F9; B = 16'h0035; #100;
A = 16'h00F9; B = 16'h0036; #100;
A = 16'h00F9; B = 16'h0037; #100;
A = 16'h00F9; B = 16'h0038; #100;
A = 16'h00F9; B = 16'h0039; #100;
A = 16'h00F9; B = 16'h003A; #100;
A = 16'h00F9; B = 16'h003B; #100;
A = 16'h00F9; B = 16'h003C; #100;
A = 16'h00F9; B = 16'h003D; #100;
A = 16'h00F9; B = 16'h003E; #100;
A = 16'h00F9; B = 16'h003F; #100;
A = 16'h00F9; B = 16'h0040; #100;
A = 16'h00F9; B = 16'h0041; #100;
A = 16'h00F9; B = 16'h0042; #100;
A = 16'h00F9; B = 16'h0043; #100;
A = 16'h00F9; B = 16'h0044; #100;
A = 16'h00F9; B = 16'h0045; #100;
A = 16'h00F9; B = 16'h0046; #100;
A = 16'h00F9; B = 16'h0047; #100;
A = 16'h00F9; B = 16'h0048; #100;
A = 16'h00F9; B = 16'h0049; #100;
A = 16'h00F9; B = 16'h004A; #100;
A = 16'h00F9; B = 16'h004B; #100;
A = 16'h00F9; B = 16'h004C; #100;
A = 16'h00F9; B = 16'h004D; #100;
A = 16'h00F9; B = 16'h004E; #100;
A = 16'h00F9; B = 16'h004F; #100;
A = 16'h00F9; B = 16'h0050; #100;
A = 16'h00F9; B = 16'h0051; #100;
A = 16'h00F9; B = 16'h0052; #100;
A = 16'h00F9; B = 16'h0053; #100;
A = 16'h00F9; B = 16'h0054; #100;
A = 16'h00F9; B = 16'h0055; #100;
A = 16'h00F9; B = 16'h0056; #100;
A = 16'h00F9; B = 16'h0057; #100;
A = 16'h00F9; B = 16'h0058; #100;
A = 16'h00F9; B = 16'h0059; #100;
A = 16'h00F9; B = 16'h005A; #100;
A = 16'h00F9; B = 16'h005B; #100;
A = 16'h00F9; B = 16'h005C; #100;
A = 16'h00F9; B = 16'h005D; #100;
A = 16'h00F9; B = 16'h005E; #100;
A = 16'h00F9; B = 16'h005F; #100;
A = 16'h00F9; B = 16'h0060; #100;
A = 16'h00F9; B = 16'h0061; #100;
A = 16'h00F9; B = 16'h0062; #100;
A = 16'h00F9; B = 16'h0063; #100;
A = 16'h00F9; B = 16'h0064; #100;
A = 16'h00F9; B = 16'h0065; #100;
A = 16'h00F9; B = 16'h0066; #100;
A = 16'h00F9; B = 16'h0067; #100;
A = 16'h00F9; B = 16'h0068; #100;
A = 16'h00F9; B = 16'h0069; #100;
A = 16'h00F9; B = 16'h006A; #100;
A = 16'h00F9; B = 16'h006B; #100;
A = 16'h00F9; B = 16'h006C; #100;
A = 16'h00F9; B = 16'h006D; #100;
A = 16'h00F9; B = 16'h006E; #100;
A = 16'h00F9; B = 16'h006F; #100;
A = 16'h00F9; B = 16'h0070; #100;
A = 16'h00F9; B = 16'h0071; #100;
A = 16'h00F9; B = 16'h0072; #100;
A = 16'h00F9; B = 16'h0073; #100;
A = 16'h00F9; B = 16'h0074; #100;
A = 16'h00F9; B = 16'h0075; #100;
A = 16'h00F9; B = 16'h0076; #100;
A = 16'h00F9; B = 16'h0077; #100;
A = 16'h00F9; B = 16'h0078; #100;
A = 16'h00F9; B = 16'h0079; #100;
A = 16'h00F9; B = 16'h007A; #100;
A = 16'h00F9; B = 16'h007B; #100;
A = 16'h00F9; B = 16'h007C; #100;
A = 16'h00F9; B = 16'h007D; #100;
A = 16'h00F9; B = 16'h007E; #100;
A = 16'h00F9; B = 16'h007F; #100;
A = 16'h00F9; B = 16'h0080; #100;
A = 16'h00F9; B = 16'h0081; #100;
A = 16'h00F9; B = 16'h0082; #100;
A = 16'h00F9; B = 16'h0083; #100;
A = 16'h00F9; B = 16'h0084; #100;
A = 16'h00F9; B = 16'h0085; #100;
A = 16'h00F9; B = 16'h0086; #100;
A = 16'h00F9; B = 16'h0087; #100;
A = 16'h00F9; B = 16'h0088; #100;
A = 16'h00F9; B = 16'h0089; #100;
A = 16'h00F9; B = 16'h008A; #100;
A = 16'h00F9; B = 16'h008B; #100;
A = 16'h00F9; B = 16'h008C; #100;
A = 16'h00F9; B = 16'h008D; #100;
A = 16'h00F9; B = 16'h008E; #100;
A = 16'h00F9; B = 16'h008F; #100;
A = 16'h00F9; B = 16'h0090; #100;
A = 16'h00F9; B = 16'h0091; #100;
A = 16'h00F9; B = 16'h0092; #100;
A = 16'h00F9; B = 16'h0093; #100;
A = 16'h00F9; B = 16'h0094; #100;
A = 16'h00F9; B = 16'h0095; #100;
A = 16'h00F9; B = 16'h0096; #100;
A = 16'h00F9; B = 16'h0097; #100;
A = 16'h00F9; B = 16'h0098; #100;
A = 16'h00F9; B = 16'h0099; #100;
A = 16'h00F9; B = 16'h009A; #100;
A = 16'h00F9; B = 16'h009B; #100;
A = 16'h00F9; B = 16'h009C; #100;
A = 16'h00F9; B = 16'h009D; #100;
A = 16'h00F9; B = 16'h009E; #100;
A = 16'h00F9; B = 16'h009F; #100;
A = 16'h00F9; B = 16'h00A0; #100;
A = 16'h00F9; B = 16'h00A1; #100;
A = 16'h00F9; B = 16'h00A2; #100;
A = 16'h00F9; B = 16'h00A3; #100;
A = 16'h00F9; B = 16'h00A4; #100;
A = 16'h00F9; B = 16'h00A5; #100;
A = 16'h00F9; B = 16'h00A6; #100;
A = 16'h00F9; B = 16'h00A7; #100;
A = 16'h00F9; B = 16'h00A8; #100;
A = 16'h00F9; B = 16'h00A9; #100;
A = 16'h00F9; B = 16'h00AA; #100;
A = 16'h00F9; B = 16'h00AB; #100;
A = 16'h00F9; B = 16'h00AC; #100;
A = 16'h00F9; B = 16'h00AD; #100;
A = 16'h00F9; B = 16'h00AE; #100;
A = 16'h00F9; B = 16'h00AF; #100;
A = 16'h00F9; B = 16'h00B0; #100;
A = 16'h00F9; B = 16'h00B1; #100;
A = 16'h00F9; B = 16'h00B2; #100;
A = 16'h00F9; B = 16'h00B3; #100;
A = 16'h00F9; B = 16'h00B4; #100;
A = 16'h00F9; B = 16'h00B5; #100;
A = 16'h00F9; B = 16'h00B6; #100;
A = 16'h00F9; B = 16'h00B7; #100;
A = 16'h00F9; B = 16'h00B8; #100;
A = 16'h00F9; B = 16'h00B9; #100;
A = 16'h00F9; B = 16'h00BA; #100;
A = 16'h00F9; B = 16'h00BB; #100;
A = 16'h00F9; B = 16'h00BC; #100;
A = 16'h00F9; B = 16'h00BD; #100;
A = 16'h00F9; B = 16'h00BE; #100;
A = 16'h00F9; B = 16'h00BF; #100;
A = 16'h00F9; B = 16'h00C0; #100;
A = 16'h00F9; B = 16'h00C1; #100;
A = 16'h00F9; B = 16'h00C2; #100;
A = 16'h00F9; B = 16'h00C3; #100;
A = 16'h00F9; B = 16'h00C4; #100;
A = 16'h00F9; B = 16'h00C5; #100;
A = 16'h00F9; B = 16'h00C6; #100;
A = 16'h00F9; B = 16'h00C7; #100;
A = 16'h00F9; B = 16'h00C8; #100;
A = 16'h00F9; B = 16'h00C9; #100;
A = 16'h00F9; B = 16'h00CA; #100;
A = 16'h00F9; B = 16'h00CB; #100;
A = 16'h00F9; B = 16'h00CC; #100;
A = 16'h00F9; B = 16'h00CD; #100;
A = 16'h00F9; B = 16'h00CE; #100;
A = 16'h00F9; B = 16'h00CF; #100;
A = 16'h00F9; B = 16'h00D0; #100;
A = 16'h00F9; B = 16'h00D1; #100;
A = 16'h00F9; B = 16'h00D2; #100;
A = 16'h00F9; B = 16'h00D3; #100;
A = 16'h00F9; B = 16'h00D4; #100;
A = 16'h00F9; B = 16'h00D5; #100;
A = 16'h00F9; B = 16'h00D6; #100;
A = 16'h00F9; B = 16'h00D7; #100;
A = 16'h00F9; B = 16'h00D8; #100;
A = 16'h00F9; B = 16'h00D9; #100;
A = 16'h00F9; B = 16'h00DA; #100;
A = 16'h00F9; B = 16'h00DB; #100;
A = 16'h00F9; B = 16'h00DC; #100;
A = 16'h00F9; B = 16'h00DD; #100;
A = 16'h00F9; B = 16'h00DE; #100;
A = 16'h00F9; B = 16'h00DF; #100;
A = 16'h00F9; B = 16'h00E0; #100;
A = 16'h00F9; B = 16'h00E1; #100;
A = 16'h00F9; B = 16'h00E2; #100;
A = 16'h00F9; B = 16'h00E3; #100;
A = 16'h00F9; B = 16'h00E4; #100;
A = 16'h00F9; B = 16'h00E5; #100;
A = 16'h00F9; B = 16'h00E6; #100;
A = 16'h00F9; B = 16'h00E7; #100;
A = 16'h00F9; B = 16'h00E8; #100;
A = 16'h00F9; B = 16'h00E9; #100;
A = 16'h00F9; B = 16'h00EA; #100;
A = 16'h00F9; B = 16'h00EB; #100;
A = 16'h00F9; B = 16'h00EC; #100;
A = 16'h00F9; B = 16'h00ED; #100;
A = 16'h00F9; B = 16'h00EE; #100;
A = 16'h00F9; B = 16'h00EF; #100;
A = 16'h00F9; B = 16'h00F0; #100;
A = 16'h00F9; B = 16'h00F1; #100;
A = 16'h00F9; B = 16'h00F2; #100;
A = 16'h00F9; B = 16'h00F3; #100;
A = 16'h00F9; B = 16'h00F4; #100;
A = 16'h00F9; B = 16'h00F5; #100;
A = 16'h00F9; B = 16'h00F6; #100;
A = 16'h00F9; B = 16'h00F7; #100;
A = 16'h00F9; B = 16'h00F8; #100;
A = 16'h00F9; B = 16'h00F9; #100;
A = 16'h00F9; B = 16'h00FA; #100;
A = 16'h00F9; B = 16'h00FB; #100;
A = 16'h00F9; B = 16'h00FC; #100;
A = 16'h00F9; B = 16'h00FD; #100;
A = 16'h00F9; B = 16'h00FE; #100;
A = 16'h00F9; B = 16'h00FF; #100;
A = 16'h00FA; B = 16'h000; #100;
A = 16'h00FA; B = 16'h001; #100;
A = 16'h00FA; B = 16'h002; #100;
A = 16'h00FA; B = 16'h003; #100;
A = 16'h00FA; B = 16'h004; #100;
A = 16'h00FA; B = 16'h005; #100;
A = 16'h00FA; B = 16'h006; #100;
A = 16'h00FA; B = 16'h007; #100;
A = 16'h00FA; B = 16'h008; #100;
A = 16'h00FA; B = 16'h009; #100;
A = 16'h00FA; B = 16'h00A; #100;
A = 16'h00FA; B = 16'h00B; #100;
A = 16'h00FA; B = 16'h00C; #100;
A = 16'h00FA; B = 16'h00D; #100;
A = 16'h00FA; B = 16'h00E; #100;
A = 16'h00FA; B = 16'h00F; #100;
A = 16'h00FA; B = 16'h0010; #100;
A = 16'h00FA; B = 16'h0011; #100;
A = 16'h00FA; B = 16'h0012; #100;
A = 16'h00FA; B = 16'h0013; #100;
A = 16'h00FA; B = 16'h0014; #100;
A = 16'h00FA; B = 16'h0015; #100;
A = 16'h00FA; B = 16'h0016; #100;
A = 16'h00FA; B = 16'h0017; #100;
A = 16'h00FA; B = 16'h0018; #100;
A = 16'h00FA; B = 16'h0019; #100;
A = 16'h00FA; B = 16'h001A; #100;
A = 16'h00FA; B = 16'h001B; #100;
A = 16'h00FA; B = 16'h001C; #100;
A = 16'h00FA; B = 16'h001D; #100;
A = 16'h00FA; B = 16'h001E; #100;
A = 16'h00FA; B = 16'h001F; #100;
A = 16'h00FA; B = 16'h0020; #100;
A = 16'h00FA; B = 16'h0021; #100;
A = 16'h00FA; B = 16'h0022; #100;
A = 16'h00FA; B = 16'h0023; #100;
A = 16'h00FA; B = 16'h0024; #100;
A = 16'h00FA; B = 16'h0025; #100;
A = 16'h00FA; B = 16'h0026; #100;
A = 16'h00FA; B = 16'h0027; #100;
A = 16'h00FA; B = 16'h0028; #100;
A = 16'h00FA; B = 16'h0029; #100;
A = 16'h00FA; B = 16'h002A; #100;
A = 16'h00FA; B = 16'h002B; #100;
A = 16'h00FA; B = 16'h002C; #100;
A = 16'h00FA; B = 16'h002D; #100;
A = 16'h00FA; B = 16'h002E; #100;
A = 16'h00FA; B = 16'h002F; #100;
A = 16'h00FA; B = 16'h0030; #100;
A = 16'h00FA; B = 16'h0031; #100;
A = 16'h00FA; B = 16'h0032; #100;
A = 16'h00FA; B = 16'h0033; #100;
A = 16'h00FA; B = 16'h0034; #100;
A = 16'h00FA; B = 16'h0035; #100;
A = 16'h00FA; B = 16'h0036; #100;
A = 16'h00FA; B = 16'h0037; #100;
A = 16'h00FA; B = 16'h0038; #100;
A = 16'h00FA; B = 16'h0039; #100;
A = 16'h00FA; B = 16'h003A; #100;
A = 16'h00FA; B = 16'h003B; #100;
A = 16'h00FA; B = 16'h003C; #100;
A = 16'h00FA; B = 16'h003D; #100;
A = 16'h00FA; B = 16'h003E; #100;
A = 16'h00FA; B = 16'h003F; #100;
A = 16'h00FA; B = 16'h0040; #100;
A = 16'h00FA; B = 16'h0041; #100;
A = 16'h00FA; B = 16'h0042; #100;
A = 16'h00FA; B = 16'h0043; #100;
A = 16'h00FA; B = 16'h0044; #100;
A = 16'h00FA; B = 16'h0045; #100;
A = 16'h00FA; B = 16'h0046; #100;
A = 16'h00FA; B = 16'h0047; #100;
A = 16'h00FA; B = 16'h0048; #100;
A = 16'h00FA; B = 16'h0049; #100;
A = 16'h00FA; B = 16'h004A; #100;
A = 16'h00FA; B = 16'h004B; #100;
A = 16'h00FA; B = 16'h004C; #100;
A = 16'h00FA; B = 16'h004D; #100;
A = 16'h00FA; B = 16'h004E; #100;
A = 16'h00FA; B = 16'h004F; #100;
A = 16'h00FA; B = 16'h0050; #100;
A = 16'h00FA; B = 16'h0051; #100;
A = 16'h00FA; B = 16'h0052; #100;
A = 16'h00FA; B = 16'h0053; #100;
A = 16'h00FA; B = 16'h0054; #100;
A = 16'h00FA; B = 16'h0055; #100;
A = 16'h00FA; B = 16'h0056; #100;
A = 16'h00FA; B = 16'h0057; #100;
A = 16'h00FA; B = 16'h0058; #100;
A = 16'h00FA; B = 16'h0059; #100;
A = 16'h00FA; B = 16'h005A; #100;
A = 16'h00FA; B = 16'h005B; #100;
A = 16'h00FA; B = 16'h005C; #100;
A = 16'h00FA; B = 16'h005D; #100;
A = 16'h00FA; B = 16'h005E; #100;
A = 16'h00FA; B = 16'h005F; #100;
A = 16'h00FA; B = 16'h0060; #100;
A = 16'h00FA; B = 16'h0061; #100;
A = 16'h00FA; B = 16'h0062; #100;
A = 16'h00FA; B = 16'h0063; #100;
A = 16'h00FA; B = 16'h0064; #100;
A = 16'h00FA; B = 16'h0065; #100;
A = 16'h00FA; B = 16'h0066; #100;
A = 16'h00FA; B = 16'h0067; #100;
A = 16'h00FA; B = 16'h0068; #100;
A = 16'h00FA; B = 16'h0069; #100;
A = 16'h00FA; B = 16'h006A; #100;
A = 16'h00FA; B = 16'h006B; #100;
A = 16'h00FA; B = 16'h006C; #100;
A = 16'h00FA; B = 16'h006D; #100;
A = 16'h00FA; B = 16'h006E; #100;
A = 16'h00FA; B = 16'h006F; #100;
A = 16'h00FA; B = 16'h0070; #100;
A = 16'h00FA; B = 16'h0071; #100;
A = 16'h00FA; B = 16'h0072; #100;
A = 16'h00FA; B = 16'h0073; #100;
A = 16'h00FA; B = 16'h0074; #100;
A = 16'h00FA; B = 16'h0075; #100;
A = 16'h00FA; B = 16'h0076; #100;
A = 16'h00FA; B = 16'h0077; #100;
A = 16'h00FA; B = 16'h0078; #100;
A = 16'h00FA; B = 16'h0079; #100;
A = 16'h00FA; B = 16'h007A; #100;
A = 16'h00FA; B = 16'h007B; #100;
A = 16'h00FA; B = 16'h007C; #100;
A = 16'h00FA; B = 16'h007D; #100;
A = 16'h00FA; B = 16'h007E; #100;
A = 16'h00FA; B = 16'h007F; #100;
A = 16'h00FA; B = 16'h0080; #100;
A = 16'h00FA; B = 16'h0081; #100;
A = 16'h00FA; B = 16'h0082; #100;
A = 16'h00FA; B = 16'h0083; #100;
A = 16'h00FA; B = 16'h0084; #100;
A = 16'h00FA; B = 16'h0085; #100;
A = 16'h00FA; B = 16'h0086; #100;
A = 16'h00FA; B = 16'h0087; #100;
A = 16'h00FA; B = 16'h0088; #100;
A = 16'h00FA; B = 16'h0089; #100;
A = 16'h00FA; B = 16'h008A; #100;
A = 16'h00FA; B = 16'h008B; #100;
A = 16'h00FA; B = 16'h008C; #100;
A = 16'h00FA; B = 16'h008D; #100;
A = 16'h00FA; B = 16'h008E; #100;
A = 16'h00FA; B = 16'h008F; #100;
A = 16'h00FA; B = 16'h0090; #100;
A = 16'h00FA; B = 16'h0091; #100;
A = 16'h00FA; B = 16'h0092; #100;
A = 16'h00FA; B = 16'h0093; #100;
A = 16'h00FA; B = 16'h0094; #100;
A = 16'h00FA; B = 16'h0095; #100;
A = 16'h00FA; B = 16'h0096; #100;
A = 16'h00FA; B = 16'h0097; #100;
A = 16'h00FA; B = 16'h0098; #100;
A = 16'h00FA; B = 16'h0099; #100;
A = 16'h00FA; B = 16'h009A; #100;
A = 16'h00FA; B = 16'h009B; #100;
A = 16'h00FA; B = 16'h009C; #100;
A = 16'h00FA; B = 16'h009D; #100;
A = 16'h00FA; B = 16'h009E; #100;
A = 16'h00FA; B = 16'h009F; #100;
A = 16'h00FA; B = 16'h00A0; #100;
A = 16'h00FA; B = 16'h00A1; #100;
A = 16'h00FA; B = 16'h00A2; #100;
A = 16'h00FA; B = 16'h00A3; #100;
A = 16'h00FA; B = 16'h00A4; #100;
A = 16'h00FA; B = 16'h00A5; #100;
A = 16'h00FA; B = 16'h00A6; #100;
A = 16'h00FA; B = 16'h00A7; #100;
A = 16'h00FA; B = 16'h00A8; #100;
A = 16'h00FA; B = 16'h00A9; #100;
A = 16'h00FA; B = 16'h00AA; #100;
A = 16'h00FA; B = 16'h00AB; #100;
A = 16'h00FA; B = 16'h00AC; #100;
A = 16'h00FA; B = 16'h00AD; #100;
A = 16'h00FA; B = 16'h00AE; #100;
A = 16'h00FA; B = 16'h00AF; #100;
A = 16'h00FA; B = 16'h00B0; #100;
A = 16'h00FA; B = 16'h00B1; #100;
A = 16'h00FA; B = 16'h00B2; #100;
A = 16'h00FA; B = 16'h00B3; #100;
A = 16'h00FA; B = 16'h00B4; #100;
A = 16'h00FA; B = 16'h00B5; #100;
A = 16'h00FA; B = 16'h00B6; #100;
A = 16'h00FA; B = 16'h00B7; #100;
A = 16'h00FA; B = 16'h00B8; #100;
A = 16'h00FA; B = 16'h00B9; #100;
A = 16'h00FA; B = 16'h00BA; #100;
A = 16'h00FA; B = 16'h00BB; #100;
A = 16'h00FA; B = 16'h00BC; #100;
A = 16'h00FA; B = 16'h00BD; #100;
A = 16'h00FA; B = 16'h00BE; #100;
A = 16'h00FA; B = 16'h00BF; #100;
A = 16'h00FA; B = 16'h00C0; #100;
A = 16'h00FA; B = 16'h00C1; #100;
A = 16'h00FA; B = 16'h00C2; #100;
A = 16'h00FA; B = 16'h00C3; #100;
A = 16'h00FA; B = 16'h00C4; #100;
A = 16'h00FA; B = 16'h00C5; #100;
A = 16'h00FA; B = 16'h00C6; #100;
A = 16'h00FA; B = 16'h00C7; #100;
A = 16'h00FA; B = 16'h00C8; #100;
A = 16'h00FA; B = 16'h00C9; #100;
A = 16'h00FA; B = 16'h00CA; #100;
A = 16'h00FA; B = 16'h00CB; #100;
A = 16'h00FA; B = 16'h00CC; #100;
A = 16'h00FA; B = 16'h00CD; #100;
A = 16'h00FA; B = 16'h00CE; #100;
A = 16'h00FA; B = 16'h00CF; #100;
A = 16'h00FA; B = 16'h00D0; #100;
A = 16'h00FA; B = 16'h00D1; #100;
A = 16'h00FA; B = 16'h00D2; #100;
A = 16'h00FA; B = 16'h00D3; #100;
A = 16'h00FA; B = 16'h00D4; #100;
A = 16'h00FA; B = 16'h00D5; #100;
A = 16'h00FA; B = 16'h00D6; #100;
A = 16'h00FA; B = 16'h00D7; #100;
A = 16'h00FA; B = 16'h00D8; #100;
A = 16'h00FA; B = 16'h00D9; #100;
A = 16'h00FA; B = 16'h00DA; #100;
A = 16'h00FA; B = 16'h00DB; #100;
A = 16'h00FA; B = 16'h00DC; #100;
A = 16'h00FA; B = 16'h00DD; #100;
A = 16'h00FA; B = 16'h00DE; #100;
A = 16'h00FA; B = 16'h00DF; #100;
A = 16'h00FA; B = 16'h00E0; #100;
A = 16'h00FA; B = 16'h00E1; #100;
A = 16'h00FA; B = 16'h00E2; #100;
A = 16'h00FA; B = 16'h00E3; #100;
A = 16'h00FA; B = 16'h00E4; #100;
A = 16'h00FA; B = 16'h00E5; #100;
A = 16'h00FA; B = 16'h00E6; #100;
A = 16'h00FA; B = 16'h00E7; #100;
A = 16'h00FA; B = 16'h00E8; #100;
A = 16'h00FA; B = 16'h00E9; #100;
A = 16'h00FA; B = 16'h00EA; #100;
A = 16'h00FA; B = 16'h00EB; #100;
A = 16'h00FA; B = 16'h00EC; #100;
A = 16'h00FA; B = 16'h00ED; #100;
A = 16'h00FA; B = 16'h00EE; #100;
A = 16'h00FA; B = 16'h00EF; #100;
A = 16'h00FA; B = 16'h00F0; #100;
A = 16'h00FA; B = 16'h00F1; #100;
A = 16'h00FA; B = 16'h00F2; #100;
A = 16'h00FA; B = 16'h00F3; #100;
A = 16'h00FA; B = 16'h00F4; #100;
A = 16'h00FA; B = 16'h00F5; #100;
A = 16'h00FA; B = 16'h00F6; #100;
A = 16'h00FA; B = 16'h00F7; #100;
A = 16'h00FA; B = 16'h00F8; #100;
A = 16'h00FA; B = 16'h00F9; #100;
A = 16'h00FA; B = 16'h00FA; #100;
A = 16'h00FA; B = 16'h00FB; #100;
A = 16'h00FA; B = 16'h00FC; #100;
A = 16'h00FA; B = 16'h00FD; #100;
A = 16'h00FA; B = 16'h00FE; #100;
A = 16'h00FA; B = 16'h00FF; #100;
A = 16'h00FB; B = 16'h000; #100;
A = 16'h00FB; B = 16'h001; #100;
A = 16'h00FB; B = 16'h002; #100;
A = 16'h00FB; B = 16'h003; #100;
A = 16'h00FB; B = 16'h004; #100;
A = 16'h00FB; B = 16'h005; #100;
A = 16'h00FB; B = 16'h006; #100;
A = 16'h00FB; B = 16'h007; #100;
A = 16'h00FB; B = 16'h008; #100;
A = 16'h00FB; B = 16'h009; #100;
A = 16'h00FB; B = 16'h00A; #100;
A = 16'h00FB; B = 16'h00B; #100;
A = 16'h00FB; B = 16'h00C; #100;
A = 16'h00FB; B = 16'h00D; #100;
A = 16'h00FB; B = 16'h00E; #100;
A = 16'h00FB; B = 16'h00F; #100;
A = 16'h00FB; B = 16'h0010; #100;
A = 16'h00FB; B = 16'h0011; #100;
A = 16'h00FB; B = 16'h0012; #100;
A = 16'h00FB; B = 16'h0013; #100;
A = 16'h00FB; B = 16'h0014; #100;
A = 16'h00FB; B = 16'h0015; #100;
A = 16'h00FB; B = 16'h0016; #100;
A = 16'h00FB; B = 16'h0017; #100;
A = 16'h00FB; B = 16'h0018; #100;
A = 16'h00FB; B = 16'h0019; #100;
A = 16'h00FB; B = 16'h001A; #100;
A = 16'h00FB; B = 16'h001B; #100;
A = 16'h00FB; B = 16'h001C; #100;
A = 16'h00FB; B = 16'h001D; #100;
A = 16'h00FB; B = 16'h001E; #100;
A = 16'h00FB; B = 16'h001F; #100;
A = 16'h00FB; B = 16'h0020; #100;
A = 16'h00FB; B = 16'h0021; #100;
A = 16'h00FB; B = 16'h0022; #100;
A = 16'h00FB; B = 16'h0023; #100;
A = 16'h00FB; B = 16'h0024; #100;
A = 16'h00FB; B = 16'h0025; #100;
A = 16'h00FB; B = 16'h0026; #100;
A = 16'h00FB; B = 16'h0027; #100;
A = 16'h00FB; B = 16'h0028; #100;
A = 16'h00FB; B = 16'h0029; #100;
A = 16'h00FB; B = 16'h002A; #100;
A = 16'h00FB; B = 16'h002B; #100;
A = 16'h00FB; B = 16'h002C; #100;
A = 16'h00FB; B = 16'h002D; #100;
A = 16'h00FB; B = 16'h002E; #100;
A = 16'h00FB; B = 16'h002F; #100;
A = 16'h00FB; B = 16'h0030; #100;
A = 16'h00FB; B = 16'h0031; #100;
A = 16'h00FB; B = 16'h0032; #100;
A = 16'h00FB; B = 16'h0033; #100;
A = 16'h00FB; B = 16'h0034; #100;
A = 16'h00FB; B = 16'h0035; #100;
A = 16'h00FB; B = 16'h0036; #100;
A = 16'h00FB; B = 16'h0037; #100;
A = 16'h00FB; B = 16'h0038; #100;
A = 16'h00FB; B = 16'h0039; #100;
A = 16'h00FB; B = 16'h003A; #100;
A = 16'h00FB; B = 16'h003B; #100;
A = 16'h00FB; B = 16'h003C; #100;
A = 16'h00FB; B = 16'h003D; #100;
A = 16'h00FB; B = 16'h003E; #100;
A = 16'h00FB; B = 16'h003F; #100;
A = 16'h00FB; B = 16'h0040; #100;
A = 16'h00FB; B = 16'h0041; #100;
A = 16'h00FB; B = 16'h0042; #100;
A = 16'h00FB; B = 16'h0043; #100;
A = 16'h00FB; B = 16'h0044; #100;
A = 16'h00FB; B = 16'h0045; #100;
A = 16'h00FB; B = 16'h0046; #100;
A = 16'h00FB; B = 16'h0047; #100;
A = 16'h00FB; B = 16'h0048; #100;
A = 16'h00FB; B = 16'h0049; #100;
A = 16'h00FB; B = 16'h004A; #100;
A = 16'h00FB; B = 16'h004B; #100;
A = 16'h00FB; B = 16'h004C; #100;
A = 16'h00FB; B = 16'h004D; #100;
A = 16'h00FB; B = 16'h004E; #100;
A = 16'h00FB; B = 16'h004F; #100;
A = 16'h00FB; B = 16'h0050; #100;
A = 16'h00FB; B = 16'h0051; #100;
A = 16'h00FB; B = 16'h0052; #100;
A = 16'h00FB; B = 16'h0053; #100;
A = 16'h00FB; B = 16'h0054; #100;
A = 16'h00FB; B = 16'h0055; #100;
A = 16'h00FB; B = 16'h0056; #100;
A = 16'h00FB; B = 16'h0057; #100;
A = 16'h00FB; B = 16'h0058; #100;
A = 16'h00FB; B = 16'h0059; #100;
A = 16'h00FB; B = 16'h005A; #100;
A = 16'h00FB; B = 16'h005B; #100;
A = 16'h00FB; B = 16'h005C; #100;
A = 16'h00FB; B = 16'h005D; #100;
A = 16'h00FB; B = 16'h005E; #100;
A = 16'h00FB; B = 16'h005F; #100;
A = 16'h00FB; B = 16'h0060; #100;
A = 16'h00FB; B = 16'h0061; #100;
A = 16'h00FB; B = 16'h0062; #100;
A = 16'h00FB; B = 16'h0063; #100;
A = 16'h00FB; B = 16'h0064; #100;
A = 16'h00FB; B = 16'h0065; #100;
A = 16'h00FB; B = 16'h0066; #100;
A = 16'h00FB; B = 16'h0067; #100;
A = 16'h00FB; B = 16'h0068; #100;
A = 16'h00FB; B = 16'h0069; #100;
A = 16'h00FB; B = 16'h006A; #100;
A = 16'h00FB; B = 16'h006B; #100;
A = 16'h00FB; B = 16'h006C; #100;
A = 16'h00FB; B = 16'h006D; #100;
A = 16'h00FB; B = 16'h006E; #100;
A = 16'h00FB; B = 16'h006F; #100;
A = 16'h00FB; B = 16'h0070; #100;
A = 16'h00FB; B = 16'h0071; #100;
A = 16'h00FB; B = 16'h0072; #100;
A = 16'h00FB; B = 16'h0073; #100;
A = 16'h00FB; B = 16'h0074; #100;
A = 16'h00FB; B = 16'h0075; #100;
A = 16'h00FB; B = 16'h0076; #100;
A = 16'h00FB; B = 16'h0077; #100;
A = 16'h00FB; B = 16'h0078; #100;
A = 16'h00FB; B = 16'h0079; #100;
A = 16'h00FB; B = 16'h007A; #100;
A = 16'h00FB; B = 16'h007B; #100;
A = 16'h00FB; B = 16'h007C; #100;
A = 16'h00FB; B = 16'h007D; #100;
A = 16'h00FB; B = 16'h007E; #100;
A = 16'h00FB; B = 16'h007F; #100;
A = 16'h00FB; B = 16'h0080; #100;
A = 16'h00FB; B = 16'h0081; #100;
A = 16'h00FB; B = 16'h0082; #100;
A = 16'h00FB; B = 16'h0083; #100;
A = 16'h00FB; B = 16'h0084; #100;
A = 16'h00FB; B = 16'h0085; #100;
A = 16'h00FB; B = 16'h0086; #100;
A = 16'h00FB; B = 16'h0087; #100;
A = 16'h00FB; B = 16'h0088; #100;
A = 16'h00FB; B = 16'h0089; #100;
A = 16'h00FB; B = 16'h008A; #100;
A = 16'h00FB; B = 16'h008B; #100;
A = 16'h00FB; B = 16'h008C; #100;
A = 16'h00FB; B = 16'h008D; #100;
A = 16'h00FB; B = 16'h008E; #100;
A = 16'h00FB; B = 16'h008F; #100;
A = 16'h00FB; B = 16'h0090; #100;
A = 16'h00FB; B = 16'h0091; #100;
A = 16'h00FB; B = 16'h0092; #100;
A = 16'h00FB; B = 16'h0093; #100;
A = 16'h00FB; B = 16'h0094; #100;
A = 16'h00FB; B = 16'h0095; #100;
A = 16'h00FB; B = 16'h0096; #100;
A = 16'h00FB; B = 16'h0097; #100;
A = 16'h00FB; B = 16'h0098; #100;
A = 16'h00FB; B = 16'h0099; #100;
A = 16'h00FB; B = 16'h009A; #100;
A = 16'h00FB; B = 16'h009B; #100;
A = 16'h00FB; B = 16'h009C; #100;
A = 16'h00FB; B = 16'h009D; #100;
A = 16'h00FB; B = 16'h009E; #100;
A = 16'h00FB; B = 16'h009F; #100;
A = 16'h00FB; B = 16'h00A0; #100;
A = 16'h00FB; B = 16'h00A1; #100;
A = 16'h00FB; B = 16'h00A2; #100;
A = 16'h00FB; B = 16'h00A3; #100;
A = 16'h00FB; B = 16'h00A4; #100;
A = 16'h00FB; B = 16'h00A5; #100;
A = 16'h00FB; B = 16'h00A6; #100;
A = 16'h00FB; B = 16'h00A7; #100;
A = 16'h00FB; B = 16'h00A8; #100;
A = 16'h00FB; B = 16'h00A9; #100;
A = 16'h00FB; B = 16'h00AA; #100;
A = 16'h00FB; B = 16'h00AB; #100;
A = 16'h00FB; B = 16'h00AC; #100;
A = 16'h00FB; B = 16'h00AD; #100;
A = 16'h00FB; B = 16'h00AE; #100;
A = 16'h00FB; B = 16'h00AF; #100;
A = 16'h00FB; B = 16'h00B0; #100;
A = 16'h00FB; B = 16'h00B1; #100;
A = 16'h00FB; B = 16'h00B2; #100;
A = 16'h00FB; B = 16'h00B3; #100;
A = 16'h00FB; B = 16'h00B4; #100;
A = 16'h00FB; B = 16'h00B5; #100;
A = 16'h00FB; B = 16'h00B6; #100;
A = 16'h00FB; B = 16'h00B7; #100;
A = 16'h00FB; B = 16'h00B8; #100;
A = 16'h00FB; B = 16'h00B9; #100;
A = 16'h00FB; B = 16'h00BA; #100;
A = 16'h00FB; B = 16'h00BB; #100;
A = 16'h00FB; B = 16'h00BC; #100;
A = 16'h00FB; B = 16'h00BD; #100;
A = 16'h00FB; B = 16'h00BE; #100;
A = 16'h00FB; B = 16'h00BF; #100;
A = 16'h00FB; B = 16'h00C0; #100;
A = 16'h00FB; B = 16'h00C1; #100;
A = 16'h00FB; B = 16'h00C2; #100;
A = 16'h00FB; B = 16'h00C3; #100;
A = 16'h00FB; B = 16'h00C4; #100;
A = 16'h00FB; B = 16'h00C5; #100;
A = 16'h00FB; B = 16'h00C6; #100;
A = 16'h00FB; B = 16'h00C7; #100;
A = 16'h00FB; B = 16'h00C8; #100;
A = 16'h00FB; B = 16'h00C9; #100;
A = 16'h00FB; B = 16'h00CA; #100;
A = 16'h00FB; B = 16'h00CB; #100;
A = 16'h00FB; B = 16'h00CC; #100;
A = 16'h00FB; B = 16'h00CD; #100;
A = 16'h00FB; B = 16'h00CE; #100;
A = 16'h00FB; B = 16'h00CF; #100;
A = 16'h00FB; B = 16'h00D0; #100;
A = 16'h00FB; B = 16'h00D1; #100;
A = 16'h00FB; B = 16'h00D2; #100;
A = 16'h00FB; B = 16'h00D3; #100;
A = 16'h00FB; B = 16'h00D4; #100;
A = 16'h00FB; B = 16'h00D5; #100;
A = 16'h00FB; B = 16'h00D6; #100;
A = 16'h00FB; B = 16'h00D7; #100;
A = 16'h00FB; B = 16'h00D8; #100;
A = 16'h00FB; B = 16'h00D9; #100;
A = 16'h00FB; B = 16'h00DA; #100;
A = 16'h00FB; B = 16'h00DB; #100;
A = 16'h00FB; B = 16'h00DC; #100;
A = 16'h00FB; B = 16'h00DD; #100;
A = 16'h00FB; B = 16'h00DE; #100;
A = 16'h00FB; B = 16'h00DF; #100;
A = 16'h00FB; B = 16'h00E0; #100;
A = 16'h00FB; B = 16'h00E1; #100;
A = 16'h00FB; B = 16'h00E2; #100;
A = 16'h00FB; B = 16'h00E3; #100;
A = 16'h00FB; B = 16'h00E4; #100;
A = 16'h00FB; B = 16'h00E5; #100;
A = 16'h00FB; B = 16'h00E6; #100;
A = 16'h00FB; B = 16'h00E7; #100;
A = 16'h00FB; B = 16'h00E8; #100;
A = 16'h00FB; B = 16'h00E9; #100;
A = 16'h00FB; B = 16'h00EA; #100;
A = 16'h00FB; B = 16'h00EB; #100;
A = 16'h00FB; B = 16'h00EC; #100;
A = 16'h00FB; B = 16'h00ED; #100;
A = 16'h00FB; B = 16'h00EE; #100;
A = 16'h00FB; B = 16'h00EF; #100;
A = 16'h00FB; B = 16'h00F0; #100;
A = 16'h00FB; B = 16'h00F1; #100;
A = 16'h00FB; B = 16'h00F2; #100;
A = 16'h00FB; B = 16'h00F3; #100;
A = 16'h00FB; B = 16'h00F4; #100;
A = 16'h00FB; B = 16'h00F5; #100;
A = 16'h00FB; B = 16'h00F6; #100;
A = 16'h00FB; B = 16'h00F7; #100;
A = 16'h00FB; B = 16'h00F8; #100;
A = 16'h00FB; B = 16'h00F9; #100;
A = 16'h00FB; B = 16'h00FA; #100;
A = 16'h00FB; B = 16'h00FB; #100;
A = 16'h00FB; B = 16'h00FC; #100;
A = 16'h00FB; B = 16'h00FD; #100;
A = 16'h00FB; B = 16'h00FE; #100;
A = 16'h00FB; B = 16'h00FF; #100;
A = 16'h00FC; B = 16'h000; #100;
A = 16'h00FC; B = 16'h001; #100;
A = 16'h00FC; B = 16'h002; #100;
A = 16'h00FC; B = 16'h003; #100;
A = 16'h00FC; B = 16'h004; #100;
A = 16'h00FC; B = 16'h005; #100;
A = 16'h00FC; B = 16'h006; #100;
A = 16'h00FC; B = 16'h007; #100;
A = 16'h00FC; B = 16'h008; #100;
A = 16'h00FC; B = 16'h009; #100;
A = 16'h00FC; B = 16'h00A; #100;
A = 16'h00FC; B = 16'h00B; #100;
A = 16'h00FC; B = 16'h00C; #100;
A = 16'h00FC; B = 16'h00D; #100;
A = 16'h00FC; B = 16'h00E; #100;
A = 16'h00FC; B = 16'h00F; #100;
A = 16'h00FC; B = 16'h0010; #100;
A = 16'h00FC; B = 16'h0011; #100;
A = 16'h00FC; B = 16'h0012; #100;
A = 16'h00FC; B = 16'h0013; #100;
A = 16'h00FC; B = 16'h0014; #100;
A = 16'h00FC; B = 16'h0015; #100;
A = 16'h00FC; B = 16'h0016; #100;
A = 16'h00FC; B = 16'h0017; #100;
A = 16'h00FC; B = 16'h0018; #100;
A = 16'h00FC; B = 16'h0019; #100;
A = 16'h00FC; B = 16'h001A; #100;
A = 16'h00FC; B = 16'h001B; #100;
A = 16'h00FC; B = 16'h001C; #100;
A = 16'h00FC; B = 16'h001D; #100;
A = 16'h00FC; B = 16'h001E; #100;
A = 16'h00FC; B = 16'h001F; #100;
A = 16'h00FC; B = 16'h0020; #100;
A = 16'h00FC; B = 16'h0021; #100;
A = 16'h00FC; B = 16'h0022; #100;
A = 16'h00FC; B = 16'h0023; #100;
A = 16'h00FC; B = 16'h0024; #100;
A = 16'h00FC; B = 16'h0025; #100;
A = 16'h00FC; B = 16'h0026; #100;
A = 16'h00FC; B = 16'h0027; #100;
A = 16'h00FC; B = 16'h0028; #100;
A = 16'h00FC; B = 16'h0029; #100;
A = 16'h00FC; B = 16'h002A; #100;
A = 16'h00FC; B = 16'h002B; #100;
A = 16'h00FC; B = 16'h002C; #100;
A = 16'h00FC; B = 16'h002D; #100;
A = 16'h00FC; B = 16'h002E; #100;
A = 16'h00FC; B = 16'h002F; #100;
A = 16'h00FC; B = 16'h0030; #100;
A = 16'h00FC; B = 16'h0031; #100;
A = 16'h00FC; B = 16'h0032; #100;
A = 16'h00FC; B = 16'h0033; #100;
A = 16'h00FC; B = 16'h0034; #100;
A = 16'h00FC; B = 16'h0035; #100;
A = 16'h00FC; B = 16'h0036; #100;
A = 16'h00FC; B = 16'h0037; #100;
A = 16'h00FC; B = 16'h0038; #100;
A = 16'h00FC; B = 16'h0039; #100;
A = 16'h00FC; B = 16'h003A; #100;
A = 16'h00FC; B = 16'h003B; #100;
A = 16'h00FC; B = 16'h003C; #100;
A = 16'h00FC; B = 16'h003D; #100;
A = 16'h00FC; B = 16'h003E; #100;
A = 16'h00FC; B = 16'h003F; #100;
A = 16'h00FC; B = 16'h0040; #100;
A = 16'h00FC; B = 16'h0041; #100;
A = 16'h00FC; B = 16'h0042; #100;
A = 16'h00FC; B = 16'h0043; #100;
A = 16'h00FC; B = 16'h0044; #100;
A = 16'h00FC; B = 16'h0045; #100;
A = 16'h00FC; B = 16'h0046; #100;
A = 16'h00FC; B = 16'h0047; #100;
A = 16'h00FC; B = 16'h0048; #100;
A = 16'h00FC; B = 16'h0049; #100;
A = 16'h00FC; B = 16'h004A; #100;
A = 16'h00FC; B = 16'h004B; #100;
A = 16'h00FC; B = 16'h004C; #100;
A = 16'h00FC; B = 16'h004D; #100;
A = 16'h00FC; B = 16'h004E; #100;
A = 16'h00FC; B = 16'h004F; #100;
A = 16'h00FC; B = 16'h0050; #100;
A = 16'h00FC; B = 16'h0051; #100;
A = 16'h00FC; B = 16'h0052; #100;
A = 16'h00FC; B = 16'h0053; #100;
A = 16'h00FC; B = 16'h0054; #100;
A = 16'h00FC; B = 16'h0055; #100;
A = 16'h00FC; B = 16'h0056; #100;
A = 16'h00FC; B = 16'h0057; #100;
A = 16'h00FC; B = 16'h0058; #100;
A = 16'h00FC; B = 16'h0059; #100;
A = 16'h00FC; B = 16'h005A; #100;
A = 16'h00FC; B = 16'h005B; #100;
A = 16'h00FC; B = 16'h005C; #100;
A = 16'h00FC; B = 16'h005D; #100;
A = 16'h00FC; B = 16'h005E; #100;
A = 16'h00FC; B = 16'h005F; #100;
A = 16'h00FC; B = 16'h0060; #100;
A = 16'h00FC; B = 16'h0061; #100;
A = 16'h00FC; B = 16'h0062; #100;
A = 16'h00FC; B = 16'h0063; #100;
A = 16'h00FC; B = 16'h0064; #100;
A = 16'h00FC; B = 16'h0065; #100;
A = 16'h00FC; B = 16'h0066; #100;
A = 16'h00FC; B = 16'h0067; #100;
A = 16'h00FC; B = 16'h0068; #100;
A = 16'h00FC; B = 16'h0069; #100;
A = 16'h00FC; B = 16'h006A; #100;
A = 16'h00FC; B = 16'h006B; #100;
A = 16'h00FC; B = 16'h006C; #100;
A = 16'h00FC; B = 16'h006D; #100;
A = 16'h00FC; B = 16'h006E; #100;
A = 16'h00FC; B = 16'h006F; #100;
A = 16'h00FC; B = 16'h0070; #100;
A = 16'h00FC; B = 16'h0071; #100;
A = 16'h00FC; B = 16'h0072; #100;
A = 16'h00FC; B = 16'h0073; #100;
A = 16'h00FC; B = 16'h0074; #100;
A = 16'h00FC; B = 16'h0075; #100;
A = 16'h00FC; B = 16'h0076; #100;
A = 16'h00FC; B = 16'h0077; #100;
A = 16'h00FC; B = 16'h0078; #100;
A = 16'h00FC; B = 16'h0079; #100;
A = 16'h00FC; B = 16'h007A; #100;
A = 16'h00FC; B = 16'h007B; #100;
A = 16'h00FC; B = 16'h007C; #100;
A = 16'h00FC; B = 16'h007D; #100;
A = 16'h00FC; B = 16'h007E; #100;
A = 16'h00FC; B = 16'h007F; #100;
A = 16'h00FC; B = 16'h0080; #100;
A = 16'h00FC; B = 16'h0081; #100;
A = 16'h00FC; B = 16'h0082; #100;
A = 16'h00FC; B = 16'h0083; #100;
A = 16'h00FC; B = 16'h0084; #100;
A = 16'h00FC; B = 16'h0085; #100;
A = 16'h00FC; B = 16'h0086; #100;
A = 16'h00FC; B = 16'h0087; #100;
A = 16'h00FC; B = 16'h0088; #100;
A = 16'h00FC; B = 16'h0089; #100;
A = 16'h00FC; B = 16'h008A; #100;
A = 16'h00FC; B = 16'h008B; #100;
A = 16'h00FC; B = 16'h008C; #100;
A = 16'h00FC; B = 16'h008D; #100;
A = 16'h00FC; B = 16'h008E; #100;
A = 16'h00FC; B = 16'h008F; #100;
A = 16'h00FC; B = 16'h0090; #100;
A = 16'h00FC; B = 16'h0091; #100;
A = 16'h00FC; B = 16'h0092; #100;
A = 16'h00FC; B = 16'h0093; #100;
A = 16'h00FC; B = 16'h0094; #100;
A = 16'h00FC; B = 16'h0095; #100;
A = 16'h00FC; B = 16'h0096; #100;
A = 16'h00FC; B = 16'h0097; #100;
A = 16'h00FC; B = 16'h0098; #100;
A = 16'h00FC; B = 16'h0099; #100;
A = 16'h00FC; B = 16'h009A; #100;
A = 16'h00FC; B = 16'h009B; #100;
A = 16'h00FC; B = 16'h009C; #100;
A = 16'h00FC; B = 16'h009D; #100;
A = 16'h00FC; B = 16'h009E; #100;
A = 16'h00FC; B = 16'h009F; #100;
A = 16'h00FC; B = 16'h00A0; #100;
A = 16'h00FC; B = 16'h00A1; #100;
A = 16'h00FC; B = 16'h00A2; #100;
A = 16'h00FC; B = 16'h00A3; #100;
A = 16'h00FC; B = 16'h00A4; #100;
A = 16'h00FC; B = 16'h00A5; #100;
A = 16'h00FC; B = 16'h00A6; #100;
A = 16'h00FC; B = 16'h00A7; #100;
A = 16'h00FC; B = 16'h00A8; #100;
A = 16'h00FC; B = 16'h00A9; #100;
A = 16'h00FC; B = 16'h00AA; #100;
A = 16'h00FC; B = 16'h00AB; #100;
A = 16'h00FC; B = 16'h00AC; #100;
A = 16'h00FC; B = 16'h00AD; #100;
A = 16'h00FC; B = 16'h00AE; #100;
A = 16'h00FC; B = 16'h00AF; #100;
A = 16'h00FC; B = 16'h00B0; #100;
A = 16'h00FC; B = 16'h00B1; #100;
A = 16'h00FC; B = 16'h00B2; #100;
A = 16'h00FC; B = 16'h00B3; #100;
A = 16'h00FC; B = 16'h00B4; #100;
A = 16'h00FC; B = 16'h00B5; #100;
A = 16'h00FC; B = 16'h00B6; #100;
A = 16'h00FC; B = 16'h00B7; #100;
A = 16'h00FC; B = 16'h00B8; #100;
A = 16'h00FC; B = 16'h00B9; #100;
A = 16'h00FC; B = 16'h00BA; #100;
A = 16'h00FC; B = 16'h00BB; #100;
A = 16'h00FC; B = 16'h00BC; #100;
A = 16'h00FC; B = 16'h00BD; #100;
A = 16'h00FC; B = 16'h00BE; #100;
A = 16'h00FC; B = 16'h00BF; #100;
A = 16'h00FC; B = 16'h00C0; #100;
A = 16'h00FC; B = 16'h00C1; #100;
A = 16'h00FC; B = 16'h00C2; #100;
A = 16'h00FC; B = 16'h00C3; #100;
A = 16'h00FC; B = 16'h00C4; #100;
A = 16'h00FC; B = 16'h00C5; #100;
A = 16'h00FC; B = 16'h00C6; #100;
A = 16'h00FC; B = 16'h00C7; #100;
A = 16'h00FC; B = 16'h00C8; #100;
A = 16'h00FC; B = 16'h00C9; #100;
A = 16'h00FC; B = 16'h00CA; #100;
A = 16'h00FC; B = 16'h00CB; #100;
A = 16'h00FC; B = 16'h00CC; #100;
A = 16'h00FC; B = 16'h00CD; #100;
A = 16'h00FC; B = 16'h00CE; #100;
A = 16'h00FC; B = 16'h00CF; #100;
A = 16'h00FC; B = 16'h00D0; #100;
A = 16'h00FC; B = 16'h00D1; #100;
A = 16'h00FC; B = 16'h00D2; #100;
A = 16'h00FC; B = 16'h00D3; #100;
A = 16'h00FC; B = 16'h00D4; #100;
A = 16'h00FC; B = 16'h00D5; #100;
A = 16'h00FC; B = 16'h00D6; #100;
A = 16'h00FC; B = 16'h00D7; #100;
A = 16'h00FC; B = 16'h00D8; #100;
A = 16'h00FC; B = 16'h00D9; #100;
A = 16'h00FC; B = 16'h00DA; #100;
A = 16'h00FC; B = 16'h00DB; #100;
A = 16'h00FC; B = 16'h00DC; #100;
A = 16'h00FC; B = 16'h00DD; #100;
A = 16'h00FC; B = 16'h00DE; #100;
A = 16'h00FC; B = 16'h00DF; #100;
A = 16'h00FC; B = 16'h00E0; #100;
A = 16'h00FC; B = 16'h00E1; #100;
A = 16'h00FC; B = 16'h00E2; #100;
A = 16'h00FC; B = 16'h00E3; #100;
A = 16'h00FC; B = 16'h00E4; #100;
A = 16'h00FC; B = 16'h00E5; #100;
A = 16'h00FC; B = 16'h00E6; #100;
A = 16'h00FC; B = 16'h00E7; #100;
A = 16'h00FC; B = 16'h00E8; #100;
A = 16'h00FC; B = 16'h00E9; #100;
A = 16'h00FC; B = 16'h00EA; #100;
A = 16'h00FC; B = 16'h00EB; #100;
A = 16'h00FC; B = 16'h00EC; #100;
A = 16'h00FC; B = 16'h00ED; #100;
A = 16'h00FC; B = 16'h00EE; #100;
A = 16'h00FC; B = 16'h00EF; #100;
A = 16'h00FC; B = 16'h00F0; #100;
A = 16'h00FC; B = 16'h00F1; #100;
A = 16'h00FC; B = 16'h00F2; #100;
A = 16'h00FC; B = 16'h00F3; #100;
A = 16'h00FC; B = 16'h00F4; #100;
A = 16'h00FC; B = 16'h00F5; #100;
A = 16'h00FC; B = 16'h00F6; #100;
A = 16'h00FC; B = 16'h00F7; #100;
A = 16'h00FC; B = 16'h00F8; #100;
A = 16'h00FC; B = 16'h00F9; #100;
A = 16'h00FC; B = 16'h00FA; #100;
A = 16'h00FC; B = 16'h00FB; #100;
A = 16'h00FC; B = 16'h00FC; #100;
A = 16'h00FC; B = 16'h00FD; #100;
A = 16'h00FC; B = 16'h00FE; #100;
A = 16'h00FC; B = 16'h00FF; #100;
A = 16'h00FD; B = 16'h000; #100;
A = 16'h00FD; B = 16'h001; #100;
A = 16'h00FD; B = 16'h002; #100;
A = 16'h00FD; B = 16'h003; #100;
A = 16'h00FD; B = 16'h004; #100;
A = 16'h00FD; B = 16'h005; #100;
A = 16'h00FD; B = 16'h006; #100;
A = 16'h00FD; B = 16'h007; #100;
A = 16'h00FD; B = 16'h008; #100;
A = 16'h00FD; B = 16'h009; #100;
A = 16'h00FD; B = 16'h00A; #100;
A = 16'h00FD; B = 16'h00B; #100;
A = 16'h00FD; B = 16'h00C; #100;
A = 16'h00FD; B = 16'h00D; #100;
A = 16'h00FD; B = 16'h00E; #100;
A = 16'h00FD; B = 16'h00F; #100;
A = 16'h00FD; B = 16'h0010; #100;
A = 16'h00FD; B = 16'h0011; #100;
A = 16'h00FD; B = 16'h0012; #100;
A = 16'h00FD; B = 16'h0013; #100;
A = 16'h00FD; B = 16'h0014; #100;
A = 16'h00FD; B = 16'h0015; #100;
A = 16'h00FD; B = 16'h0016; #100;
A = 16'h00FD; B = 16'h0017; #100;
A = 16'h00FD; B = 16'h0018; #100;
A = 16'h00FD; B = 16'h0019; #100;
A = 16'h00FD; B = 16'h001A; #100;
A = 16'h00FD; B = 16'h001B; #100;
A = 16'h00FD; B = 16'h001C; #100;
A = 16'h00FD; B = 16'h001D; #100;
A = 16'h00FD; B = 16'h001E; #100;
A = 16'h00FD; B = 16'h001F; #100;
A = 16'h00FD; B = 16'h0020; #100;
A = 16'h00FD; B = 16'h0021; #100;
A = 16'h00FD; B = 16'h0022; #100;
A = 16'h00FD; B = 16'h0023; #100;
A = 16'h00FD; B = 16'h0024; #100;
A = 16'h00FD; B = 16'h0025; #100;
A = 16'h00FD; B = 16'h0026; #100;
A = 16'h00FD; B = 16'h0027; #100;
A = 16'h00FD; B = 16'h0028; #100;
A = 16'h00FD; B = 16'h0029; #100;
A = 16'h00FD; B = 16'h002A; #100;
A = 16'h00FD; B = 16'h002B; #100;
A = 16'h00FD; B = 16'h002C; #100;
A = 16'h00FD; B = 16'h002D; #100;
A = 16'h00FD; B = 16'h002E; #100;
A = 16'h00FD; B = 16'h002F; #100;
A = 16'h00FD; B = 16'h0030; #100;
A = 16'h00FD; B = 16'h0031; #100;
A = 16'h00FD; B = 16'h0032; #100;
A = 16'h00FD; B = 16'h0033; #100;
A = 16'h00FD; B = 16'h0034; #100;
A = 16'h00FD; B = 16'h0035; #100;
A = 16'h00FD; B = 16'h0036; #100;
A = 16'h00FD; B = 16'h0037; #100;
A = 16'h00FD; B = 16'h0038; #100;
A = 16'h00FD; B = 16'h0039; #100;
A = 16'h00FD; B = 16'h003A; #100;
A = 16'h00FD; B = 16'h003B; #100;
A = 16'h00FD; B = 16'h003C; #100;
A = 16'h00FD; B = 16'h003D; #100;
A = 16'h00FD; B = 16'h003E; #100;
A = 16'h00FD; B = 16'h003F; #100;
A = 16'h00FD; B = 16'h0040; #100;
A = 16'h00FD; B = 16'h0041; #100;
A = 16'h00FD; B = 16'h0042; #100;
A = 16'h00FD; B = 16'h0043; #100;
A = 16'h00FD; B = 16'h0044; #100;
A = 16'h00FD; B = 16'h0045; #100;
A = 16'h00FD; B = 16'h0046; #100;
A = 16'h00FD; B = 16'h0047; #100;
A = 16'h00FD; B = 16'h0048; #100;
A = 16'h00FD; B = 16'h0049; #100;
A = 16'h00FD; B = 16'h004A; #100;
A = 16'h00FD; B = 16'h004B; #100;
A = 16'h00FD; B = 16'h004C; #100;
A = 16'h00FD; B = 16'h004D; #100;
A = 16'h00FD; B = 16'h004E; #100;
A = 16'h00FD; B = 16'h004F; #100;
A = 16'h00FD; B = 16'h0050; #100;
A = 16'h00FD; B = 16'h0051; #100;
A = 16'h00FD; B = 16'h0052; #100;
A = 16'h00FD; B = 16'h0053; #100;
A = 16'h00FD; B = 16'h0054; #100;
A = 16'h00FD; B = 16'h0055; #100;
A = 16'h00FD; B = 16'h0056; #100;
A = 16'h00FD; B = 16'h0057; #100;
A = 16'h00FD; B = 16'h0058; #100;
A = 16'h00FD; B = 16'h0059; #100;
A = 16'h00FD; B = 16'h005A; #100;
A = 16'h00FD; B = 16'h005B; #100;
A = 16'h00FD; B = 16'h005C; #100;
A = 16'h00FD; B = 16'h005D; #100;
A = 16'h00FD; B = 16'h005E; #100;
A = 16'h00FD; B = 16'h005F; #100;
A = 16'h00FD; B = 16'h0060; #100;
A = 16'h00FD; B = 16'h0061; #100;
A = 16'h00FD; B = 16'h0062; #100;
A = 16'h00FD; B = 16'h0063; #100;
A = 16'h00FD; B = 16'h0064; #100;
A = 16'h00FD; B = 16'h0065; #100;
A = 16'h00FD; B = 16'h0066; #100;
A = 16'h00FD; B = 16'h0067; #100;
A = 16'h00FD; B = 16'h0068; #100;
A = 16'h00FD; B = 16'h0069; #100;
A = 16'h00FD; B = 16'h006A; #100;
A = 16'h00FD; B = 16'h006B; #100;
A = 16'h00FD; B = 16'h006C; #100;
A = 16'h00FD; B = 16'h006D; #100;
A = 16'h00FD; B = 16'h006E; #100;
A = 16'h00FD; B = 16'h006F; #100;
A = 16'h00FD; B = 16'h0070; #100;
A = 16'h00FD; B = 16'h0071; #100;
A = 16'h00FD; B = 16'h0072; #100;
A = 16'h00FD; B = 16'h0073; #100;
A = 16'h00FD; B = 16'h0074; #100;
A = 16'h00FD; B = 16'h0075; #100;
A = 16'h00FD; B = 16'h0076; #100;
A = 16'h00FD; B = 16'h0077; #100;
A = 16'h00FD; B = 16'h0078; #100;
A = 16'h00FD; B = 16'h0079; #100;
A = 16'h00FD; B = 16'h007A; #100;
A = 16'h00FD; B = 16'h007B; #100;
A = 16'h00FD; B = 16'h007C; #100;
A = 16'h00FD; B = 16'h007D; #100;
A = 16'h00FD; B = 16'h007E; #100;
A = 16'h00FD; B = 16'h007F; #100;
A = 16'h00FD; B = 16'h0080; #100;
A = 16'h00FD; B = 16'h0081; #100;
A = 16'h00FD; B = 16'h0082; #100;
A = 16'h00FD; B = 16'h0083; #100;
A = 16'h00FD; B = 16'h0084; #100;
A = 16'h00FD; B = 16'h0085; #100;
A = 16'h00FD; B = 16'h0086; #100;
A = 16'h00FD; B = 16'h0087; #100;
A = 16'h00FD; B = 16'h0088; #100;
A = 16'h00FD; B = 16'h0089; #100;
A = 16'h00FD; B = 16'h008A; #100;
A = 16'h00FD; B = 16'h008B; #100;
A = 16'h00FD; B = 16'h008C; #100;
A = 16'h00FD; B = 16'h008D; #100;
A = 16'h00FD; B = 16'h008E; #100;
A = 16'h00FD; B = 16'h008F; #100;
A = 16'h00FD; B = 16'h0090; #100;
A = 16'h00FD; B = 16'h0091; #100;
A = 16'h00FD; B = 16'h0092; #100;
A = 16'h00FD; B = 16'h0093; #100;
A = 16'h00FD; B = 16'h0094; #100;
A = 16'h00FD; B = 16'h0095; #100;
A = 16'h00FD; B = 16'h0096; #100;
A = 16'h00FD; B = 16'h0097; #100;
A = 16'h00FD; B = 16'h0098; #100;
A = 16'h00FD; B = 16'h0099; #100;
A = 16'h00FD; B = 16'h009A; #100;
A = 16'h00FD; B = 16'h009B; #100;
A = 16'h00FD; B = 16'h009C; #100;
A = 16'h00FD; B = 16'h009D; #100;
A = 16'h00FD; B = 16'h009E; #100;
A = 16'h00FD; B = 16'h009F; #100;
A = 16'h00FD; B = 16'h00A0; #100;
A = 16'h00FD; B = 16'h00A1; #100;
A = 16'h00FD; B = 16'h00A2; #100;
A = 16'h00FD; B = 16'h00A3; #100;
A = 16'h00FD; B = 16'h00A4; #100;
A = 16'h00FD; B = 16'h00A5; #100;
A = 16'h00FD; B = 16'h00A6; #100;
A = 16'h00FD; B = 16'h00A7; #100;
A = 16'h00FD; B = 16'h00A8; #100;
A = 16'h00FD; B = 16'h00A9; #100;
A = 16'h00FD; B = 16'h00AA; #100;
A = 16'h00FD; B = 16'h00AB; #100;
A = 16'h00FD; B = 16'h00AC; #100;
A = 16'h00FD; B = 16'h00AD; #100;
A = 16'h00FD; B = 16'h00AE; #100;
A = 16'h00FD; B = 16'h00AF; #100;
A = 16'h00FD; B = 16'h00B0; #100;
A = 16'h00FD; B = 16'h00B1; #100;
A = 16'h00FD; B = 16'h00B2; #100;
A = 16'h00FD; B = 16'h00B3; #100;
A = 16'h00FD; B = 16'h00B4; #100;
A = 16'h00FD; B = 16'h00B5; #100;
A = 16'h00FD; B = 16'h00B6; #100;
A = 16'h00FD; B = 16'h00B7; #100;
A = 16'h00FD; B = 16'h00B8; #100;
A = 16'h00FD; B = 16'h00B9; #100;
A = 16'h00FD; B = 16'h00BA; #100;
A = 16'h00FD; B = 16'h00BB; #100;
A = 16'h00FD; B = 16'h00BC; #100;
A = 16'h00FD; B = 16'h00BD; #100;
A = 16'h00FD; B = 16'h00BE; #100;
A = 16'h00FD; B = 16'h00BF; #100;
A = 16'h00FD; B = 16'h00C0; #100;
A = 16'h00FD; B = 16'h00C1; #100;
A = 16'h00FD; B = 16'h00C2; #100;
A = 16'h00FD; B = 16'h00C3; #100;
A = 16'h00FD; B = 16'h00C4; #100;
A = 16'h00FD; B = 16'h00C5; #100;
A = 16'h00FD; B = 16'h00C6; #100;
A = 16'h00FD; B = 16'h00C7; #100;
A = 16'h00FD; B = 16'h00C8; #100;
A = 16'h00FD; B = 16'h00C9; #100;
A = 16'h00FD; B = 16'h00CA; #100;
A = 16'h00FD; B = 16'h00CB; #100;
A = 16'h00FD; B = 16'h00CC; #100;
A = 16'h00FD; B = 16'h00CD; #100;
A = 16'h00FD; B = 16'h00CE; #100;
A = 16'h00FD; B = 16'h00CF; #100;
A = 16'h00FD; B = 16'h00D0; #100;
A = 16'h00FD; B = 16'h00D1; #100;
A = 16'h00FD; B = 16'h00D2; #100;
A = 16'h00FD; B = 16'h00D3; #100;
A = 16'h00FD; B = 16'h00D4; #100;
A = 16'h00FD; B = 16'h00D5; #100;
A = 16'h00FD; B = 16'h00D6; #100;
A = 16'h00FD; B = 16'h00D7; #100;
A = 16'h00FD; B = 16'h00D8; #100;
A = 16'h00FD; B = 16'h00D9; #100;
A = 16'h00FD; B = 16'h00DA; #100;
A = 16'h00FD; B = 16'h00DB; #100;
A = 16'h00FD; B = 16'h00DC; #100;
A = 16'h00FD; B = 16'h00DD; #100;
A = 16'h00FD; B = 16'h00DE; #100;
A = 16'h00FD; B = 16'h00DF; #100;
A = 16'h00FD; B = 16'h00E0; #100;
A = 16'h00FD; B = 16'h00E1; #100;
A = 16'h00FD; B = 16'h00E2; #100;
A = 16'h00FD; B = 16'h00E3; #100;
A = 16'h00FD; B = 16'h00E4; #100;
A = 16'h00FD; B = 16'h00E5; #100;
A = 16'h00FD; B = 16'h00E6; #100;
A = 16'h00FD; B = 16'h00E7; #100;
A = 16'h00FD; B = 16'h00E8; #100;
A = 16'h00FD; B = 16'h00E9; #100;
A = 16'h00FD; B = 16'h00EA; #100;
A = 16'h00FD; B = 16'h00EB; #100;
A = 16'h00FD; B = 16'h00EC; #100;
A = 16'h00FD; B = 16'h00ED; #100;
A = 16'h00FD; B = 16'h00EE; #100;
A = 16'h00FD; B = 16'h00EF; #100;
A = 16'h00FD; B = 16'h00F0; #100;
A = 16'h00FD; B = 16'h00F1; #100;
A = 16'h00FD; B = 16'h00F2; #100;
A = 16'h00FD; B = 16'h00F3; #100;
A = 16'h00FD; B = 16'h00F4; #100;
A = 16'h00FD; B = 16'h00F5; #100;
A = 16'h00FD; B = 16'h00F6; #100;
A = 16'h00FD; B = 16'h00F7; #100;
A = 16'h00FD; B = 16'h00F8; #100;
A = 16'h00FD; B = 16'h00F9; #100;
A = 16'h00FD; B = 16'h00FA; #100;
A = 16'h00FD; B = 16'h00FB; #100;
A = 16'h00FD; B = 16'h00FC; #100;
A = 16'h00FD; B = 16'h00FD; #100;
A = 16'h00FD; B = 16'h00FE; #100;
A = 16'h00FD; B = 16'h00FF; #100;
A = 16'h00FE; B = 16'h000; #100;
A = 16'h00FE; B = 16'h001; #100;
A = 16'h00FE; B = 16'h002; #100;
A = 16'h00FE; B = 16'h003; #100;
A = 16'h00FE; B = 16'h004; #100;
A = 16'h00FE; B = 16'h005; #100;
A = 16'h00FE; B = 16'h006; #100;
A = 16'h00FE; B = 16'h007; #100;
A = 16'h00FE; B = 16'h008; #100;
A = 16'h00FE; B = 16'h009; #100;
A = 16'h00FE; B = 16'h00A; #100;
A = 16'h00FE; B = 16'h00B; #100;
A = 16'h00FE; B = 16'h00C; #100;
A = 16'h00FE; B = 16'h00D; #100;
A = 16'h00FE; B = 16'h00E; #100;
A = 16'h00FE; B = 16'h00F; #100;
A = 16'h00FE; B = 16'h0010; #100;
A = 16'h00FE; B = 16'h0011; #100;
A = 16'h00FE; B = 16'h0012; #100;
A = 16'h00FE; B = 16'h0013; #100;
A = 16'h00FE; B = 16'h0014; #100;
A = 16'h00FE; B = 16'h0015; #100;
A = 16'h00FE; B = 16'h0016; #100;
A = 16'h00FE; B = 16'h0017; #100;
A = 16'h00FE; B = 16'h0018; #100;
A = 16'h00FE; B = 16'h0019; #100;
A = 16'h00FE; B = 16'h001A; #100;
A = 16'h00FE; B = 16'h001B; #100;
A = 16'h00FE; B = 16'h001C; #100;
A = 16'h00FE; B = 16'h001D; #100;
A = 16'h00FE; B = 16'h001E; #100;
A = 16'h00FE; B = 16'h001F; #100;
A = 16'h00FE; B = 16'h0020; #100;
A = 16'h00FE; B = 16'h0021; #100;
A = 16'h00FE; B = 16'h0022; #100;
A = 16'h00FE; B = 16'h0023; #100;
A = 16'h00FE; B = 16'h0024; #100;
A = 16'h00FE; B = 16'h0025; #100;
A = 16'h00FE; B = 16'h0026; #100;
A = 16'h00FE; B = 16'h0027; #100;
A = 16'h00FE; B = 16'h0028; #100;
A = 16'h00FE; B = 16'h0029; #100;
A = 16'h00FE; B = 16'h002A; #100;
A = 16'h00FE; B = 16'h002B; #100;
A = 16'h00FE; B = 16'h002C; #100;
A = 16'h00FE; B = 16'h002D; #100;
A = 16'h00FE; B = 16'h002E; #100;
A = 16'h00FE; B = 16'h002F; #100;
A = 16'h00FE; B = 16'h0030; #100;
A = 16'h00FE; B = 16'h0031; #100;
A = 16'h00FE; B = 16'h0032; #100;
A = 16'h00FE; B = 16'h0033; #100;
A = 16'h00FE; B = 16'h0034; #100;
A = 16'h00FE; B = 16'h0035; #100;
A = 16'h00FE; B = 16'h0036; #100;
A = 16'h00FE; B = 16'h0037; #100;
A = 16'h00FE; B = 16'h0038; #100;
A = 16'h00FE; B = 16'h0039; #100;
A = 16'h00FE; B = 16'h003A; #100;
A = 16'h00FE; B = 16'h003B; #100;
A = 16'h00FE; B = 16'h003C; #100;
A = 16'h00FE; B = 16'h003D; #100;
A = 16'h00FE; B = 16'h003E; #100;
A = 16'h00FE; B = 16'h003F; #100;
A = 16'h00FE; B = 16'h0040; #100;
A = 16'h00FE; B = 16'h0041; #100;
A = 16'h00FE; B = 16'h0042; #100;
A = 16'h00FE; B = 16'h0043; #100;
A = 16'h00FE; B = 16'h0044; #100;
A = 16'h00FE; B = 16'h0045; #100;
A = 16'h00FE; B = 16'h0046; #100;
A = 16'h00FE; B = 16'h0047; #100;
A = 16'h00FE; B = 16'h0048; #100;
A = 16'h00FE; B = 16'h0049; #100;
A = 16'h00FE; B = 16'h004A; #100;
A = 16'h00FE; B = 16'h004B; #100;
A = 16'h00FE; B = 16'h004C; #100;
A = 16'h00FE; B = 16'h004D; #100;
A = 16'h00FE; B = 16'h004E; #100;
A = 16'h00FE; B = 16'h004F; #100;
A = 16'h00FE; B = 16'h0050; #100;
A = 16'h00FE; B = 16'h0051; #100;
A = 16'h00FE; B = 16'h0052; #100;
A = 16'h00FE; B = 16'h0053; #100;
A = 16'h00FE; B = 16'h0054; #100;
A = 16'h00FE; B = 16'h0055; #100;
A = 16'h00FE; B = 16'h0056; #100;
A = 16'h00FE; B = 16'h0057; #100;
A = 16'h00FE; B = 16'h0058; #100;
A = 16'h00FE; B = 16'h0059; #100;
A = 16'h00FE; B = 16'h005A; #100;
A = 16'h00FE; B = 16'h005B; #100;
A = 16'h00FE; B = 16'h005C; #100;
A = 16'h00FE; B = 16'h005D; #100;
A = 16'h00FE; B = 16'h005E; #100;
A = 16'h00FE; B = 16'h005F; #100;
A = 16'h00FE; B = 16'h0060; #100;
A = 16'h00FE; B = 16'h0061; #100;
A = 16'h00FE; B = 16'h0062; #100;
A = 16'h00FE; B = 16'h0063; #100;
A = 16'h00FE; B = 16'h0064; #100;
A = 16'h00FE; B = 16'h0065; #100;
A = 16'h00FE; B = 16'h0066; #100;
A = 16'h00FE; B = 16'h0067; #100;
A = 16'h00FE; B = 16'h0068; #100;
A = 16'h00FE; B = 16'h0069; #100;
A = 16'h00FE; B = 16'h006A; #100;
A = 16'h00FE; B = 16'h006B; #100;
A = 16'h00FE; B = 16'h006C; #100;
A = 16'h00FE; B = 16'h006D; #100;
A = 16'h00FE; B = 16'h006E; #100;
A = 16'h00FE; B = 16'h006F; #100;
A = 16'h00FE; B = 16'h0070; #100;
A = 16'h00FE; B = 16'h0071; #100;
A = 16'h00FE; B = 16'h0072; #100;
A = 16'h00FE; B = 16'h0073; #100;
A = 16'h00FE; B = 16'h0074; #100;
A = 16'h00FE; B = 16'h0075; #100;
A = 16'h00FE; B = 16'h0076; #100;
A = 16'h00FE; B = 16'h0077; #100;
A = 16'h00FE; B = 16'h0078; #100;
A = 16'h00FE; B = 16'h0079; #100;
A = 16'h00FE; B = 16'h007A; #100;
A = 16'h00FE; B = 16'h007B; #100;
A = 16'h00FE; B = 16'h007C; #100;
A = 16'h00FE; B = 16'h007D; #100;
A = 16'h00FE; B = 16'h007E; #100;
A = 16'h00FE; B = 16'h007F; #100;
A = 16'h00FE; B = 16'h0080; #100;
A = 16'h00FE; B = 16'h0081; #100;
A = 16'h00FE; B = 16'h0082; #100;
A = 16'h00FE; B = 16'h0083; #100;
A = 16'h00FE; B = 16'h0084; #100;
A = 16'h00FE; B = 16'h0085; #100;
A = 16'h00FE; B = 16'h0086; #100;
A = 16'h00FE; B = 16'h0087; #100;
A = 16'h00FE; B = 16'h0088; #100;
A = 16'h00FE; B = 16'h0089; #100;
A = 16'h00FE; B = 16'h008A; #100;
A = 16'h00FE; B = 16'h008B; #100;
A = 16'h00FE; B = 16'h008C; #100;
A = 16'h00FE; B = 16'h008D; #100;
A = 16'h00FE; B = 16'h008E; #100;
A = 16'h00FE; B = 16'h008F; #100;
A = 16'h00FE; B = 16'h0090; #100;
A = 16'h00FE; B = 16'h0091; #100;
A = 16'h00FE; B = 16'h0092; #100;
A = 16'h00FE; B = 16'h0093; #100;
A = 16'h00FE; B = 16'h0094; #100;
A = 16'h00FE; B = 16'h0095; #100;
A = 16'h00FE; B = 16'h0096; #100;
A = 16'h00FE; B = 16'h0097; #100;
A = 16'h00FE; B = 16'h0098; #100;
A = 16'h00FE; B = 16'h0099; #100;
A = 16'h00FE; B = 16'h009A; #100;
A = 16'h00FE; B = 16'h009B; #100;
A = 16'h00FE; B = 16'h009C; #100;
A = 16'h00FE; B = 16'h009D; #100;
A = 16'h00FE; B = 16'h009E; #100;
A = 16'h00FE; B = 16'h009F; #100;
A = 16'h00FE; B = 16'h00A0; #100;
A = 16'h00FE; B = 16'h00A1; #100;
A = 16'h00FE; B = 16'h00A2; #100;
A = 16'h00FE; B = 16'h00A3; #100;
A = 16'h00FE; B = 16'h00A4; #100;
A = 16'h00FE; B = 16'h00A5; #100;
A = 16'h00FE; B = 16'h00A6; #100;
A = 16'h00FE; B = 16'h00A7; #100;
A = 16'h00FE; B = 16'h00A8; #100;
A = 16'h00FE; B = 16'h00A9; #100;
A = 16'h00FE; B = 16'h00AA; #100;
A = 16'h00FE; B = 16'h00AB; #100;
A = 16'h00FE; B = 16'h00AC; #100;
A = 16'h00FE; B = 16'h00AD; #100;
A = 16'h00FE; B = 16'h00AE; #100;
A = 16'h00FE; B = 16'h00AF; #100;
A = 16'h00FE; B = 16'h00B0; #100;
A = 16'h00FE; B = 16'h00B1; #100;
A = 16'h00FE; B = 16'h00B2; #100;
A = 16'h00FE; B = 16'h00B3; #100;
A = 16'h00FE; B = 16'h00B4; #100;
A = 16'h00FE; B = 16'h00B5; #100;
A = 16'h00FE; B = 16'h00B6; #100;
A = 16'h00FE; B = 16'h00B7; #100;
A = 16'h00FE; B = 16'h00B8; #100;
A = 16'h00FE; B = 16'h00B9; #100;
A = 16'h00FE; B = 16'h00BA; #100;
A = 16'h00FE; B = 16'h00BB; #100;
A = 16'h00FE; B = 16'h00BC; #100;
A = 16'h00FE; B = 16'h00BD; #100;
A = 16'h00FE; B = 16'h00BE; #100;
A = 16'h00FE; B = 16'h00BF; #100;
A = 16'h00FE; B = 16'h00C0; #100;
A = 16'h00FE; B = 16'h00C1; #100;
A = 16'h00FE; B = 16'h00C2; #100;
A = 16'h00FE; B = 16'h00C3; #100;
A = 16'h00FE; B = 16'h00C4; #100;
A = 16'h00FE; B = 16'h00C5; #100;
A = 16'h00FE; B = 16'h00C6; #100;
A = 16'h00FE; B = 16'h00C7; #100;
A = 16'h00FE; B = 16'h00C8; #100;
A = 16'h00FE; B = 16'h00C9; #100;
A = 16'h00FE; B = 16'h00CA; #100;
A = 16'h00FE; B = 16'h00CB; #100;
A = 16'h00FE; B = 16'h00CC; #100;
A = 16'h00FE; B = 16'h00CD; #100;
A = 16'h00FE; B = 16'h00CE; #100;
A = 16'h00FE; B = 16'h00CF; #100;
A = 16'h00FE; B = 16'h00D0; #100;
A = 16'h00FE; B = 16'h00D1; #100;
A = 16'h00FE; B = 16'h00D2; #100;
A = 16'h00FE; B = 16'h00D3; #100;
A = 16'h00FE; B = 16'h00D4; #100;
A = 16'h00FE; B = 16'h00D5; #100;
A = 16'h00FE; B = 16'h00D6; #100;
A = 16'h00FE; B = 16'h00D7; #100;
A = 16'h00FE; B = 16'h00D8; #100;
A = 16'h00FE; B = 16'h00D9; #100;
A = 16'h00FE; B = 16'h00DA; #100;
A = 16'h00FE; B = 16'h00DB; #100;
A = 16'h00FE; B = 16'h00DC; #100;
A = 16'h00FE; B = 16'h00DD; #100;
A = 16'h00FE; B = 16'h00DE; #100;
A = 16'h00FE; B = 16'h00DF; #100;
A = 16'h00FE; B = 16'h00E0; #100;
A = 16'h00FE; B = 16'h00E1; #100;
A = 16'h00FE; B = 16'h00E2; #100;
A = 16'h00FE; B = 16'h00E3; #100;
A = 16'h00FE; B = 16'h00E4; #100;
A = 16'h00FE; B = 16'h00E5; #100;
A = 16'h00FE; B = 16'h00E6; #100;
A = 16'h00FE; B = 16'h00E7; #100;
A = 16'h00FE; B = 16'h00E8; #100;
A = 16'h00FE; B = 16'h00E9; #100;
A = 16'h00FE; B = 16'h00EA; #100;
A = 16'h00FE; B = 16'h00EB; #100;
A = 16'h00FE; B = 16'h00EC; #100;
A = 16'h00FE; B = 16'h00ED; #100;
A = 16'h00FE; B = 16'h00EE; #100;
A = 16'h00FE; B = 16'h00EF; #100;
A = 16'h00FE; B = 16'h00F0; #100;
A = 16'h00FE; B = 16'h00F1; #100;
A = 16'h00FE; B = 16'h00F2; #100;
A = 16'h00FE; B = 16'h00F3; #100;
A = 16'h00FE; B = 16'h00F4; #100;
A = 16'h00FE; B = 16'h00F5; #100;
A = 16'h00FE; B = 16'h00F6; #100;
A = 16'h00FE; B = 16'h00F7; #100;
A = 16'h00FE; B = 16'h00F8; #100;
A = 16'h00FE; B = 16'h00F9; #100;
A = 16'h00FE; B = 16'h00FA; #100;
A = 16'h00FE; B = 16'h00FB; #100;
A = 16'h00FE; B = 16'h00FC; #100;
A = 16'h00FE; B = 16'h00FD; #100;
A = 16'h00FE; B = 16'h00FE; #100;
A = 16'h00FE; B = 16'h00FF; #100;
A = 16'h00FF; B = 16'h000; #100;
A = 16'h00FF; B = 16'h001; #100;
A = 16'h00FF; B = 16'h002; #100;
A = 16'h00FF; B = 16'h003; #100;
A = 16'h00FF; B = 16'h004; #100;
A = 16'h00FF; B = 16'h005; #100;
A = 16'h00FF; B = 16'h006; #100;
A = 16'h00FF; B = 16'h007; #100;
A = 16'h00FF; B = 16'h008; #100;
A = 16'h00FF; B = 16'h009; #100;
A = 16'h00FF; B = 16'h00A; #100;
A = 16'h00FF; B = 16'h00B; #100;
A = 16'h00FF; B = 16'h00C; #100;
A = 16'h00FF; B = 16'h00D; #100;
A = 16'h00FF; B = 16'h00E; #100;
A = 16'h00FF; B = 16'h00F; #100;
A = 16'h00FF; B = 16'h0010; #100;
A = 16'h00FF; B = 16'h0011; #100;
A = 16'h00FF; B = 16'h0012; #100;
A = 16'h00FF; B = 16'h0013; #100;
A = 16'h00FF; B = 16'h0014; #100;
A = 16'h00FF; B = 16'h0015; #100;
A = 16'h00FF; B = 16'h0016; #100;
A = 16'h00FF; B = 16'h0017; #100;
A = 16'h00FF; B = 16'h0018; #100;
A = 16'h00FF; B = 16'h0019; #100;
A = 16'h00FF; B = 16'h001A; #100;
A = 16'h00FF; B = 16'h001B; #100;
A = 16'h00FF; B = 16'h001C; #100;
A = 16'h00FF; B = 16'h001D; #100;
A = 16'h00FF; B = 16'h001E; #100;
A = 16'h00FF; B = 16'h001F; #100;
A = 16'h00FF; B = 16'h0020; #100;
A = 16'h00FF; B = 16'h0021; #100;
A = 16'h00FF; B = 16'h0022; #100;
A = 16'h00FF; B = 16'h0023; #100;
A = 16'h00FF; B = 16'h0024; #100;
A = 16'h00FF; B = 16'h0025; #100;
A = 16'h00FF; B = 16'h0026; #100;
A = 16'h00FF; B = 16'h0027; #100;
A = 16'h00FF; B = 16'h0028; #100;
A = 16'h00FF; B = 16'h0029; #100;
A = 16'h00FF; B = 16'h002A; #100;
A = 16'h00FF; B = 16'h002B; #100;
A = 16'h00FF; B = 16'h002C; #100;
A = 16'h00FF; B = 16'h002D; #100;
A = 16'h00FF; B = 16'h002E; #100;
A = 16'h00FF; B = 16'h002F; #100;
A = 16'h00FF; B = 16'h0030; #100;
A = 16'h00FF; B = 16'h0031; #100;
A = 16'h00FF; B = 16'h0032; #100;
A = 16'h00FF; B = 16'h0033; #100;
A = 16'h00FF; B = 16'h0034; #100;
A = 16'h00FF; B = 16'h0035; #100;
A = 16'h00FF; B = 16'h0036; #100;
A = 16'h00FF; B = 16'h0037; #100;
A = 16'h00FF; B = 16'h0038; #100;
A = 16'h00FF; B = 16'h0039; #100;
A = 16'h00FF; B = 16'h003A; #100;
A = 16'h00FF; B = 16'h003B; #100;
A = 16'h00FF; B = 16'h003C; #100;
A = 16'h00FF; B = 16'h003D; #100;
A = 16'h00FF; B = 16'h003E; #100;
A = 16'h00FF; B = 16'h003F; #100;
A = 16'h00FF; B = 16'h0040; #100;
A = 16'h00FF; B = 16'h0041; #100;
A = 16'h00FF; B = 16'h0042; #100;
A = 16'h00FF; B = 16'h0043; #100;
A = 16'h00FF; B = 16'h0044; #100;
A = 16'h00FF; B = 16'h0045; #100;
A = 16'h00FF; B = 16'h0046; #100;
A = 16'h00FF; B = 16'h0047; #100;
A = 16'h00FF; B = 16'h0048; #100;
A = 16'h00FF; B = 16'h0049; #100;
A = 16'h00FF; B = 16'h004A; #100;
A = 16'h00FF; B = 16'h004B; #100;
A = 16'h00FF; B = 16'h004C; #100;
A = 16'h00FF; B = 16'h004D; #100;
A = 16'h00FF; B = 16'h004E; #100;
A = 16'h00FF; B = 16'h004F; #100;
A = 16'h00FF; B = 16'h0050; #100;
A = 16'h00FF; B = 16'h0051; #100;
A = 16'h00FF; B = 16'h0052; #100;
A = 16'h00FF; B = 16'h0053; #100;
A = 16'h00FF; B = 16'h0054; #100;
A = 16'h00FF; B = 16'h0055; #100;
A = 16'h00FF; B = 16'h0056; #100;
A = 16'h00FF; B = 16'h0057; #100;
A = 16'h00FF; B = 16'h0058; #100;
A = 16'h00FF; B = 16'h0059; #100;
A = 16'h00FF; B = 16'h005A; #100;
A = 16'h00FF; B = 16'h005B; #100;
A = 16'h00FF; B = 16'h005C; #100;
A = 16'h00FF; B = 16'h005D; #100;
A = 16'h00FF; B = 16'h005E; #100;
A = 16'h00FF; B = 16'h005F; #100;
A = 16'h00FF; B = 16'h0060; #100;
A = 16'h00FF; B = 16'h0061; #100;
A = 16'h00FF; B = 16'h0062; #100;
A = 16'h00FF; B = 16'h0063; #100;
A = 16'h00FF; B = 16'h0064; #100;
A = 16'h00FF; B = 16'h0065; #100;
A = 16'h00FF; B = 16'h0066; #100;
A = 16'h00FF; B = 16'h0067; #100;
A = 16'h00FF; B = 16'h0068; #100;
A = 16'h00FF; B = 16'h0069; #100;
A = 16'h00FF; B = 16'h006A; #100;
A = 16'h00FF; B = 16'h006B; #100;
A = 16'h00FF; B = 16'h006C; #100;
A = 16'h00FF; B = 16'h006D; #100;
A = 16'h00FF; B = 16'h006E; #100;
A = 16'h00FF; B = 16'h006F; #100;
A = 16'h00FF; B = 16'h0070; #100;
A = 16'h00FF; B = 16'h0071; #100;
A = 16'h00FF; B = 16'h0072; #100;
A = 16'h00FF; B = 16'h0073; #100;
A = 16'h00FF; B = 16'h0074; #100;
A = 16'h00FF; B = 16'h0075; #100;
A = 16'h00FF; B = 16'h0076; #100;
A = 16'h00FF; B = 16'h0077; #100;
A = 16'h00FF; B = 16'h0078; #100;
A = 16'h00FF; B = 16'h0079; #100;
A = 16'h00FF; B = 16'h007A; #100;
A = 16'h00FF; B = 16'h007B; #100;
A = 16'h00FF; B = 16'h007C; #100;
A = 16'h00FF; B = 16'h007D; #100;
A = 16'h00FF; B = 16'h007E; #100;
A = 16'h00FF; B = 16'h007F; #100;
A = 16'h00FF; B = 16'h0080; #100;
A = 16'h00FF; B = 16'h0081; #100;
A = 16'h00FF; B = 16'h0082; #100;
A = 16'h00FF; B = 16'h0083; #100;
A = 16'h00FF; B = 16'h0084; #100;
A = 16'h00FF; B = 16'h0085; #100;
A = 16'h00FF; B = 16'h0086; #100;
A = 16'h00FF; B = 16'h0087; #100;
A = 16'h00FF; B = 16'h0088; #100;
A = 16'h00FF; B = 16'h0089; #100;
A = 16'h00FF; B = 16'h008A; #100;
A = 16'h00FF; B = 16'h008B; #100;
A = 16'h00FF; B = 16'h008C; #100;
A = 16'h00FF; B = 16'h008D; #100;
A = 16'h00FF; B = 16'h008E; #100;
A = 16'h00FF; B = 16'h008F; #100;
A = 16'h00FF; B = 16'h0090; #100;
A = 16'h00FF; B = 16'h0091; #100;
A = 16'h00FF; B = 16'h0092; #100;
A = 16'h00FF; B = 16'h0093; #100;
A = 16'h00FF; B = 16'h0094; #100;
A = 16'h00FF; B = 16'h0095; #100;
A = 16'h00FF; B = 16'h0096; #100;
A = 16'h00FF; B = 16'h0097; #100;
A = 16'h00FF; B = 16'h0098; #100;
A = 16'h00FF; B = 16'h0099; #100;
A = 16'h00FF; B = 16'h009A; #100;
A = 16'h00FF; B = 16'h009B; #100;
A = 16'h00FF; B = 16'h009C; #100;
A = 16'h00FF; B = 16'h009D; #100;
A = 16'h00FF; B = 16'h009E; #100;
A = 16'h00FF; B = 16'h009F; #100;
A = 16'h00FF; B = 16'h00A0; #100;
A = 16'h00FF; B = 16'h00A1; #100;
A = 16'h00FF; B = 16'h00A2; #100;
A = 16'h00FF; B = 16'h00A3; #100;
A = 16'h00FF; B = 16'h00A4; #100;
A = 16'h00FF; B = 16'h00A5; #100;
A = 16'h00FF; B = 16'h00A6; #100;
A = 16'h00FF; B = 16'h00A7; #100;
A = 16'h00FF; B = 16'h00A8; #100;
A = 16'h00FF; B = 16'h00A9; #100;
A = 16'h00FF; B = 16'h00AA; #100;
A = 16'h00FF; B = 16'h00AB; #100;
A = 16'h00FF; B = 16'h00AC; #100;
A = 16'h00FF; B = 16'h00AD; #100;
A = 16'h00FF; B = 16'h00AE; #100;
A = 16'h00FF; B = 16'h00AF; #100;
A = 16'h00FF; B = 16'h00B0; #100;
A = 16'h00FF; B = 16'h00B1; #100;
A = 16'h00FF; B = 16'h00B2; #100;
A = 16'h00FF; B = 16'h00B3; #100;
A = 16'h00FF; B = 16'h00B4; #100;
A = 16'h00FF; B = 16'h00B5; #100;
A = 16'h00FF; B = 16'h00B6; #100;
A = 16'h00FF; B = 16'h00B7; #100;
A = 16'h00FF; B = 16'h00B8; #100;
A = 16'h00FF; B = 16'h00B9; #100;
A = 16'h00FF; B = 16'h00BA; #100;
A = 16'h00FF; B = 16'h00BB; #100;
A = 16'h00FF; B = 16'h00BC; #100;
A = 16'h00FF; B = 16'h00BD; #100;
A = 16'h00FF; B = 16'h00BE; #100;
A = 16'h00FF; B = 16'h00BF; #100;
A = 16'h00FF; B = 16'h00C0; #100;
A = 16'h00FF; B = 16'h00C1; #100;
A = 16'h00FF; B = 16'h00C2; #100;
A = 16'h00FF; B = 16'h00C3; #100;
A = 16'h00FF; B = 16'h00C4; #100;
A = 16'h00FF; B = 16'h00C5; #100;
A = 16'h00FF; B = 16'h00C6; #100;
A = 16'h00FF; B = 16'h00C7; #100;
A = 16'h00FF; B = 16'h00C8; #100;
A = 16'h00FF; B = 16'h00C9; #100;
A = 16'h00FF; B = 16'h00CA; #100;
A = 16'h00FF; B = 16'h00CB; #100;
A = 16'h00FF; B = 16'h00CC; #100;
A = 16'h00FF; B = 16'h00CD; #100;
A = 16'h00FF; B = 16'h00CE; #100;
A = 16'h00FF; B = 16'h00CF; #100;
A = 16'h00FF; B = 16'h00D0; #100;
A = 16'h00FF; B = 16'h00D1; #100;
A = 16'h00FF; B = 16'h00D2; #100;
A = 16'h00FF; B = 16'h00D3; #100;
A = 16'h00FF; B = 16'h00D4; #100;
A = 16'h00FF; B = 16'h00D5; #100;
A = 16'h00FF; B = 16'h00D6; #100;
A = 16'h00FF; B = 16'h00D7; #100;
A = 16'h00FF; B = 16'h00D8; #100;
A = 16'h00FF; B = 16'h00D9; #100;
A = 16'h00FF; B = 16'h00DA; #100;
A = 16'h00FF; B = 16'h00DB; #100;
A = 16'h00FF; B = 16'h00DC; #100;
A = 16'h00FF; B = 16'h00DD; #100;
A = 16'h00FF; B = 16'h00DE; #100;
A = 16'h00FF; B = 16'h00DF; #100;
A = 16'h00FF; B = 16'h00E0; #100;
A = 16'h00FF; B = 16'h00E1; #100;
A = 16'h00FF; B = 16'h00E2; #100;
A = 16'h00FF; B = 16'h00E3; #100;
A = 16'h00FF; B = 16'h00E4; #100;
A = 16'h00FF; B = 16'h00E5; #100;
A = 16'h00FF; B = 16'h00E6; #100;
A = 16'h00FF; B = 16'h00E7; #100;
A = 16'h00FF; B = 16'h00E8; #100;
A = 16'h00FF; B = 16'h00E9; #100;
A = 16'h00FF; B = 16'h00EA; #100;
A = 16'h00FF; B = 16'h00EB; #100;
A = 16'h00FF; B = 16'h00EC; #100;
A = 16'h00FF; B = 16'h00ED; #100;
A = 16'h00FF; B = 16'h00EE; #100;
A = 16'h00FF; B = 16'h00EF; #100;
A = 16'h00FF; B = 16'h00F0; #100;
A = 16'h00FF; B = 16'h00F1; #100;
A = 16'h00FF; B = 16'h00F2; #100;
A = 16'h00FF; B = 16'h00F3; #100;
A = 16'h00FF; B = 16'h00F4; #100;
A = 16'h00FF; B = 16'h00F5; #100;
A = 16'h00FF; B = 16'h00F6; #100;
A = 16'h00FF; B = 16'h00F7; #100;
A = 16'h00FF; B = 16'h00F8; #100;
A = 16'h00FF; B = 16'h00F9; #100;
A = 16'h00FF; B = 16'h00FA; #100;
A = 16'h00FF; B = 16'h00FB; #100;
A = 16'h00FF; B = 16'h00FC; #100;
A = 16'h00FF; B = 16'h00FD; #100;
A = 16'h00FF; B = 16'h00FE; #100;
A = 16'h00FF; B = 16'h00FF; #100;
A = 16'hFFFF; B = 16'h0001; #100;  // Desbordamiento, resultado esperado: 0x0000, Cout = 1
A = 16'h8000; B = 16'h8000; #100;  // Suma de valores m�ximos en signo negativo, resultado esperado: 0x0000, Cout = 1
A = 16'h7FFF; B = 16'h0001; #100;  // Desbordamiento en positivo, resultado esperado: 0x8000, Cout = 0
A = 16'hFFFF; B = 16'hFFFF; #100;  // Caso de todos unos, resultado esperado: 0xFFFE, Cout = 1
A = 16'h1234; B = 16'h4321; #100;  // Suma arbitraria, resultado esperado: 0x5555, Cout = 0
A = 16'hFFFF; B = 16'h7FFF; #100;  // Desbordamiento sin acarreo, resultado esperado: 0x7FFE, Cout = 1
A = 16'h8000; B = 16'h7FFF; #100;  // Valores m�ximos y m�nimos, resultado esperado: 0xFFFF, Cout = 0
A = 16'h0001; B = 16'hFFFF; #100;  // Desbordamiento en un extremo, resultado esperado: 0x0000, Cout = 1
A = 16'hAAAA; B = 16'h5555; #100;  // Alternancia de bits, resultado esperado: 0xFFFF, Cout = 0





	$stop;
end


endmodule 